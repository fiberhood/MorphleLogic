VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 2.400 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 2.400 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 2.400 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 2.400 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 2.400 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 2.400 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 2.400 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 2.400 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 2.400 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 2.400 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 2.400 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 2.400 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 2.400 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 468.095 2910.335 469.645 ;
      LAYER mcon ;
        RECT 2910.105 468.265 2910.275 468.435 ;
      LAYER met1 ;
        RECT 2910.045 468.420 2910.335 468.465 ;
        RECT 2906.300 468.280 2910.335 468.420 ;
        RECT 2910.045 468.235 2910.335 468.280 ;
      LAYER met3 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2906.300 204.870 2924.800 205.170 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 2774.655 2910.335 2776.205 ;
      LAYER mcon ;
        RECT 2910.105 2774.825 2910.275 2774.995 ;
      LAYER met1 ;
        RECT 2910.045 2774.980 2910.335 2775.025 ;
        RECT 2906.300 2774.840 2910.335 2774.980 ;
        RECT 2910.045 2774.795 2910.335 2774.840 ;
      LAYER met3 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2906.300 2551.550 2924.800 2551.850 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 2627.775 2910.335 2629.325 ;
      LAYER mcon ;
        RECT 2910.105 2628.625 2910.275 2628.795 ;
      LAYER met1 ;
        RECT 2910.045 2628.780 2910.335 2628.825 ;
        RECT 2906.300 2628.640 2910.335 2628.780 ;
        RECT 2910.045 2628.595 2910.335 2628.640 ;
      LAYER met3 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2906.300 2786.150 2924.800 2786.450 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2911.195 2914.035 2911.715 2915.585 ;
      LAYER mcon ;
        RECT 2911.485 2915.245 2911.655 2915.415 ;
      LAYER met1 ;
        RECT 2911.425 2915.400 2911.715 2915.445 ;
        RECT 2906.300 2915.260 2911.715 2915.400 ;
        RECT 2911.425 2915.215 2911.715 2915.260 ;
      LAYER met3 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2906.300 3020.750 2924.800 3021.050 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2911.195 3202.355 2911.715 3203.905 ;
      LAYER mcon ;
        RECT 2911.485 3203.565 2911.655 3203.735 ;
      LAYER met1 ;
        RECT 2911.410 3203.720 2911.730 3203.780 ;
        RECT 2911.215 3203.580 2911.730 3203.720 ;
        RECT 2911.410 3203.520 2911.730 3203.580 ;
      LAYER via ;
        RECT 2911.440 3203.520 2911.700 3203.780 ;
      LAYER met2 ;
        RECT 2911.430 3255.315 2911.710 3255.685 ;
        RECT 2911.500 3203.810 2911.640 3255.315 ;
        RECT 2911.440 3203.490 2911.700 3203.810 ;
      LAYER via2 ;
        RECT 2911.430 3255.360 2911.710 3255.640 ;
      LAYER met3 ;
        RECT 2911.405 3255.650 2911.735 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2911.405 3255.350 2924.800 3255.650 ;
        RECT 2911.405 3255.335 2911.735 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 3095.615 2910.335 3097.165 ;
      LAYER mcon ;
        RECT 2910.105 3096.805 2910.275 3096.975 ;
      LAYER met1 ;
        RECT 2910.045 3096.960 2910.335 3097.005 ;
        RECT 2906.300 3096.820 2910.335 3096.960 ;
        RECT 2910.045 3096.775 2910.335 3096.820 ;
      LAYER met3 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2906.300 3489.950 2924.800 3490.250 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2911.195 3503.615 2911.715 3505.165 ;
      LAYER mcon ;
        RECT 2911.485 3504.465 2911.655 3504.635 ;
      LAYER met1 ;
        RECT 2911.425 3504.620 2911.715 3504.665 ;
        RECT 2906.300 3504.480 2911.715 3504.620 ;
        RECT 2911.425 3504.435 2911.715 3504.480 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3506.300 2636.100 3517.600 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3506.300 2311.800 3517.600 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3506.300 1987.500 3517.600 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3506.300 1662.740 3517.600 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3506.300 1338.440 3517.600 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 288.575 2910.335 290.125 ;
      LAYER mcon ;
        RECT 2910.105 289.425 2910.275 289.595 ;
      LAYER met1 ;
        RECT 2910.045 289.580 2910.335 289.625 ;
        RECT 2906.300 289.440 2910.335 289.580 ;
        RECT 2910.045 289.395 2910.335 289.440 ;
      LAYER met3 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2906.300 439.470 2924.800 439.770 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3506.300 1014.140 3517.600 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3506.300 689.380 3517.600 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3509.890 365.080 3517.600 ;
        RECT 363.100 3509.750 365.080 3509.890 ;
        RECT 363.100 3506.300 363.240 3509.750 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 11.815 3503.615 12.335 3505.165 ;
      LAYER mcon ;
        RECT 12.105 3504.805 12.275 3504.975 ;
      LAYER met1 ;
        RECT 12.045 3504.960 12.335 3505.005 ;
        RECT 12.045 3504.820 13.700 3504.960 ;
        RECT 12.045 3504.775 12.335 3504.820 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3506.300 40.780 3517.600 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 2970.495 10.035 2972.045 ;
      LAYER mcon ;
        RECT 9.805 2971.685 9.975 2971.855 ;
      LAYER met1 ;
        RECT 9.745 2971.840 10.035 2971.885 ;
        RECT 9.745 2971.700 13.700 2971.840 ;
        RECT 9.745 2971.655 10.035 2971.700 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT -4.800 3267.590 13.700 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 3011.955 10.035 3013.505 ;
      LAYER mcon ;
        RECT 9.805 3012.145 9.975 3012.315 ;
      LAYER met1 ;
        RECT 9.730 3012.300 10.050 3012.360 ;
        RECT 9.535 3012.160 10.050 3012.300 ;
        RECT 9.730 3012.100 10.050 3012.160 ;
      LAYER via ;
        RECT 9.760 3012.100 10.020 3012.360 ;
      LAYER met2 ;
        RECT 9.760 3012.070 10.020 3012.390 ;
        RECT 9.820 2980.285 9.960 3012.070 ;
        RECT 9.750 2979.915 10.030 2980.285 ;
      LAYER via2 ;
        RECT 9.750 2979.960 10.030 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 9.725 2980.250 10.055 2980.265 ;
        RECT -4.800 2979.950 10.055 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 9.725 2979.935 10.055 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 2870.515 10.035 2872.065 ;
      LAYER mcon ;
        RECT 9.805 2870.705 9.975 2870.875 ;
      LAYER met1 ;
        RECT 9.745 2870.860 10.035 2870.905 ;
        RECT 9.745 2870.720 13.700 2870.860 ;
        RECT 9.745 2870.675 10.035 2870.720 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT -4.800 2692.990 13.700 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 2500.595 10.035 2502.145 ;
      LAYER mcon ;
        RECT 9.805 2500.785 9.975 2500.955 ;
      LAYER met1 ;
        RECT 9.745 2500.940 10.035 2500.985 ;
        RECT 9.745 2500.800 13.700 2500.940 ;
        RECT 9.745 2500.755 10.035 2500.800 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT -4.800 2405.350 13.700 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1983.795 10.035 1985.345 ;
      LAYER mcon ;
        RECT 9.805 1985.005 9.975 1985.175 ;
      LAYER met1 ;
        RECT 9.745 1985.160 10.035 1985.205 ;
        RECT 9.745 1985.020 13.700 1985.160 ;
        RECT 9.745 1984.975 10.035 1985.020 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT -4.800 2118.390 13.700 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1706.355 10.035 1707.905 ;
      LAYER mcon ;
        RECT 9.805 1707.565 9.975 1707.735 ;
      LAYER met1 ;
        RECT 9.745 1707.720 10.035 1707.765 ;
        RECT 9.745 1707.580 13.700 1707.720 ;
        RECT 9.745 1707.535 10.035 1707.580 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT -4.800 1830.750 13.700 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 734.655 2910.335 736.205 ;
      LAYER mcon ;
        RECT 2910.105 734.825 2910.275 734.995 ;
      LAYER met1 ;
        RECT 2910.045 734.980 2910.335 735.025 ;
        RECT 2906.300 734.840 2910.335 734.980 ;
        RECT 2910.045 734.795 2910.335 734.840 ;
      LAYER met3 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2906.300 674.070 2924.800 674.370 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1581.235 10.035 1582.785 ;
      LAYER mcon ;
        RECT 9.805 1581.425 9.975 1581.595 ;
      LAYER met1 ;
        RECT 9.730 1581.580 10.050 1581.640 ;
        RECT 9.535 1581.440 10.050 1581.580 ;
        RECT 9.730 1581.380 10.050 1581.440 ;
      LAYER via ;
        RECT 9.760 1581.380 10.020 1581.640 ;
      LAYER met2 ;
        RECT 9.760 1581.350 10.020 1581.670 ;
        RECT 9.820 1544.125 9.960 1581.350 ;
        RECT 9.750 1543.755 10.030 1544.125 ;
      LAYER via2 ;
        RECT 9.750 1543.800 10.030 1544.080 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 9.725 1544.090 10.055 1544.105 ;
        RECT -4.800 1543.790 10.055 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 9.725 1543.775 10.055 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1273.215 10.035 1274.765 ;
      LAYER mcon ;
        RECT 9.805 1274.405 9.975 1274.575 ;
      LAYER met1 ;
        RECT 9.730 1274.560 10.050 1274.620 ;
        RECT 9.535 1274.420 10.050 1274.560 ;
        RECT 9.730 1274.360 10.050 1274.420 ;
      LAYER via ;
        RECT 9.760 1274.360 10.020 1274.620 ;
      LAYER met2 ;
        RECT 9.750 1328.195 10.030 1328.565 ;
        RECT 9.820 1274.650 9.960 1328.195 ;
        RECT 9.760 1274.330 10.020 1274.650 ;
      LAYER via2 ;
        RECT 9.750 1328.240 10.030 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 9.725 1328.530 10.055 1328.545 ;
        RECT -4.800 1328.230 10.055 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 9.725 1328.215 10.055 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1033.855 10.035 1035.405 ;
      LAYER mcon ;
        RECT 9.805 1034.705 9.975 1034.875 ;
      LAYER met1 ;
        RECT 9.270 1034.860 9.590 1034.920 ;
        RECT 9.745 1034.860 10.035 1034.905 ;
        RECT 9.270 1034.720 10.035 1034.860 ;
        RECT 9.270 1034.660 9.590 1034.720 ;
        RECT 9.745 1034.675 10.035 1034.720 ;
      LAYER via ;
        RECT 9.300 1034.660 9.560 1034.920 ;
      LAYER met2 ;
        RECT 9.290 1112.635 9.570 1113.005 ;
        RECT 9.360 1034.950 9.500 1112.635 ;
        RECT 9.300 1034.630 9.560 1034.950 ;
      LAYER via2 ;
        RECT 9.290 1112.680 9.570 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 9.265 1112.970 9.595 1112.985 ;
        RECT -4.800 1112.670 9.595 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 9.265 1112.655 9.595 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 629.235 10.035 630.785 ;
      LAYER mcon ;
        RECT 9.805 630.445 9.975 630.615 ;
      LAYER met1 ;
        RECT 9.745 630.600 10.035 630.645 ;
        RECT 9.745 630.460 13.700 630.600 ;
        RECT 9.745 630.415 10.035 630.460 ;
      LAYER met3 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT -4.800 897.110 13.700 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 313.715 10.035 315.265 ;
      LAYER mcon ;
        RECT 9.805 314.925 9.975 315.095 ;
      LAYER met1 ;
        RECT 9.745 315.080 10.035 315.125 ;
        RECT 9.745 314.940 13.700 315.080 ;
        RECT 9.745 314.895 10.035 314.940 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT -4.800 681.550 13.700 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 438.835 10.035 440.385 ;
      LAYER mcon ;
        RECT 9.805 440.045 9.975 440.215 ;
      LAYER met1 ;
        RECT 9.745 440.200 10.035 440.245 ;
        RECT 9.745 440.060 13.700 440.200 ;
        RECT 9.745 440.015 10.035 440.060 ;
      LAYER met3 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT -4.800 465.990 13.700 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 440.895 10.035 442.445 ;
      LAYER mcon ;
        RECT 9.805 441.745 9.975 441.915 ;
      LAYER met1 ;
        RECT 9.745 441.900 10.035 441.945 ;
        RECT 9.745 441.760 13.700 441.900 ;
        RECT 9.745 441.715 10.035 441.760 ;
      LAYER met3 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT -4.800 250.430 13.700 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 391.935 10.035 393.485 ;
      LAYER mcon ;
        RECT 9.805 392.105 9.975 392.275 ;
      LAYER met1 ;
        RECT 9.745 392.260 10.035 392.305 ;
        RECT 9.745 392.120 13.700 392.260 ;
        RECT 9.745 392.075 10.035 392.120 ;
      LAYER met3 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT -4.800 35.550 13.700 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 810.815 2910.335 812.365 ;
      LAYER mcon ;
        RECT 2910.105 812.005 2910.275 812.175 ;
      LAYER met1 ;
        RECT 2910.045 812.160 2910.335 812.205 ;
        RECT 2906.300 812.020 2910.335 812.160 ;
        RECT 2910.045 811.975 2910.335 812.020 ;
      LAYER met3 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2906.300 909.350 2924.800 909.650 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 1006.655 2910.335 1008.205 ;
      LAYER mcon ;
        RECT 2910.105 1007.845 2910.275 1008.015 ;
      LAYER met1 ;
        RECT 2910.045 1008.000 2910.335 1008.045 ;
        RECT 2906.300 1007.860 2910.335 1008.000 ;
        RECT 2910.045 1007.815 2910.335 1007.860 ;
      LAYER met3 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2906.300 1143.950 2924.800 1144.250 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 1265.715 2910.335 1267.265 ;
      LAYER mcon ;
        RECT 2910.105 1266.925 2910.275 1267.095 ;
      LAYER met1 ;
        RECT 2910.045 1267.080 2910.335 1267.125 ;
        RECT 2906.300 1266.940 2910.335 1267.080 ;
        RECT 2910.045 1266.895 2910.335 1266.940 ;
      LAYER met3 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2906.300 1378.550 2924.800 1378.850 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 1670.335 2910.335 1671.885 ;
      LAYER mcon ;
        RECT 2910.105 1670.505 2910.275 1670.675 ;
      LAYER met1 ;
        RECT 2910.045 1670.660 2910.335 1670.705 ;
        RECT 2906.300 1670.520 2910.335 1670.660 ;
        RECT 2910.045 1670.475 2910.335 1670.520 ;
      LAYER met3 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2906.300 1613.150 2924.800 1613.450 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 2116.415 2910.335 2117.965 ;
      LAYER mcon ;
        RECT 2910.105 2116.585 2910.275 2116.755 ;
      LAYER met1 ;
        RECT 2910.045 2116.740 2910.335 2116.785 ;
        RECT 2906.300 2116.600 2910.335 2116.740 ;
        RECT 2910.045 2116.555 2910.335 2116.600 ;
      LAYER met3 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2906.300 1847.750 2924.800 1848.050 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 2263.295 2910.335 2264.845 ;
      LAYER mcon ;
        RECT 2910.105 2263.465 2910.275 2263.635 ;
      LAYER met1 ;
        RECT 2910.045 2263.620 2910.335 2263.665 ;
        RECT 2906.300 2263.480 2910.335 2263.620 ;
        RECT 2910.045 2263.435 2910.335 2263.480 ;
      LAYER met3 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2906.300 2082.350 2924.800 2082.650 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 2386.355 2910.335 2387.905 ;
      LAYER mcon ;
        RECT 2910.105 2386.545 2910.275 2386.715 ;
      LAYER met1 ;
        RECT 2910.045 2386.700 2910.335 2386.745 ;
        RECT 2906.300 2386.560 2910.335 2386.700 ;
        RECT 2910.045 2386.515 2910.335 2386.560 ;
      LAYER met3 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2906.300 2316.950 2924.800 2317.250 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 60.095 2910.335 61.645 ;
      LAYER mcon ;
        RECT 2910.105 61.285 2910.275 61.455 ;
      LAYER met1 ;
        RECT 2910.030 61.440 2910.350 61.500 ;
        RECT 2909.835 61.300 2910.350 61.440 ;
        RECT 2910.030 61.240 2910.350 61.300 ;
      LAYER via ;
        RECT 2910.060 61.240 2910.320 61.500 ;
      LAYER met2 ;
        RECT 2910.050 146.355 2910.330 146.725 ;
        RECT 2910.120 61.530 2910.260 146.355 ;
        RECT 2910.060 61.210 2910.320 61.530 ;
      LAYER via2 ;
        RECT 2910.050 146.400 2910.330 146.680 ;
      LAYER met3 ;
        RECT 2910.025 146.690 2910.355 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2910.025 146.390 2924.800 146.690 ;
        RECT 2910.025 146.375 2910.355 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 2431.935 2910.335 2433.485 ;
      LAYER mcon ;
        RECT 2910.105 2433.125 2910.275 2433.295 ;
      LAYER met1 ;
        RECT 2910.030 2433.280 2910.350 2433.340 ;
        RECT 2909.835 2433.140 2910.350 2433.280 ;
        RECT 2910.030 2433.080 2910.350 2433.140 ;
      LAYER via ;
        RECT 2910.060 2433.080 2910.320 2433.340 ;
      LAYER met2 ;
        RECT 2910.050 2493.035 2910.330 2493.405 ;
        RECT 2910.120 2433.370 2910.260 2493.035 ;
        RECT 2910.060 2433.050 2910.320 2433.370 ;
      LAYER via2 ;
        RECT 2910.050 2493.080 2910.330 2493.360 ;
      LAYER met3 ;
        RECT 2910.025 2493.370 2910.355 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2910.025 2493.070 2924.800 2493.370 ;
        RECT 2910.025 2493.055 2910.355 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 2600.575 2910.335 2602.125 ;
      LAYER mcon ;
        RECT 2910.105 2601.765 2910.275 2601.935 ;
      LAYER met1 ;
        RECT 2910.045 2601.920 2910.335 2601.965 ;
        RECT 2906.300 2601.780 2910.335 2601.920 ;
        RECT 2910.045 2601.735 2910.335 2601.780 ;
      LAYER met3 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2906.300 2727.670 2924.800 2727.970 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2911.195 3365.555 2911.715 3367.105 ;
      LAYER mcon ;
        RECT 2911.485 3365.745 2911.655 3365.915 ;
      LAYER met1 ;
        RECT 2911.425 3365.900 2911.715 3365.945 ;
        RECT 2906.300 3365.760 2911.715 3365.900 ;
        RECT 2911.425 3365.715 2911.715 3365.760 ;
      LAYER met3 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2906.300 2962.270 2924.800 2962.570 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 3400.255 2910.335 3401.805 ;
      LAYER mcon ;
        RECT 2910.105 3400.425 2910.275 3400.595 ;
      LAYER met1 ;
        RECT 2910.045 3400.580 2910.335 3400.625 ;
        RECT 2906.300 3400.440 2910.335 3400.580 ;
        RECT 2910.045 3400.395 2910.335 3400.440 ;
      LAYER met3 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2906.300 3196.870 2924.800 3197.170 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 3503.615 2910.335 3505.165 ;
      LAYER mcon ;
        RECT 2910.105 3503.785 2910.275 3503.955 ;
      LAYER met1 ;
        RECT 2910.045 3503.940 2910.335 3503.985 ;
        RECT 2906.300 3503.800 2910.335 3503.940 ;
        RECT 2910.045 3503.755 2910.335 3503.800 ;
      LAYER met3 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2906.300 3431.470 2924.800 3431.770 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3506.300 2717.520 3517.600 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3506.300 2392.760 3517.600 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3506.300 2068.460 3517.600 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3506.300 1744.160 3517.600 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3506.300 1419.400 3517.600 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2911.195 232.115 2911.715 233.665 ;
      LAYER mcon ;
        RECT 2911.485 233.325 2911.655 233.495 ;
      LAYER met1 ;
        RECT 2911.425 233.480 2911.715 233.525 ;
        RECT 2906.300 233.340 2911.715 233.480 ;
        RECT 2911.425 233.295 2911.715 233.340 ;
      LAYER met3 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2906.300 380.990 2924.800 381.290 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3506.300 1095.100 3517.600 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3517.370 770.800 3517.600 ;
        RECT 770.660 3517.230 772.640 3517.370 ;
        RECT 772.500 3506.300 772.640 3517.230 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3506.300 446.040 3517.600 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 10.435 3503.615 10.955 3505.165 ;
      LAYER mcon ;
        RECT 10.725 3504.125 10.895 3504.295 ;
      LAYER met1 ;
        RECT 10.665 3504.280 10.955 3504.325 ;
        RECT 10.665 3504.140 13.700 3504.280 ;
        RECT 10.665 3504.095 10.955 3504.140 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3506.300 121.740 3517.600 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 3224.115 10.035 3225.665 ;
      LAYER mcon ;
        RECT 9.805 3225.325 9.975 3225.495 ;
      LAYER met1 ;
        RECT 9.745 3225.480 10.035 3225.525 ;
        RECT 9.745 3225.340 13.700 3225.480 ;
        RECT 9.745 3225.295 10.035 3225.340 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT -4.800 3339.670 13.700 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 2954.175 10.035 2955.725 ;
      LAYER mcon ;
        RECT 9.805 2955.365 9.975 2955.535 ;
      LAYER met1 ;
        RECT 9.745 2955.520 10.035 2955.565 ;
        RECT 9.745 2955.380 13.700 2955.520 ;
        RECT 9.745 2955.335 10.035 2955.380 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT -4.800 3052.030 13.700 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 2883.455 10.035 2885.005 ;
      LAYER mcon ;
        RECT 9.805 2884.305 9.975 2884.475 ;
      LAYER met1 ;
        RECT 9.745 2884.460 10.035 2884.505 ;
        RECT 9.745 2884.320 13.700 2884.460 ;
        RECT 9.745 2884.275 10.035 2884.320 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT -4.800 2765.070 13.700 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 2380.915 10.035 2382.465 ;
      LAYER mcon ;
        RECT 9.805 2382.125 9.975 2382.295 ;
      LAYER met1 ;
        RECT 9.745 2382.280 10.035 2382.325 ;
        RECT 9.745 2382.140 13.700 2382.280 ;
        RECT 9.745 2382.095 10.035 2382.140 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT -4.800 2477.430 13.700 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1777.075 10.035 1778.625 ;
      LAYER mcon ;
        RECT 9.805 1778.285 9.975 1778.455 ;
      LAYER met1 ;
        RECT 9.745 1778.440 10.035 1778.485 ;
        RECT 9.745 1778.300 13.700 1778.440 ;
        RECT 9.745 1778.255 10.035 1778.300 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT -4.800 2189.790 13.700 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1953.215 10.035 1954.765 ;
      LAYER mcon ;
        RECT 9.805 1953.385 9.975 1953.555 ;
      LAYER met1 ;
        RECT 9.745 1953.540 10.035 1953.585 ;
        RECT 9.745 1953.400 13.700 1953.540 ;
        RECT 9.745 1953.355 10.035 1953.400 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT -4.800 1902.830 13.700 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2911.195 449.715 2911.715 451.265 ;
      LAYER mcon ;
        RECT 2911.485 450.925 2911.655 451.095 ;
      LAYER met1 ;
        RECT 2911.425 451.080 2911.715 451.125 ;
        RECT 2906.300 450.940 2911.715 451.080 ;
        RECT 2911.425 450.895 2911.715 450.940 ;
      LAYER met3 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2906.300 615.590 2924.800 615.890 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1216.755 10.035 1218.305 ;
      LAYER mcon ;
        RECT 9.805 1217.965 9.975 1218.135 ;
      LAYER met1 ;
        RECT 9.745 1218.120 10.035 1218.165 ;
        RECT 9.745 1217.980 13.700 1218.120 ;
        RECT 9.745 1217.935 10.035 1217.980 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT -4.800 1615.190 13.700 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1327.615 10.035 1329.165 ;
      LAYER mcon ;
        RECT 9.805 1328.805 9.975 1328.975 ;
      LAYER met1 ;
        RECT 9.745 1328.960 10.035 1329.005 ;
        RECT 9.745 1328.820 13.700 1328.960 ;
        RECT 9.745 1328.775 10.035 1328.820 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT -4.800 1400.310 13.700 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1110.015 10.035 1111.565 ;
      LAYER mcon ;
        RECT 9.805 1110.525 9.975 1110.695 ;
      LAYER met1 ;
        RECT 9.730 1110.680 10.050 1110.740 ;
        RECT 9.535 1110.540 10.050 1110.680 ;
        RECT 9.730 1110.480 10.050 1110.540 ;
      LAYER via ;
        RECT 9.760 1110.480 10.020 1110.740 ;
      LAYER met2 ;
        RECT 9.750 1184.715 10.030 1185.085 ;
        RECT 9.820 1110.770 9.960 1184.715 ;
        RECT 9.760 1110.450 10.020 1110.770 ;
      LAYER via2 ;
        RECT 9.750 1184.760 10.030 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 9.725 1185.050 10.055 1185.065 ;
        RECT -4.800 1184.750 10.055 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 9.725 1184.735 10.055 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 1284.095 10.035 1285.645 ;
      LAYER mcon ;
        RECT 9.805 1284.265 9.975 1284.435 ;
      LAYER met1 ;
        RECT 9.745 1284.420 10.035 1284.465 ;
        RECT 9.745 1284.280 13.700 1284.420 ;
        RECT 9.745 1284.235 10.035 1284.280 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT -4.800 969.190 13.700 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 602.035 10.035 603.585 ;
      LAYER mcon ;
        RECT 9.805 603.245 9.975 603.415 ;
      LAYER met1 ;
        RECT 9.745 603.400 10.035 603.445 ;
        RECT 9.745 603.260 13.700 603.400 ;
        RECT 9.745 603.215 10.035 603.260 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT -4.800 753.630 13.700 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 721.715 10.035 723.265 ;
      LAYER mcon ;
        RECT 9.805 721.905 9.975 722.075 ;
      LAYER met1 ;
        RECT 9.745 722.060 10.035 722.105 ;
        RECT 9.745 721.920 13.700 722.060 ;
        RECT 9.745 721.875 10.035 721.920 ;
      LAYER met3 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT -4.800 538.070 13.700 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 10.895 11.135 11.415 12.685 ;
      LAYER mcon ;
        RECT 11.185 12.325 11.355 12.495 ;
      LAYER met1 ;
        RECT 11.125 12.480 11.415 12.525 ;
        RECT 15.710 12.480 16.030 12.540 ;
        RECT 11.125 12.340 16.030 12.480 ;
        RECT 11.125 12.295 11.415 12.340 ;
        RECT 15.710 12.280 16.030 12.340 ;
      LAYER via ;
        RECT 15.740 12.280 16.000 12.540 ;
      LAYER met2 ;
        RECT 15.800 12.570 15.940 13.700 ;
        RECT 15.740 12.250 16.000 12.570 ;
      LAYER met3 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT -4.800 322.510 13.700 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 9.515 400.755 10.035 402.305 ;
      LAYER mcon ;
        RECT 9.805 400.945 9.975 401.115 ;
      LAYER met1 ;
        RECT 9.745 401.100 10.035 401.145 ;
        RECT 9.745 400.960 13.700 401.100 ;
        RECT 9.745 400.915 10.035 400.960 ;
      LAYER met3 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT -4.800 106.950 13.700 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 995.775 2910.335 997.325 ;
      LAYER mcon ;
        RECT 2910.105 995.945 2910.275 996.115 ;
      LAYER met1 ;
        RECT 2910.045 996.100 2910.335 996.145 ;
        RECT 2906.300 995.960 2910.335 996.100 ;
        RECT 2910.045 995.915 2910.335 995.960 ;
      LAYER met3 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2906.300 850.190 2924.800 850.490 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 1300.415 2910.335 1301.965 ;
      LAYER mcon ;
        RECT 2910.105 1300.585 2910.275 1300.755 ;
      LAYER met1 ;
        RECT 2910.045 1300.740 2910.335 1300.785 ;
        RECT 2906.300 1300.600 2910.335 1300.740 ;
        RECT 2910.045 1300.555 2910.335 1300.600 ;
      LAYER met3 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2906.300 1084.790 2924.800 1085.090 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 1526.835 2910.335 1528.385 ;
      LAYER mcon ;
        RECT 2910.105 1527.025 2910.275 1527.195 ;
      LAYER met1 ;
        RECT 2910.045 1527.180 2910.335 1527.225 ;
        RECT 2906.300 1527.040 2910.335 1527.180 ;
        RECT 2910.045 1526.995 2910.335 1527.040 ;
      LAYER met3 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2906.300 1319.390 2924.800 1319.690 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 1472.435 2910.335 1473.985 ;
      LAYER mcon ;
        RECT 2910.105 1473.645 2910.275 1473.815 ;
      LAYER met1 ;
        RECT 2910.045 1473.800 2910.335 1473.845 ;
        RECT 2906.300 1473.660 2910.335 1473.800 ;
        RECT 2910.045 1473.615 2910.335 1473.660 ;
      LAYER met3 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2906.300 1553.990 2924.800 1554.290 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 1515.955 2910.335 1517.505 ;
      LAYER mcon ;
        RECT 2910.105 1517.165 2910.275 1517.335 ;
      LAYER met1 ;
        RECT 2910.045 1517.320 2910.335 1517.365 ;
        RECT 2906.300 1517.180 2910.335 1517.320 ;
        RECT 2910.045 1517.135 2910.335 1517.180 ;
      LAYER met3 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2906.300 1789.270 2924.800 1789.570 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 1934.835 2910.335 1936.385 ;
      LAYER mcon ;
        RECT 2910.105 1936.045 2910.275 1936.215 ;
      LAYER met1 ;
        RECT 2910.030 1936.200 2910.350 1936.260 ;
        RECT 2909.835 1936.060 2910.350 1936.200 ;
        RECT 2910.030 1936.000 2910.350 1936.060 ;
      LAYER via ;
        RECT 2910.060 1936.000 2910.320 1936.260 ;
      LAYER met2 ;
        RECT 2910.050 2023.835 2910.330 2024.205 ;
        RECT 2910.120 1936.290 2910.260 2023.835 ;
        RECT 2910.060 1935.970 2910.320 1936.290 ;
      LAYER via2 ;
        RECT 2910.050 2023.880 2910.330 2024.160 ;
      LAYER met3 ;
        RECT 2910.025 2024.170 2910.355 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2910.025 2023.870 2924.800 2024.170 ;
        RECT 2910.025 2023.855 2910.355 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 2462.515 2910.335 2464.065 ;
      LAYER mcon ;
        RECT 2910.105 2462.705 2910.275 2462.875 ;
      LAYER met1 ;
        RECT 2910.045 2462.860 2910.335 2462.905 ;
        RECT 2906.300 2462.720 2910.335 2462.860 ;
        RECT 2910.045 2462.675 2910.335 2462.720 ;
      LAYER met3 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2906.300 2258.470 2924.800 2258.770 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.460 2.400 2417.600 13.700 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2433.560 9.930 2433.700 13.700 ;
        RECT 2433.560 9.790 2435.080 9.930 ;
        RECT 2434.940 2.400 2435.080 9.790 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.880 2.400 2453.020 13.700 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.820 2.400 2470.960 13.700 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.760 2.400 2488.900 13.700 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.240 2.400 2506.380 13.700 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.720 9.930 2523.860 13.700 ;
        RECT 2523.720 9.790 2524.320 9.930 ;
        RECT 2524.180 2.400 2524.320 9.790 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2542.120 2.400 2542.260 13.700 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2560.060 2.400 2560.200 13.700 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2578.000 2.400 2578.140 13.700 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.480 2.400 2595.620 13.700 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.420 2.400 2613.560 13.700 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.360 2.400 2631.500 13.700 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.300 2.400 2649.440 13.700 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.840 2.400 1774.980 13.700 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.780 2.400 1792.920 13.700 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.720 2.400 1810.860 13.700 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.660 2.400 1828.800 13.700 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1846.140 2.400 1846.280 13.700 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1864.080 2.400 1864.220 13.700 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1882.020 2.400 1882.160 13.700 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.960 2.400 1900.100 13.700 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.900 2.400 1918.040 13.700 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.380 2.400 1935.520 13.700 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.320 2.400 1953.460 13.700 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.260 2.400 1971.400 13.700 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1989.200 2.400 1989.340 13.700 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.680 2.400 2006.820 13.700 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.620 2.400 2024.760 13.700 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.560 2.400 2042.700 13.700 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.500 2.400 2060.640 13.700 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.440 2.400 2078.580 13.700 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.920 2.400 2096.060 13.700 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.860 2.400 2114.000 13.700 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.800 2.400 2131.940 13.700 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.740 2.400 2149.880 13.700 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2167.665 2.805 2167.835 13.700 ;
      LAYER met1 ;
        RECT 2167.590 2.960 2167.910 3.020 ;
        RECT 2167.395 2.820 2167.910 2.960 ;
        RECT 2167.590 2.760 2167.910 2.820 ;
      LAYER via ;
        RECT 2167.620 2.760 2167.880 3.020 ;
      LAYER met2 ;
        RECT 2167.620 2.730 2167.880 3.050 ;
        RECT 2167.680 2.400 2167.820 2.730 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2185.160 2.400 2185.300 13.700 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2203.100 2.400 2203.240 13.700 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2221.040 2.400 2221.180 13.700 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.980 2.400 2239.120 13.700 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2257.380 9.930 2257.520 13.700 ;
        RECT 2256.460 9.790 2257.520 9.930 ;
        RECT 2256.460 2.400 2256.600 9.790 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.400 2.400 2274.540 13.700 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.340 2.400 2292.480 13.700 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.280 2.400 2310.420 13.700 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.220 2.400 2328.360 13.700 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2343.400 9.930 2343.540 13.700 ;
        RECT 2343.400 9.790 2345.840 9.930 ;
        RECT 2345.700 2.400 2345.840 9.790 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.640 2.400 2363.780 13.700 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.580 2.400 2381.720 13.700 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.520 2.400 2399.660 13.700 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 639.100 2.400 639.240 13.700 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.980 2.400 2423.120 13.700 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.920 2.400 2441.060 13.700 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.860 2.400 2459.000 13.700 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.800 2.400 2476.940 13.700 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.740 2.400 2494.880 13.700 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.220 2.400 2512.360 13.700 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2530.160 2.400 2530.300 13.700 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2548.100 2.400 2548.240 13.700 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2566.040 2.400 2566.180 13.700 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.980 2.400 2584.120 13.700 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.580 2.400 817.720 13.700 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.460 2.400 2601.600 13.700 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.400 2.400 2619.540 13.700 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.340 2.400 2637.480 13.700 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.280 2.400 2655.420 13.700 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 11.135 2910.335 12.685 ;
      LAYER mcon ;
        RECT 2910.105 11.305 2910.275 11.475 ;
      LAYER met1 ;
        RECT 2672.670 11.460 2672.990 11.520 ;
        RECT 2910.045 11.460 2910.335 11.505 ;
        RECT 2672.670 11.320 2910.335 11.460 ;
        RECT 2672.670 11.260 2672.990 11.320 ;
        RECT 2910.045 11.275 2910.335 11.320 ;
      LAYER via ;
        RECT 2672.700 11.260 2672.960 11.520 ;
      LAYER met2 ;
        RECT 2672.700 11.230 2672.960 11.550 ;
        RECT 2672.760 2.400 2672.900 11.230 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2911.195 16.575 2911.715 18.125 ;
      LAYER mcon ;
        RECT 2911.485 17.425 2911.655 17.595 ;
      LAYER met1 ;
        RECT 2911.425 17.580 2911.715 17.625 ;
        RECT 2906.300 17.440 2911.715 17.580 ;
        RECT 2911.425 17.395 2911.715 17.440 ;
      LAYER met2 ;
        RECT 2690.700 2.400 2690.840 13.700 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2907.975 14.515 2908.495 16.065 ;
      LAYER mcon ;
        RECT 2908.265 15.725 2908.435 15.895 ;
      LAYER met1 ;
        RECT 2908.205 15.880 2908.495 15.925 ;
        RECT 2906.300 15.740 2908.495 15.880 ;
        RECT 2908.205 15.695 2908.495 15.740 ;
      LAYER met2 ;
        RECT 2708.640 2.400 2708.780 13.700 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.580 2.400 2726.720 13.700 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.520 2.400 2744.660 13.700 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2762.000 2.400 2762.140 13.700 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.520 2.400 835.660 13.700 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.940 2.400 2780.080 13.700 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.880 2.400 2798.020 13.700 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.820 2.400 2815.960 13.700 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.760 2.400 2833.900 13.700 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.815 16.575 2910.335 18.125 ;
      LAYER mcon ;
        RECT 2910.105 16.745 2910.275 16.915 ;
      LAYER met1 ;
        RECT 2910.045 16.900 2910.335 16.945 ;
        RECT 2906.300 16.760 2910.335 16.900 ;
        RECT 2910.045 16.715 2910.335 16.760 ;
      LAYER met2 ;
        RECT 2851.240 2.400 2851.380 13.700 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2909.355 14.515 2909.875 16.065 ;
      LAYER mcon ;
        RECT 2909.645 14.705 2909.815 14.875 ;
      LAYER met1 ;
        RECT 2909.585 14.675 2909.875 14.905 ;
        RECT 2909.660 14.520 2909.800 14.675 ;
        RECT 2906.300 14.380 2909.800 14.520 ;
      LAYER met2 ;
        RECT 2869.180 2.400 2869.320 13.700 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2911.195 14.515 2911.715 16.065 ;
      LAYER mcon ;
        RECT 2911.485 15.045 2911.655 15.215 ;
      LAYER met1 ;
        RECT 2911.425 15.200 2911.715 15.245 ;
        RECT 2906.300 15.060 2911.715 15.200 ;
        RECT 2911.425 15.015 2911.715 15.060 ;
      LAYER met2 ;
        RECT 2887.120 2.400 2887.260 13.700 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2905.060 2.400 2905.200 13.700 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 853.000 2.400 853.140 13.700 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.940 2.400 871.080 13.700 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 889.800 3.130 889.940 13.700 ;
        RECT 888.880 2.990 889.940 3.130 ;
        RECT 888.880 2.400 889.020 2.990 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 907.280 9.930 907.420 13.700 ;
        RECT 906.820 9.790 907.420 9.930 ;
        RECT 906.820 2.400 906.960 9.790 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.300 2.400 924.440 13.700 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.240 2.400 942.380 13.700 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.180 2.400 960.320 13.700 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.120 2.400 978.260 13.700 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.040 2.400 657.180 13.700 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.440 9.930 997.580 13.700 ;
        RECT 996.060 9.790 997.580 9.930 ;
        RECT 996.060 2.400 996.200 9.790 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.540 2.400 1013.680 13.700 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.480 2.400 1031.620 13.700 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.420 2.400 1049.560 13.700 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.360 2.400 1067.500 13.700 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1087.140 8.570 1087.280 13.700 ;
        RECT 1085.300 8.430 1087.280 8.570 ;
        RECT 1085.300 2.400 1085.440 8.430 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.780 2.400 1102.920 13.700 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.720 2.400 1120.860 13.700 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.660 2.400 1138.800 13.700 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.600 2.400 1156.740 13.700 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 674.520 2.400 674.660 13.700 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.620 9.250 1173.760 13.700 ;
        RECT 1173.620 9.110 1174.220 9.250 ;
        RECT 1174.080 2.400 1174.220 9.110 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1191.930 2.960 1192.250 3.020 ;
        RECT 1193.310 2.960 1193.630 3.020 ;
        RECT 1191.930 2.820 1193.630 2.960 ;
        RECT 1191.930 2.760 1192.250 2.820 ;
        RECT 1193.310 2.760 1193.630 2.820 ;
      LAYER via ;
        RECT 1191.960 2.760 1192.220 3.020 ;
        RECT 1193.340 2.760 1193.600 3.020 ;
      LAYER met2 ;
        RECT 1193.400 3.050 1193.540 13.700 ;
        RECT 1191.960 2.730 1192.220 3.050 ;
        RECT 1193.340 2.730 1193.600 3.050 ;
        RECT 1192.020 2.400 1192.160 2.730 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.960 2.400 1210.100 13.700 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.900 2.400 1228.040 13.700 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.840 2.400 1245.980 13.700 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.320 2.400 1263.460 13.700 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.260 2.400 1281.400 13.700 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1300.580 3.130 1300.720 13.700 ;
        RECT 1299.200 2.990 1300.720 3.130 ;
        RECT 1299.200 2.400 1299.340 2.990 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1317.140 2.400 1317.280 13.700 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1335.080 2.400 1335.220 13.700 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.460 2.400 692.600 13.700 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.560 2.400 1352.700 13.700 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.500 2.400 1370.640 13.700 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.440 2.400 1388.580 13.700 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.380 2.400 1406.520 13.700 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.860 2.400 1424.000 13.700 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.800 2.400 1441.940 13.700 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.740 2.400 1459.880 13.700 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.680 2.400 1477.820 13.700 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1496.540 7.890 1496.680 13.700 ;
        RECT 1495.620 7.750 1496.680 7.890 ;
        RECT 1495.620 2.400 1495.760 7.750 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1513.100 2.400 1513.240 13.700 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.400 2.400 710.540 13.700 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1531.040 2.400 1531.180 13.700 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.980 2.400 1549.120 13.700 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.920 2.400 1567.060 13.700 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1577.945 12.665 1578.115 13.700 ;
      LAYER met1 ;
        RECT 1577.885 12.820 1578.175 12.865 ;
        RECT 1584.770 12.820 1585.090 12.880 ;
        RECT 1577.885 12.680 1585.090 12.820 ;
        RECT 1577.885 12.635 1578.175 12.680 ;
        RECT 1584.770 12.620 1585.090 12.680 ;
      LAYER via ;
        RECT 1584.800 12.620 1585.060 12.880 ;
      LAYER met2 ;
        RECT 1584.800 12.590 1585.060 12.910 ;
        RECT 1584.860 2.400 1585.000 12.590 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1577.485 13.005 1577.655 13.700 ;
        RECT 1580.705 13.005 1580.875 13.700 ;
      LAYER met1 ;
        RECT 1577.425 13.160 1577.715 13.205 ;
        RECT 1580.645 13.160 1580.935 13.205 ;
        RECT 1577.425 13.020 1580.935 13.160 ;
        RECT 1577.425 12.975 1577.715 13.020 ;
        RECT 1580.645 12.975 1580.935 13.020 ;
      LAYER met2 ;
        RECT 1602.340 2.400 1602.480 13.700 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1580.245 12.325 1580.415 13.700 ;
      LAYER met1 ;
        RECT 1580.185 12.480 1580.475 12.525 ;
        RECT 1620.190 12.480 1620.510 12.540 ;
        RECT 1580.185 12.340 1620.510 12.480 ;
        RECT 1580.185 12.295 1580.475 12.340 ;
        RECT 1620.190 12.280 1620.510 12.340 ;
      LAYER via ;
        RECT 1620.220 12.280 1620.480 12.540 ;
      LAYER met2 ;
        RECT 1620.220 12.250 1620.480 12.570 ;
        RECT 1620.280 2.400 1620.420 12.250 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1587.605 13.005 1587.775 13.700 ;
        RECT 1603.705 13.005 1603.875 13.700 ;
      LAYER met1 ;
        RECT 1587.545 13.160 1587.835 13.205 ;
        RECT 1603.645 13.160 1603.935 13.205 ;
        RECT 1587.545 13.020 1603.935 13.160 ;
        RECT 1587.545 12.975 1587.835 13.020 ;
        RECT 1603.645 12.975 1603.935 13.020 ;
      LAYER met2 ;
        RECT 1638.220 2.400 1638.360 13.700 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1656.160 2.400 1656.300 13.700 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.640 2.400 1673.780 13.700 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.580 2.400 1691.720 13.700 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.340 2.400 728.480 13.700 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.520 2.400 1709.660 13.700 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.460 2.400 1727.600 13.700 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.400 2.400 1745.540 13.700 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.880 2.400 1763.020 13.700 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.820 2.400 1780.960 13.700 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.760 2.400 1798.900 13.700 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.700 2.400 1816.840 13.700 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.640 2.400 1834.780 13.700 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1852.120 2.400 1852.260 13.700 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1870.060 2.400 1870.200 13.700 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.280 2.400 746.420 13.700 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1888.000 2.400 1888.140 13.700 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.940 2.400 1906.080 13.700 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.420 2.400 1923.560 13.700 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1942.280 7.890 1942.420 13.700 ;
        RECT 1941.360 7.750 1942.420 7.890 ;
        RECT 1941.360 2.400 1941.500 7.750 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.300 2.400 1959.440 13.700 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.240 2.400 1977.380 13.700 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1995.180 2.400 1995.320 13.700 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.660 2.400 2012.800 13.700 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2062.325 13.005 2062.495 13.700 ;
        RECT 2075.665 13.005 2075.835 13.700 ;
      LAYER met1 ;
        RECT 2062.265 13.160 2062.555 13.205 ;
        RECT 2075.605 13.160 2075.895 13.205 ;
        RECT 2062.265 13.020 2075.895 13.160 ;
        RECT 2062.265 12.975 2062.555 13.020 ;
        RECT 2075.605 12.975 2075.895 13.020 ;
      LAYER met2 ;
        RECT 2032.440 6.530 2032.580 13.700 ;
        RECT 2030.600 6.390 2032.580 6.530 ;
        RECT 2030.600 2.400 2030.740 6.390 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.540 2.400 2048.680 13.700 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.600 3.130 765.740 13.700 ;
        RECT 763.760 2.990 765.740 3.130 ;
        RECT 763.760 2.400 763.900 2.990 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.480 2.400 2066.620 13.700 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.420 2.400 2084.560 13.700 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.900 2.400 2102.040 13.700 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2214.125 13.005 2214.295 13.700 ;
        RECT 2227.465 13.005 2227.635 13.700 ;
      LAYER met1 ;
        RECT 2214.065 13.160 2214.355 13.205 ;
        RECT 2227.405 13.160 2227.695 13.205 ;
        RECT 2214.065 13.020 2227.695 13.160 ;
        RECT 2214.065 12.975 2214.355 13.020 ;
        RECT 2227.405 12.975 2227.695 13.020 ;
      LAYER met2 ;
        RECT 2122.140 9.250 2122.280 13.700 ;
        RECT 2119.840 9.110 2122.280 9.250 ;
        RECT 2119.840 2.400 2119.980 9.110 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.780 2.400 2137.920 13.700 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.720 2.400 2155.860 13.700 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.740 13.330 2172.880 13.700 ;
        RECT 2172.740 13.190 2173.340 13.330 ;
        RECT 2173.200 2.400 2173.340 13.190 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2191.140 2.400 2191.280 13.700 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.620 7.210 2208.760 13.700 ;
        RECT 2208.620 7.070 2209.220 7.210 ;
        RECT 2209.080 2.400 2209.220 7.070 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2227.020 2.400 2227.160 13.700 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.700 2.400 781.840 13.700 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.960 2.400 2245.100 13.700 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.440 2.400 2262.580 13.700 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.380 2.400 2280.520 13.700 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.320 2.400 2298.460 13.700 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.260 2.400 2316.400 13.700 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2334.200 2.400 2334.340 13.700 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.680 2.400 2351.820 13.700 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.620 2.400 2369.760 13.700 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.560 2.400 2387.700 13.700 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.500 2.400 2405.640 13.700 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 800.100 3.130 800.240 13.700 ;
        RECT 799.640 2.990 800.240 3.130 ;
        RECT 799.640 2.400 799.780 2.990 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.954000 ;
    PORT
      LAYER li1 ;
        RECT 6.990 126.215 7.340 126.865 ;
        RECT 6.990 41.775 7.340 42.425 ;
        RECT 6.990 17.415 7.340 18.065 ;
        RECT 6.990 14.575 7.340 15.225 ;
        RECT 81.970 11.975 82.320 12.625 ;
        RECT 391.090 11.975 391.440 12.625 ;
      LAYER mcon ;
        RECT 7.045 126.225 7.215 126.395 ;
        RECT 7.045 42.245 7.215 42.415 ;
        RECT 7.045 17.425 7.215 17.595 ;
        RECT 7.045 14.705 7.215 14.875 ;
        RECT 82.025 12.325 82.195 12.495 ;
        RECT 391.145 11.985 391.315 12.155 ;
      LAYER met1 ;
        RECT 7.060 126.580 13.700 126.720 ;
        RECT 7.060 126.440 7.200 126.580 ;
        RECT 6.970 126.380 7.290 126.440 ;
        RECT 6.775 126.240 7.290 126.380 ;
        RECT 6.970 126.180 7.290 126.240 ;
        RECT 6.970 42.400 7.290 42.460 ;
        RECT 6.775 42.260 7.290 42.400 ;
        RECT 6.970 42.200 7.290 42.260 ;
        RECT 6.970 17.580 7.290 17.640 ;
        RECT 6.775 17.440 7.290 17.580 ;
        RECT 6.970 17.380 7.290 17.440 ;
        RECT 6.970 16.900 7.290 16.960 ;
        RECT 6.970 16.760 13.700 16.900 ;
        RECT 6.970 16.700 7.290 16.760 ;
        RECT 2.830 14.860 3.150 14.920 ;
        RECT 6.970 14.860 7.290 14.920 ;
        RECT 2.830 14.720 7.290 14.860 ;
        RECT 2.830 14.660 3.150 14.720 ;
        RECT 6.970 14.660 7.290 14.720 ;
        RECT 81.965 12.480 82.255 12.525 ;
        RECT 82.410 12.480 82.730 12.540 ;
        RECT 81.965 12.340 82.730 12.480 ;
        RECT 81.965 12.295 82.255 12.340 ;
        RECT 82.410 12.280 82.730 12.340 ;
        RECT 390.610 12.140 390.930 12.200 ;
        RECT 391.085 12.140 391.375 12.185 ;
        RECT 395.670 12.140 395.990 12.200 ;
        RECT 390.610 12.000 395.990 12.140 ;
        RECT 390.610 11.940 390.930 12.000 ;
        RECT 391.085 11.955 391.375 12.000 ;
        RECT 395.670 11.940 395.990 12.000 ;
      LAYER via ;
        RECT 7.000 126.180 7.260 126.440 ;
        RECT 7.000 42.200 7.260 42.460 ;
        RECT 7.000 17.380 7.260 17.640 ;
        RECT 7.000 16.700 7.260 16.960 ;
        RECT 2.860 14.660 3.120 14.920 ;
        RECT 7.000 14.660 7.260 14.920 ;
        RECT 82.440 12.280 82.700 12.540 ;
        RECT 390.640 11.940 390.900 12.200 ;
        RECT 395.700 11.940 395.960 12.200 ;
      LAYER met2 ;
        RECT 7.000 126.150 7.260 126.470 ;
        RECT 7.060 42.490 7.200 126.150 ;
        RECT 7.000 42.170 7.260 42.490 ;
        RECT 7.060 17.670 7.200 42.170 ;
        RECT 7.000 17.350 7.260 17.670 ;
        RECT 7.060 16.990 7.200 17.350 ;
        RECT 7.000 16.670 7.260 16.990 ;
        RECT 7.060 14.950 7.200 16.670 ;
        RECT 2.860 14.630 3.120 14.950 ;
        RECT 7.000 14.630 7.260 14.950 ;
        RECT 2.920 2.400 3.060 14.630 ;
        RECT 82.500 12.570 82.640 13.700 ;
        RECT 82.440 12.250 82.700 12.570 ;
        RECT 390.700 12.230 390.840 13.700 ;
        RECT 395.760 12.230 395.900 13.700 ;
        RECT 390.640 11.910 390.900 12.230 ;
        RECT 395.700 12.085 395.960 12.230 ;
        RECT 425.660 12.085 425.800 13.700 ;
        RECT 395.690 11.715 395.970 12.085 ;
        RECT 425.590 11.715 425.870 12.085 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 395.690 11.760 395.970 12.040 ;
        RECT 425.590 11.760 425.870 12.040 ;
      LAYER met3 ;
        RECT 395.665 12.050 395.995 12.065 ;
        RECT 425.565 12.050 425.895 12.065 ;
        RECT 395.665 11.750 425.895 12.050 ;
        RECT 395.665 11.735 395.995 11.750 ;
        RECT 425.565 11.735 425.895 11.750 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 9.360 17.780 13.700 17.920 ;
        RECT 9.360 17.640 9.500 17.780 ;
        RECT 9.270 17.380 9.590 17.640 ;
      LAYER via ;
        RECT 9.300 17.380 9.560 17.640 ;
      LAYER met2 ;
        RECT 9.300 17.350 9.560 17.670 ;
        RECT 9.360 9.250 9.500 17.350 ;
        RECT 8.440 9.110 9.500 9.250 ;
        RECT 8.440 2.400 8.580 9.110 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 88.865 12.870 89.200 13.295 ;
        RECT 89.720 12.870 90.055 13.295 ;
        RECT 88.865 12.700 90.535 12.870 ;
        RECT 8.845 12.275 9.175 12.525 ;
        RECT 12.565 10.285 12.735 12.155 ;
        RECT 90.290 12.135 90.535 12.700 ;
        RECT 88.865 11.965 90.535 12.135 ;
        RECT 58.565 10.285 58.735 11.475 ;
        RECT 88.865 11.205 89.200 11.965 ;
        RECT 89.720 11.205 90.050 11.965 ;
      LAYER mcon ;
        RECT 8.885 12.325 9.055 12.495 ;
        RECT 12.565 11.985 12.735 12.155 ;
        RECT 58.565 11.305 58.735 11.475 ;
        RECT 88.925 11.305 89.095 11.475 ;
      LAYER met1 ;
        RECT 8.825 12.295 9.115 12.525 ;
        RECT 8.900 12.140 9.040 12.295 ;
        RECT 12.505 12.140 12.795 12.185 ;
        RECT 8.900 12.000 12.795 12.140 ;
        RECT 12.505 11.955 12.795 12.000 ;
        RECT 58.505 11.460 58.795 11.505 ;
        RECT 88.865 11.460 89.155 11.505 ;
        RECT 58.505 11.320 89.155 11.460 ;
        RECT 58.505 11.275 58.795 11.320 ;
        RECT 88.865 11.275 89.155 11.320 ;
        RECT 12.505 10.440 12.795 10.485 ;
        RECT 14.330 10.440 14.650 10.500 ;
        RECT 58.505 10.440 58.795 10.485 ;
        RECT 12.505 10.300 58.795 10.440 ;
        RECT 12.505 10.255 12.795 10.300 ;
        RECT 14.330 10.240 14.650 10.300 ;
        RECT 58.505 10.255 58.795 10.300 ;
      LAYER via ;
        RECT 14.360 10.240 14.620 10.500 ;
      LAYER met2 ;
        RECT 14.360 10.210 14.620 10.530 ;
        RECT 14.420 2.400 14.560 10.210 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.400 2.400 20.540 13.700 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.320 2.400 44.460 13.700 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.720 2.400 246.860 13.700 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.200 2.400 264.340 13.700 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.140 2.400 282.280 13.700 ;
        RECT 354.360 13.445 354.500 13.700 ;
        RECT 354.290 13.075 354.570 13.445 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 354.290 13.120 354.570 13.400 ;
      LAYER met3 ;
        RECT 346.230 13.410 346.530 13.700 ;
        RECT 354.265 13.410 354.595 13.425 ;
        RECT 346.230 13.110 354.595 13.410 ;
        RECT 354.265 13.095 354.595 13.110 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.080 2.400 300.220 13.700 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.020 2.400 318.160 13.700 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 205.705 12.155 206.195 12.525 ;
        RECT 207.135 12.355 207.515 12.525 ;
        RECT 207.135 12.155 207.305 12.355 ;
        RECT 204.385 10.285 204.555 12.155 ;
        RECT 205.705 11.985 207.305 12.155 ;
      LAYER mcon ;
        RECT 204.385 11.985 204.555 12.155 ;
        RECT 205.765 11.985 205.935 12.155 ;
      LAYER met1 ;
        RECT 204.325 12.140 204.615 12.185 ;
        RECT 205.705 12.140 205.995 12.185 ;
        RECT 204.325 12.000 205.995 12.140 ;
        RECT 204.325 11.955 204.615 12.000 ;
        RECT 205.705 11.955 205.995 12.000 ;
        RECT 204.325 10.440 204.615 10.485 ;
        RECT 335.870 10.440 336.190 10.500 ;
        RECT 204.325 10.300 336.190 10.440 ;
        RECT 204.325 10.255 204.615 10.300 ;
        RECT 335.870 10.240 336.190 10.300 ;
      LAYER via ;
        RECT 335.900 10.240 336.160 10.500 ;
      LAYER met2 ;
        RECT 335.900 10.210 336.160 10.530 ;
        RECT 335.960 2.400 336.100 10.210 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 351.510 2.960 351.830 3.020 ;
        RECT 353.350 2.960 353.670 3.020 ;
        RECT 351.510 2.820 353.670 2.960 ;
        RECT 351.510 2.760 351.830 2.820 ;
        RECT 353.350 2.760 353.670 2.820 ;
      LAYER via ;
        RECT 351.540 2.760 351.800 3.020 ;
        RECT 353.380 2.760 353.640 3.020 ;
      LAYER met2 ;
        RECT 351.600 3.050 351.740 13.700 ;
        RECT 351.540 2.730 351.800 3.050 ;
        RECT 353.380 2.730 353.640 3.050 ;
        RECT 353.440 2.400 353.580 2.730 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.380 2.400 371.520 13.700 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.320 2.400 389.460 13.700 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.260 2.400 407.400 13.700 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.985 20.485 8.585 20.655 ;
        RECT 6.985 20.115 7.475 20.485 ;
        RECT 8.415 20.315 8.585 20.485 ;
        RECT 8.415 20.285 8.595 20.315 ;
        RECT 8.415 20.115 8.795 20.285 ;
      LAYER mcon ;
        RECT 8.425 20.145 8.595 20.315 ;
      LAYER met1 ;
        RECT 8.365 20.115 8.655 20.345 ;
        RECT 8.440 19.960 8.580 20.115 ;
        RECT 8.440 19.820 13.700 19.960 ;
      LAYER met2 ;
        RECT 68.240 2.400 68.380 13.700 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.740 2.400 424.880 13.700 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.680 2.400 442.820 13.700 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.620 2.400 460.760 13.700 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.560 2.400 478.700 13.700 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.500 2.400 496.640 13.700 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.980 2.400 514.120 13.700 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.920 2.400 532.060 13.700 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.860 2.400 550.000 13.700 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.800 2.400 567.940 13.700 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.740 2.400 585.880 13.700 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 91.610 2.960 91.930 3.020 ;
        RECT 93.450 2.960 93.770 3.020 ;
        RECT 91.610 2.820 93.770 2.960 ;
        RECT 91.610 2.760 91.930 2.820 ;
        RECT 93.450 2.760 93.770 2.820 ;
      LAYER via ;
        RECT 91.640 2.760 91.900 3.020 ;
        RECT 93.480 2.760 93.740 3.020 ;
      LAYER met2 ;
        RECT 93.540 3.050 93.680 13.700 ;
        RECT 91.640 2.730 91.900 3.050 ;
        RECT 93.480 2.730 93.740 3.050 ;
        RECT 91.700 2.400 91.840 2.730 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 603.220 2.400 603.360 13.700 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 621.160 2.400 621.300 13.700 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.620 2.400 115.760 13.700 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.620 12.650 138.760 13.700 ;
        RECT 138.620 12.510 139.680 12.650 ;
        RECT 139.540 2.400 139.680 12.510 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 158.860 13.330 159.000 13.700 ;
        RECT 157.480 13.190 159.000 13.330 ;
        RECT 157.480 2.400 157.620 13.190 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.960 2.400 175.100 13.700 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 192.885 13.005 193.055 13.700 ;
        RECT 203.005 11.985 203.175 13.700 ;
      LAYER met1 ;
        RECT 192.810 13.160 193.130 13.220 ;
        RECT 192.615 13.020 193.130 13.160 ;
        RECT 192.810 12.960 193.130 13.020 ;
        RECT 193.730 12.140 194.050 12.200 ;
        RECT 202.945 12.140 203.235 12.185 ;
        RECT 193.730 12.000 203.235 12.140 ;
        RECT 193.730 11.940 194.050 12.000 ;
        RECT 202.945 11.955 203.235 12.000 ;
      LAYER via ;
        RECT 192.840 12.960 193.100 13.220 ;
        RECT 193.760 11.940 194.020 12.200 ;
      LAYER met2 ;
        RECT 192.840 12.930 193.100 13.250 ;
        RECT 192.900 2.400 193.040 12.930 ;
        RECT 193.820 12.230 193.960 13.700 ;
        RECT 193.760 11.910 194.020 12.230 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.920 7.210 210.060 13.700 ;
        RECT 209.920 7.070 210.980 7.210 ;
        RECT 210.840 2.400 210.980 7.070 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.860 7.210 228.000 13.700 ;
        RECT 227.860 7.070 228.920 7.210 ;
        RECT 228.780 2.400 228.920 7.070 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.460 12.650 48.600 13.700 ;
        RECT 48.460 12.510 50.440 12.650 ;
        RECT 50.300 2.400 50.440 12.510 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 64.470 7.720 64.790 7.780 ;
        RECT 252.610 7.720 252.930 7.780 ;
        RECT 64.470 7.580 252.930 7.720 ;
        RECT 64.470 7.520 64.790 7.580 ;
        RECT 252.610 7.520 252.930 7.580 ;
      LAYER via ;
        RECT 64.500 7.520 64.760 7.780 ;
        RECT 252.640 7.520 252.900 7.780 ;
      LAYER met2 ;
        RECT 64.560 7.810 64.700 13.700 ;
        RECT 252.700 7.810 252.840 13.700 ;
        RECT 64.500 7.490 64.760 7.810 ;
        RECT 252.640 7.490 252.900 7.810 ;
        RECT 252.700 2.400 252.840 7.490 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.180 2.400 270.320 13.700 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 170.730 7.040 171.050 7.100 ;
        RECT 249.850 7.040 250.170 7.100 ;
        RECT 288.030 7.040 288.350 7.100 ;
        RECT 170.730 6.900 288.350 7.040 ;
        RECT 170.730 6.840 171.050 6.900 ;
        RECT 249.850 6.840 250.170 6.900 ;
        RECT 288.030 6.840 288.350 6.900 ;
      LAYER via ;
        RECT 170.760 6.840 171.020 7.100 ;
        RECT 249.880 6.840 250.140 7.100 ;
        RECT 288.060 6.840 288.320 7.100 ;
      LAYER met2 ;
        RECT 170.820 7.130 170.960 13.700 ;
        RECT 249.940 7.130 250.080 13.700 ;
        RECT 170.760 6.810 171.020 7.130 ;
        RECT 249.880 6.810 250.140 7.130 ;
        RECT 288.060 6.810 288.320 7.130 ;
        RECT 288.120 2.400 288.260 6.810 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 138.070 9.420 138.390 9.480 ;
        RECT 305.970 9.420 306.290 9.480 ;
        RECT 138.070 9.280 306.290 9.420 ;
        RECT 138.070 9.220 138.390 9.280 ;
        RECT 305.970 9.220 306.290 9.280 ;
        RECT 305.970 7.380 306.290 7.440 ;
        RECT 310.110 7.380 310.430 7.440 ;
        RECT 305.970 7.240 310.430 7.380 ;
        RECT 305.970 7.180 306.290 7.240 ;
        RECT 310.110 7.180 310.430 7.240 ;
      LAYER via ;
        RECT 138.100 9.220 138.360 9.480 ;
        RECT 306.000 9.220 306.260 9.480 ;
        RECT 306.000 7.180 306.260 7.440 ;
        RECT 310.140 7.180 310.400 7.440 ;
      LAYER met2 ;
        RECT 138.160 9.510 138.300 13.700 ;
        RECT 138.100 9.190 138.360 9.510 ;
        RECT 306.000 9.190 306.260 9.510 ;
        RECT 306.060 7.470 306.200 9.190 ;
        RECT 310.200 7.470 310.340 13.700 ;
        RECT 306.000 7.150 306.260 7.470 ;
        RECT 310.140 7.150 310.400 7.470 ;
        RECT 306.060 2.400 306.200 7.150 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 324.460 13.330 324.600 13.700 ;
        RECT 324.000 13.190 324.600 13.330 ;
        RECT 324.000 2.400 324.140 13.190 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 10.440 341.710 10.500 ;
        RECT 367.610 10.440 367.930 10.500 ;
        RECT 341.390 10.300 367.930 10.440 ;
        RECT 341.390 10.240 341.710 10.300 ;
        RECT 367.610 10.240 367.930 10.300 ;
      LAYER via ;
        RECT 341.420 10.240 341.680 10.500 ;
        RECT 367.640 10.240 367.900 10.500 ;
      LAYER met2 ;
        RECT 341.480 10.530 341.620 13.700 ;
        RECT 367.700 10.530 367.840 13.700 ;
        RECT 341.420 10.210 341.680 10.530 ;
        RECT 367.640 10.210 367.900 10.530 ;
        RECT 341.480 2.400 341.620 10.210 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.240 12.085 91.380 13.700 ;
        RECT 359.420 12.085 359.560 13.700 ;
        RECT 91.170 11.715 91.450 12.085 ;
        RECT 359.350 11.715 359.630 12.085 ;
        RECT 359.420 2.400 359.560 11.715 ;
        RECT 359.210 -4.800 359.770 2.400 ;
      LAYER via2 ;
        RECT 91.170 11.760 91.450 12.040 ;
        RECT 359.350 11.760 359.630 12.040 ;
      LAYER met3 ;
        RECT 91.145 12.050 91.475 12.065 ;
        RECT 359.325 12.050 359.655 12.065 ;
        RECT 91.145 11.750 359.655 12.050 ;
        RECT 91.145 11.735 91.475 11.750 ;
        RECT 359.325 11.735 359.655 11.750 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 267.560 12.325 268.055 12.525 ;
        RECT 285.805 9.945 285.975 12.495 ;
      LAYER mcon ;
        RECT 267.865 12.325 268.035 12.495 ;
        RECT 285.805 12.325 285.975 12.495 ;
      LAYER met1 ;
        RECT 267.805 12.480 268.095 12.525 ;
        RECT 285.745 12.480 286.035 12.525 ;
        RECT 267.805 12.340 286.035 12.480 ;
        RECT 267.805 12.295 268.095 12.340 ;
        RECT 285.745 12.295 286.035 12.340 ;
        RECT 379.110 10.440 379.430 10.500 ;
        RECT 375.060 10.300 379.430 10.440 ;
        RECT 285.745 10.100 286.035 10.145 ;
        RECT 375.060 10.100 375.200 10.300 ;
        RECT 379.110 10.240 379.430 10.300 ;
        RECT 285.745 9.960 375.200 10.100 ;
        RECT 285.745 9.915 286.035 9.960 ;
        RECT 375.060 9.760 375.200 9.960 ;
        RECT 377.270 9.760 377.590 9.820 ;
        RECT 375.060 9.620 377.590 9.760 ;
        RECT 377.270 9.560 377.590 9.620 ;
      LAYER via ;
        RECT 379.140 10.240 379.400 10.500 ;
        RECT 377.300 9.560 377.560 9.820 ;
      LAYER met2 ;
        RECT 379.200 10.530 379.340 13.700 ;
        RECT 379.140 10.210 379.400 10.530 ;
        RECT 377.300 9.530 377.560 9.850 ;
        RECT 377.360 2.400 377.500 9.530 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 6.360 395.530 6.420 ;
        RECT 398.430 6.360 398.750 6.420 ;
        RECT 395.210 6.220 398.750 6.360 ;
        RECT 395.210 6.160 395.530 6.220 ;
        RECT 398.430 6.160 398.750 6.220 ;
      LAYER via ;
        RECT 395.240 6.160 395.500 6.420 ;
        RECT 398.460 6.160 398.720 6.420 ;
      LAYER met2 ;
        RECT 398.520 6.450 398.660 13.700 ;
        RECT 395.240 6.130 395.500 6.450 ;
        RECT 398.460 6.130 398.720 6.450 ;
        RECT 395.300 2.400 395.440 6.130 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 278.905 13.005 279.995 13.175 ;
        RECT 230.300 12.325 230.795 12.525 ;
        RECT 278.905 11.645 279.075 13.005 ;
        RECT 279.825 12.665 279.995 13.005 ;
        RECT 304.205 12.325 307.135 12.495 ;
        RECT 304.205 11.985 304.375 12.325 ;
        RECT 306.965 11.985 307.135 12.325 ;
      LAYER mcon ;
        RECT 230.605 12.325 230.775 12.495 ;
      LAYER met1 ;
        RECT 375.980 13.020 395.900 13.160 ;
        RECT 279.765 12.820 280.055 12.865 ;
        RECT 279.765 12.680 286.420 12.820 ;
        RECT 279.765 12.635 280.055 12.680 ;
        RECT 230.545 12.295 230.835 12.525 ;
        RECT 286.280 12.480 286.420 12.680 ;
        RECT 286.280 12.340 290.100 12.480 ;
        RECT 230.620 11.800 230.760 12.295 ;
        RECT 289.960 12.140 290.100 12.340 ;
        RECT 304.145 12.140 304.435 12.185 ;
        RECT 289.960 12.000 304.435 12.140 ;
        RECT 304.145 11.955 304.435 12.000 ;
        RECT 306.905 12.140 307.195 12.185 ;
        RECT 375.980 12.140 376.120 13.020 ;
        RECT 395.760 12.820 395.900 13.020 ;
        RECT 413.610 12.820 413.930 12.880 ;
        RECT 395.760 12.680 413.930 12.820 ;
        RECT 413.610 12.620 413.930 12.680 ;
        RECT 306.905 12.000 376.120 12.140 ;
        RECT 306.905 11.955 307.195 12.000 ;
        RECT 278.845 11.800 279.135 11.845 ;
        RECT 230.620 11.660 279.135 11.800 ;
        RECT 278.845 11.615 279.135 11.660 ;
      LAYER via ;
        RECT 413.640 12.620 413.900 12.880 ;
      LAYER met2 ;
        RECT 413.700 12.910 413.840 13.700 ;
        RECT 413.640 12.590 413.900 12.910 ;
        RECT 413.700 12.140 413.840 12.590 ;
        RECT 413.240 12.000 413.840 12.140 ;
        RECT 413.240 2.400 413.380 12.000 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 74.130 10.100 74.450 10.160 ;
        RECT 224.090 10.100 224.410 10.160 ;
        RECT 74.130 9.960 224.410 10.100 ;
        RECT 74.130 9.900 74.450 9.960 ;
        RECT 224.090 9.900 224.410 9.960 ;
      LAYER via ;
        RECT 74.160 9.900 74.420 10.160 ;
        RECT 224.120 9.900 224.380 10.160 ;
      LAYER met2 ;
        RECT 224.180 10.190 224.320 13.700 ;
        RECT 74.160 9.870 74.420 10.190 ;
        RECT 224.120 9.870 224.380 10.190 ;
        RECT 74.220 2.400 74.360 9.870 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 455.700 12.325 456.195 12.525 ;
      LAYER mcon ;
        RECT 456.005 12.325 456.175 12.495 ;
      LAYER met1 ;
        RECT 455.930 12.480 456.250 12.540 ;
        RECT 455.735 12.340 456.250 12.480 ;
        RECT 455.930 12.280 456.250 12.340 ;
      LAYER via ;
        RECT 455.960 12.280 456.220 12.540 ;
      LAYER met2 ;
        RECT 430.720 2.400 430.860 13.700 ;
        RECT 456.020 12.570 456.160 13.700 ;
        RECT 455.960 12.250 456.220 12.570 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.660 2.400 448.800 13.700 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 397.985 12.870 398.320 13.295 ;
        RECT 398.840 12.870 399.175 13.295 ;
        RECT 397.985 12.700 399.655 12.870 ;
        RECT 399.410 12.135 399.655 12.700 ;
        RECT 397.985 11.965 399.655 12.135 ;
        RECT 397.985 11.205 398.320 11.965 ;
        RECT 398.840 11.205 399.170 11.965 ;
      LAYER mcon ;
        RECT 399.425 11.985 399.595 12.155 ;
      LAYER met1 ;
        RECT 399.365 12.140 399.655 12.185 ;
        RECT 399.365 12.000 400.960 12.140 ;
        RECT 399.365 11.955 399.655 12.000 ;
        RECT 400.820 11.460 400.960 12.000 ;
        RECT 466.510 11.460 466.830 11.520 ;
        RECT 468.350 11.460 468.670 11.520 ;
        RECT 400.820 11.320 468.670 11.460 ;
        RECT 466.510 11.260 466.830 11.320 ;
        RECT 468.350 11.260 468.670 11.320 ;
      LAYER via ;
        RECT 466.540 11.260 466.800 11.520 ;
        RECT 468.380 11.260 468.640 11.520 ;
      LAYER met2 ;
        RECT 468.440 11.550 468.580 13.700 ;
        RECT 466.540 11.230 466.800 11.550 ;
        RECT 468.380 11.230 468.640 11.550 ;
        RECT 466.600 2.400 466.740 11.230 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.540 2.400 484.680 13.700 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.480 2.400 502.620 13.700 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 519.945 2.805 520.115 13.700 ;
      LAYER met1 ;
        RECT 519.870 2.960 520.190 3.020 ;
        RECT 519.675 2.820 520.190 2.960 ;
        RECT 519.870 2.760 520.190 2.820 ;
      LAYER via ;
        RECT 519.900 2.760 520.160 3.020 ;
      LAYER met2 ;
        RECT 519.900 2.730 520.160 3.050 ;
        RECT 519.960 2.400 520.100 2.730 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.900 2.400 538.040 13.700 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.840 2.400 555.980 13.700 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.780 2.400 573.920 13.700 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.180 12.650 592.320 13.700 ;
        RECT 591.260 12.510 592.320 12.650 ;
        RECT 591.260 2.400 591.400 12.510 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.680 2.400 97.820 13.700 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 609.200 2.400 609.340 13.700 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.140 2.400 627.280 13.700 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.050 13.160 121.370 13.220 ;
        RECT 221.790 13.160 222.110 13.220 ;
        RECT 121.050 13.020 171.880 13.160 ;
        RECT 121.050 12.960 121.370 13.020 ;
        RECT 171.740 12.820 171.880 13.020 ;
        RECT 193.360 13.020 222.110 13.160 ;
        RECT 193.360 12.820 193.500 13.020 ;
        RECT 221.790 12.960 222.110 13.020 ;
        RECT 171.740 12.680 193.500 12.820 ;
      LAYER via ;
        RECT 121.080 12.960 121.340 13.220 ;
        RECT 221.820 12.960 222.080 13.220 ;
      LAYER met2 ;
        RECT 121.140 13.250 121.280 13.700 ;
        RECT 221.880 13.250 222.020 13.700 ;
        RECT 121.080 12.930 121.340 13.250 ;
        RECT 221.820 12.930 222.080 13.250 ;
        RECT 121.140 7.210 121.280 12.930 ;
        RECT 121.140 7.070 121.740 7.210 ;
        RECT 121.600 2.400 121.740 7.070 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 9.760 145.750 9.820 ;
        RECT 331.730 9.760 332.050 9.820 ;
        RECT 145.430 9.620 332.050 9.760 ;
        RECT 145.430 9.560 145.750 9.620 ;
        RECT 331.730 9.560 332.050 9.620 ;
      LAYER via ;
        RECT 145.460 9.560 145.720 9.820 ;
        RECT 331.760 9.560 332.020 9.820 ;
      LAYER met2 ;
        RECT 146.440 10.610 146.580 13.700 ;
        RECT 145.520 10.470 146.580 10.610 ;
        RECT 145.520 9.850 145.660 10.470 ;
        RECT 331.820 9.850 331.960 13.700 ;
        RECT 145.460 9.530 145.720 9.850 ;
        RECT 331.760 9.530 332.020 9.850 ;
        RECT 145.520 2.400 145.660 9.530 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.840 7.210 164.980 13.700 ;
        RECT 163.460 7.070 164.980 7.210 ;
        RECT 163.460 2.400 163.600 7.070 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.940 2.400 181.080 13.700 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.880 2.400 199.020 13.700 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 9.080 217.050 9.140 ;
        RECT 328.510 9.080 328.830 9.140 ;
        RECT 216.730 8.940 328.830 9.080 ;
        RECT 216.730 8.880 217.050 8.940 ;
        RECT 328.510 8.880 328.830 8.940 ;
      LAYER via ;
        RECT 216.760 8.880 217.020 9.140 ;
        RECT 328.540 8.880 328.800 9.140 ;
      LAYER met2 ;
        RECT 216.820 9.170 216.960 13.700 ;
        RECT 328.600 9.170 328.740 13.700 ;
        RECT 216.760 8.850 217.020 9.170 ;
        RECT 328.540 8.850 328.800 9.170 ;
        RECT 216.820 2.400 216.960 8.850 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.760 2.400 234.900 13.700 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.280 2.400 56.420 13.700 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.200 2.400 80.340 13.700 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 116.065 5.525 116.235 13.700 ;
        RECT 151.945 11.985 152.115 13.700 ;
        RECT 171.725 11.985 171.895 13.700 ;
      LAYER met1 ;
        RECT 151.885 12.140 152.175 12.185 ;
        RECT 171.665 12.140 171.955 12.185 ;
        RECT 151.885 12.000 171.955 12.140 ;
        RECT 151.885 11.955 152.175 12.000 ;
        RECT 171.665 11.955 171.955 12.000 ;
        RECT 103.570 5.680 103.890 5.740 ;
        RECT 116.005 5.680 116.295 5.725 ;
        RECT 103.570 5.540 116.295 5.680 ;
        RECT 103.570 5.480 103.890 5.540 ;
        RECT 116.005 5.495 116.295 5.540 ;
      LAYER via ;
        RECT 103.600 5.480 103.860 5.740 ;
      LAYER met2 ;
        RECT 103.600 5.450 103.860 5.770 ;
        RECT 103.660 2.400 103.800 5.450 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 241.645 12.275 242.020 12.605 ;
        RECT 244.865 7.225 245.035 12.495 ;
      LAYER mcon ;
        RECT 241.645 12.325 241.815 12.495 ;
        RECT 244.865 12.325 245.035 12.495 ;
      LAYER met1 ;
        RECT 241.585 12.480 241.875 12.525 ;
        RECT 244.805 12.480 245.095 12.525 ;
        RECT 241.585 12.340 245.095 12.480 ;
        RECT 241.585 12.295 241.875 12.340 ;
        RECT 244.805 12.295 245.095 12.340 ;
        RECT 127.490 7.380 127.810 7.440 ;
        RECT 244.805 7.380 245.095 7.425 ;
        RECT 127.490 7.240 245.095 7.380 ;
        RECT 127.490 7.180 127.810 7.240 ;
        RECT 244.805 7.195 245.095 7.240 ;
      LAYER via ;
        RECT 127.520 7.180 127.780 7.440 ;
      LAYER met2 ;
        RECT 127.520 7.150 127.780 7.470 ;
        RECT 127.580 2.400 127.720 7.150 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.380 2.400 26.520 13.700 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 241.185 12.260 241.475 12.855 ;
      LAYER mcon ;
        RECT 241.185 12.325 241.355 12.495 ;
      LAYER met1 ;
        RECT 227.310 12.820 227.630 12.880 ;
        RECT 227.310 12.680 231.220 12.820 ;
        RECT 227.310 12.620 227.630 12.680 ;
        RECT 231.080 12.140 231.220 12.680 ;
        RECT 241.125 12.295 241.415 12.525 ;
        RECT 241.200 12.140 241.340 12.295 ;
        RECT 231.080 12.000 241.340 12.140 ;
      LAYER via ;
        RECT 227.340 12.620 227.600 12.880 ;
      LAYER met2 ;
        RECT 32.360 2.400 32.500 13.700 ;
        RECT 227.400 12.910 227.540 13.700 ;
        RECT 227.340 12.590 227.600 12.910 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    ANTENNAGATEAREA 834.613953 ;
    ANTENNADIFFAREA 1339.223389 ;
    PORT
      LAYER nwell ;
        RECT 19.590 3507.385 20.430 3508.990 ;
        RECT 33.850 3507.385 34.690 3508.990 ;
        RECT 48.110 3507.385 48.950 3508.990 ;
        RECT 62.370 3507.385 63.210 3508.990 ;
        RECT 76.630 3507.385 77.470 3508.990 ;
        RECT 90.890 3507.385 91.730 3508.990 ;
        RECT 105.150 3507.385 105.990 3508.990 ;
        RECT 119.410 3507.385 120.250 3508.990 ;
        RECT 133.670 3507.385 134.510 3508.990 ;
        RECT 147.930 3507.385 148.770 3508.990 ;
        RECT 162.190 3507.385 163.030 3508.990 ;
        RECT 176.450 3507.385 177.290 3508.990 ;
        RECT 190.710 3507.385 191.550 3508.990 ;
        RECT 204.970 3507.385 205.810 3508.990 ;
        RECT 219.230 3507.385 220.070 3508.990 ;
        RECT 233.490 3507.385 234.330 3508.990 ;
        RECT 247.750 3507.385 248.590 3508.990 ;
        RECT 262.010 3507.385 262.850 3508.990 ;
        RECT 276.270 3507.385 277.110 3508.990 ;
        RECT 290.530 3507.385 291.370 3508.990 ;
        RECT 304.790 3507.385 305.630 3508.990 ;
        RECT 319.050 3507.385 319.890 3508.990 ;
        RECT 333.310 3507.385 334.150 3508.990 ;
        RECT 347.570 3507.385 348.410 3508.990 ;
        RECT 361.830 3507.385 362.670 3508.990 ;
        RECT 376.090 3507.385 376.930 3508.990 ;
        RECT 390.350 3507.385 391.190 3508.990 ;
        RECT 404.610 3507.385 405.450 3508.990 ;
        RECT 418.870 3507.385 419.710 3508.990 ;
        RECT 433.130 3507.385 433.970 3508.990 ;
        RECT 447.390 3507.385 448.230 3508.990 ;
        RECT 461.650 3507.385 462.490 3508.990 ;
        RECT 475.910 3507.385 476.750 3508.990 ;
        RECT 490.170 3507.385 491.010 3508.990 ;
        RECT 504.430 3507.385 505.270 3508.990 ;
        RECT 518.690 3507.385 519.530 3508.990 ;
        RECT 532.950 3507.385 533.790 3508.990 ;
        RECT 547.210 3507.385 548.050 3508.990 ;
        RECT 561.470 3507.385 562.310 3508.990 ;
        RECT 575.730 3507.385 576.570 3508.990 ;
        RECT 589.990 3507.385 590.830 3508.990 ;
        RECT 604.250 3507.385 605.090 3508.990 ;
        RECT 618.510 3507.385 619.350 3508.990 ;
        RECT 632.770 3507.385 633.610 3508.990 ;
        RECT 647.030 3507.385 647.870 3508.990 ;
        RECT 661.290 3507.385 662.130 3508.990 ;
        RECT 675.550 3507.385 676.390 3508.990 ;
        RECT 689.810 3507.385 690.650 3508.990 ;
        RECT 704.070 3507.385 704.910 3508.990 ;
        RECT 718.330 3507.385 719.170 3508.990 ;
        RECT 732.590 3507.385 733.430 3508.990 ;
        RECT 746.850 3507.385 747.690 3508.990 ;
        RECT 761.110 3507.385 761.950 3508.990 ;
        RECT 775.370 3507.385 776.210 3508.990 ;
        RECT 789.630 3507.385 790.470 3508.990 ;
        RECT 803.890 3507.385 804.730 3508.990 ;
        RECT 818.150 3507.385 818.990 3508.990 ;
        RECT 832.410 3507.385 833.250 3508.990 ;
        RECT 846.670 3507.385 847.510 3508.990 ;
        RECT 860.930 3507.385 861.770 3508.990 ;
        RECT 875.190 3507.385 876.030 3508.990 ;
        RECT 889.450 3507.385 890.290 3508.990 ;
        RECT 903.710 3507.385 904.550 3508.990 ;
        RECT 917.970 3507.385 918.810 3508.990 ;
        RECT 932.230 3507.385 933.070 3508.990 ;
        RECT 946.490 3507.385 947.330 3508.990 ;
        RECT 960.750 3507.385 961.590 3508.990 ;
        RECT 975.010 3507.385 975.850 3508.990 ;
        RECT 989.270 3507.385 990.110 3508.990 ;
        RECT 1003.530 3507.385 1004.370 3508.990 ;
        RECT 1017.790 3507.385 1018.630 3508.990 ;
        RECT 1032.050 3507.385 1032.890 3508.990 ;
        RECT 1046.310 3507.385 1047.150 3508.990 ;
        RECT 1060.570 3507.385 1061.410 3508.990 ;
        RECT 1074.830 3507.385 1075.670 3508.990 ;
        RECT 1089.090 3507.385 1089.930 3508.990 ;
        RECT 1103.350 3507.385 1104.190 3508.990 ;
        RECT 1117.610 3507.385 1118.450 3508.990 ;
        RECT 1131.870 3507.385 1132.710 3508.990 ;
        RECT 1146.130 3507.385 1146.970 3508.990 ;
        RECT 1160.390 3507.385 1161.230 3508.990 ;
        RECT 1174.650 3507.385 1175.490 3508.990 ;
        RECT 1188.910 3507.385 1189.750 3508.990 ;
        RECT 1203.170 3507.385 1204.010 3508.990 ;
        RECT 1217.430 3507.385 1218.270 3508.990 ;
        RECT 1231.690 3507.385 1232.530 3508.990 ;
        RECT 1245.950 3507.385 1246.790 3508.990 ;
        RECT 1260.210 3507.385 1261.050 3508.990 ;
        RECT 1274.470 3507.385 1275.310 3508.990 ;
        RECT 1288.730 3507.385 1289.570 3508.990 ;
        RECT 1302.990 3507.385 1303.830 3508.990 ;
        RECT 1317.250 3507.385 1318.090 3508.990 ;
        RECT 1331.510 3507.385 1332.350 3508.990 ;
        RECT 1345.770 3507.385 1346.610 3508.990 ;
        RECT 1360.030 3507.385 1360.870 3508.990 ;
        RECT 1374.290 3507.385 1375.130 3508.990 ;
        RECT 1388.550 3507.385 1389.390 3508.990 ;
        RECT 1402.810 3507.385 1403.650 3508.990 ;
        RECT 1417.070 3507.385 1417.910 3508.990 ;
        RECT 1431.330 3507.385 1432.170 3508.990 ;
        RECT 1445.590 3507.385 1446.430 3508.990 ;
        RECT 1459.850 3507.385 1460.690 3508.990 ;
        RECT 1474.110 3507.385 1474.950 3508.990 ;
        RECT 1488.370 3507.385 1489.210 3508.990 ;
        RECT 1502.630 3507.385 1503.470 3508.990 ;
        RECT 1516.890 3507.385 1517.730 3508.990 ;
        RECT 1531.150 3507.385 1531.990 3508.990 ;
        RECT 1545.410 3507.385 1546.250 3508.990 ;
        RECT 1559.670 3507.385 1560.510 3508.990 ;
        RECT 1573.930 3507.385 1574.770 3508.990 ;
        RECT 1588.190 3507.385 1589.030 3508.990 ;
        RECT 1602.450 3507.385 1603.290 3508.990 ;
        RECT 1616.710 3507.385 1617.550 3508.990 ;
        RECT 1630.970 3507.385 1631.810 3508.990 ;
        RECT 1645.230 3507.385 1646.070 3508.990 ;
        RECT 1659.490 3507.385 1660.330 3508.990 ;
        RECT 1673.750 3507.385 1674.590 3508.990 ;
        RECT 1688.010 3507.385 1688.850 3508.990 ;
        RECT 1702.270 3507.385 1703.110 3508.990 ;
        RECT 1716.530 3507.385 1717.370 3508.990 ;
        RECT 1730.790 3507.385 1731.630 3508.990 ;
        RECT 1745.050 3507.385 1745.890 3508.990 ;
        RECT 1759.310 3507.385 1760.150 3508.990 ;
        RECT 1773.570 3507.385 1774.410 3508.990 ;
        RECT 1787.830 3507.385 1788.670 3508.990 ;
        RECT 1802.090 3507.385 1802.930 3508.990 ;
        RECT 1816.350 3507.385 1817.190 3508.990 ;
        RECT 1830.610 3507.385 1831.450 3508.990 ;
        RECT 1844.870 3507.385 1845.710 3508.990 ;
        RECT 1859.130 3507.385 1859.970 3508.990 ;
        RECT 1873.390 3507.385 1874.230 3508.990 ;
        RECT 1887.650 3507.385 1888.490 3508.990 ;
        RECT 1901.910 3507.385 1902.750 3508.990 ;
        RECT 1916.170 3507.385 1917.010 3508.990 ;
        RECT 1930.430 3507.385 1931.270 3508.990 ;
        RECT 1944.690 3507.385 1945.530 3508.990 ;
        RECT 1958.950 3507.385 1959.790 3508.990 ;
        RECT 1973.210 3507.385 1974.050 3508.990 ;
        RECT 1987.470 3507.385 1988.310 3508.990 ;
        RECT 2001.730 3507.385 2002.570 3508.990 ;
        RECT 2015.990 3507.385 2016.830 3508.990 ;
        RECT 2030.250 3507.385 2031.090 3508.990 ;
        RECT 2044.510 3507.385 2045.350 3508.990 ;
        RECT 2058.770 3507.385 2059.610 3508.990 ;
        RECT 2073.030 3507.385 2073.870 3508.990 ;
        RECT 2087.290 3507.385 2088.130 3508.990 ;
        RECT 2101.550 3507.385 2102.390 3508.990 ;
        RECT 2115.810 3507.385 2116.650 3508.990 ;
        RECT 2130.070 3507.385 2130.910 3508.990 ;
        RECT 2144.330 3507.385 2145.170 3508.990 ;
        RECT 2158.590 3507.385 2159.430 3508.990 ;
        RECT 2172.850 3507.385 2173.690 3508.990 ;
        RECT 2187.110 3507.385 2187.950 3508.990 ;
        RECT 2201.370 3507.385 2202.210 3508.990 ;
        RECT 2215.630 3507.385 2216.470 3508.990 ;
        RECT 2229.890 3507.385 2230.730 3508.990 ;
        RECT 2244.150 3507.385 2244.990 3508.990 ;
        RECT 2258.410 3507.385 2259.250 3508.990 ;
        RECT 2272.670 3507.385 2273.510 3508.990 ;
        RECT 2286.930 3507.385 2287.770 3508.990 ;
        RECT 2301.190 3507.385 2302.030 3508.990 ;
        RECT 2315.450 3507.385 2316.290 3508.990 ;
        RECT 2329.710 3507.385 2330.550 3508.990 ;
        RECT 2343.970 3507.385 2344.810 3508.990 ;
        RECT 2358.230 3507.385 2359.070 3508.990 ;
        RECT 2372.490 3507.385 2373.330 3508.990 ;
        RECT 2386.750 3507.385 2387.590 3508.990 ;
        RECT 2401.010 3507.385 2401.850 3508.990 ;
        RECT 2415.270 3507.385 2416.110 3508.990 ;
        RECT 2429.530 3507.385 2430.370 3508.990 ;
        RECT 2443.790 3507.385 2444.630 3508.990 ;
        RECT 2458.050 3507.385 2458.890 3508.990 ;
        RECT 2472.310 3507.385 2473.150 3508.990 ;
        RECT 2486.570 3507.385 2487.410 3508.990 ;
        RECT 2500.830 3507.385 2501.670 3508.990 ;
        RECT 2515.090 3507.385 2515.930 3508.990 ;
        RECT 2529.350 3507.385 2530.190 3508.990 ;
        RECT 2543.610 3507.385 2544.450 3508.990 ;
        RECT 2557.870 3507.385 2558.710 3508.990 ;
        RECT 2572.130 3507.385 2572.970 3508.990 ;
        RECT 2586.390 3507.385 2587.230 3508.990 ;
        RECT 2600.650 3507.385 2601.490 3508.990 ;
        RECT 2614.910 3507.385 2615.750 3508.990 ;
        RECT 2629.170 3507.385 2630.010 3508.990 ;
        RECT 2643.430 3507.385 2644.270 3508.990 ;
        RECT 2657.690 3507.385 2658.530 3508.990 ;
        RECT 2671.950 3507.385 2672.790 3508.990 ;
        RECT 2686.210 3507.385 2687.050 3508.990 ;
        RECT 2700.470 3507.385 2701.310 3508.990 ;
        RECT 2714.730 3507.385 2715.570 3508.990 ;
        RECT 2728.990 3507.385 2729.830 3508.990 ;
        RECT 2743.250 3507.385 2744.090 3508.990 ;
        RECT 2757.510 3507.385 2758.350 3508.990 ;
        RECT 2771.770 3507.385 2772.610 3508.990 ;
        RECT 2786.030 3507.385 2786.870 3508.990 ;
        RECT 2800.290 3507.385 2801.130 3508.990 ;
        RECT 2814.550 3507.385 2815.390 3508.990 ;
        RECT 2828.810 3507.385 2829.650 3508.990 ;
        RECT 2843.070 3507.385 2843.910 3508.990 ;
        RECT 2857.330 3507.385 2858.170 3508.990 ;
        RECT 2871.590 3507.385 2872.430 3508.990 ;
        RECT 2885.850 3507.385 2886.690 3508.990 ;
        RECT 2900.110 3507.385 2900.950 3508.990 ;
        RECT 2908.850 3503.170 2911.990 3504.775 ;
        RECT 2909.770 3501.945 2910.610 3503.170 ;
        RECT 2909.770 3496.505 2910.610 3498.110 ;
        RECT 2909.770 3491.065 2910.610 3492.670 ;
        RECT 2909.770 3485.625 2910.610 3487.230 ;
        RECT 2909.770 3480.185 2910.610 3481.790 ;
        RECT 2909.770 3474.745 2910.610 3476.350 ;
        RECT 2909.770 3469.305 2910.610 3470.910 ;
        RECT 2909.770 3463.865 2910.610 3465.470 ;
        RECT 2909.770 3458.425 2910.610 3460.030 ;
        RECT 2909.770 3452.985 2910.610 3454.590 ;
        RECT 2909.770 3447.545 2910.610 3449.150 ;
        RECT 2909.770 3442.105 2910.610 3443.710 ;
        RECT 2909.770 3436.665 2910.610 3438.270 ;
        RECT 2909.770 3431.225 2910.610 3432.830 ;
        RECT 2909.770 3425.785 2910.610 3427.390 ;
        RECT 2909.770 3420.345 2910.610 3421.950 ;
        RECT 2909.770 3414.905 2910.610 3416.510 ;
        RECT 2909.770 3409.465 2910.610 3411.070 ;
        RECT 2909.770 3404.025 2910.610 3405.630 ;
        RECT 2908.850 3399.810 2910.610 3401.415 ;
        RECT 2909.770 3398.585 2910.610 3399.810 ;
        RECT 2909.770 3393.145 2910.610 3394.750 ;
        RECT 2909.770 3387.705 2910.610 3389.310 ;
        RECT 2909.770 3382.265 2910.610 3383.870 ;
        RECT 2909.770 3376.825 2910.610 3378.430 ;
        RECT 2909.770 3371.385 2910.610 3372.990 ;
        RECT 2909.770 3365.945 2911.990 3367.550 ;
        RECT 2909.770 3360.505 2910.610 3362.110 ;
        RECT 2909.770 3355.065 2910.610 3356.670 ;
        RECT 2909.770 3349.625 2910.610 3351.230 ;
        RECT 2909.770 3344.185 2910.610 3345.790 ;
        RECT 2909.770 3338.745 2910.610 3340.350 ;
        RECT 2909.770 3333.305 2910.610 3334.910 ;
        RECT 2909.770 3327.865 2910.610 3329.470 ;
        RECT 2909.770 3322.425 2910.610 3324.030 ;
        RECT 2909.770 3316.985 2910.610 3318.590 ;
        RECT 2909.770 3311.545 2910.610 3313.150 ;
        RECT 2909.770 3306.105 2910.610 3307.710 ;
        RECT 2909.770 3300.665 2910.610 3302.270 ;
        RECT 2909.770 3295.225 2910.610 3296.830 ;
        RECT 2909.770 3289.785 2910.610 3291.390 ;
        RECT 2909.770 3284.345 2910.610 3285.950 ;
        RECT 2909.770 3278.905 2910.610 3280.510 ;
        RECT 2909.770 3273.465 2910.610 3275.070 ;
        RECT 2909.770 3268.025 2910.610 3269.630 ;
        RECT 2909.770 3262.585 2910.610 3264.190 ;
        RECT 2909.770 3257.145 2910.610 3258.750 ;
        RECT 2909.770 3251.705 2910.610 3253.310 ;
        RECT 2909.770 3246.265 2910.610 3247.870 ;
        RECT 2909.770 3240.825 2910.610 3242.430 ;
        RECT 2909.770 3235.385 2910.610 3236.990 ;
        RECT 2909.770 3229.945 2910.610 3231.550 ;
        RECT 2909.770 3224.505 2910.610 3226.110 ;
        RECT 2909.770 3219.065 2910.610 3220.670 ;
        RECT 2909.770 3213.625 2910.610 3215.230 ;
        RECT 2909.770 3208.185 2910.610 3209.790 ;
        RECT 2909.770 3202.745 2911.990 3204.350 ;
        RECT 2909.770 3197.305 2910.610 3198.910 ;
        RECT 2909.770 3191.865 2910.610 3193.470 ;
        RECT 2909.770 3186.425 2910.610 3188.030 ;
        RECT 2909.770 3180.985 2910.610 3182.590 ;
        RECT 2909.770 3175.545 2910.610 3177.150 ;
        RECT 2909.770 3170.105 2910.610 3171.710 ;
        RECT 2909.770 3164.665 2910.610 3166.270 ;
        RECT 2909.770 3159.225 2910.610 3160.830 ;
        RECT 2909.770 3153.785 2910.610 3155.390 ;
        RECT 2909.770 3148.345 2910.610 3149.950 ;
        RECT 2909.770 3142.905 2910.610 3144.510 ;
        RECT 2909.770 3137.465 2910.610 3139.070 ;
        RECT 2909.770 3132.025 2910.610 3133.630 ;
        RECT 2909.770 3126.585 2910.610 3128.190 ;
        RECT 2909.770 3121.145 2910.610 3122.750 ;
        RECT 2909.770 3115.705 2910.610 3117.310 ;
        RECT 2909.770 3110.265 2910.610 3111.870 ;
        RECT 2909.770 3104.825 2910.610 3106.430 ;
        RECT 2909.770 3099.385 2910.610 3100.990 ;
        RECT 2908.850 3095.170 2910.610 3096.775 ;
        RECT 2909.770 3093.945 2910.610 3095.170 ;
        RECT 2909.770 3088.505 2910.610 3090.110 ;
        RECT 2909.770 3083.065 2910.610 3084.670 ;
        RECT 2909.770 3077.625 2910.610 3079.230 ;
        RECT 2909.770 3072.185 2910.610 3073.790 ;
        RECT 2909.770 3066.745 2910.610 3068.350 ;
        RECT 2909.770 3061.305 2910.610 3062.910 ;
        RECT 2909.770 3055.865 2910.610 3057.470 ;
        RECT 2909.770 3050.425 2910.610 3052.030 ;
        RECT 2909.770 3044.985 2910.610 3046.590 ;
        RECT 2909.770 3039.545 2910.610 3041.150 ;
        RECT 2909.770 3034.105 2910.610 3035.710 ;
        RECT 2909.770 3028.665 2910.610 3030.270 ;
        RECT 2909.770 3023.225 2910.610 3024.830 ;
        RECT 2909.770 3017.785 2910.610 3019.390 ;
        RECT 2909.770 3012.345 2910.610 3013.950 ;
        RECT 2909.770 3006.905 2910.610 3008.510 ;
        RECT 2909.770 3001.465 2910.610 3003.070 ;
        RECT 2909.770 2996.025 2910.610 2997.630 ;
        RECT 2909.770 2990.585 2910.610 2992.190 ;
        RECT 2909.770 2985.145 2910.610 2986.750 ;
        RECT 2909.770 2979.705 2910.610 2981.310 ;
        RECT 2909.770 2974.265 2910.610 2975.870 ;
        RECT 2909.770 2968.825 2910.610 2970.430 ;
        RECT 2909.770 2963.385 2910.610 2964.990 ;
        RECT 2909.770 2957.945 2910.610 2959.550 ;
        RECT 2909.770 2952.505 2910.610 2954.110 ;
        RECT 2909.770 2947.065 2910.610 2948.670 ;
        RECT 2909.770 2941.625 2910.610 2943.230 ;
        RECT 2909.770 2936.185 2910.610 2937.790 ;
        RECT 2909.770 2930.745 2910.610 2932.350 ;
        RECT 2909.770 2925.305 2910.610 2926.910 ;
        RECT 2909.770 2919.865 2910.610 2921.470 ;
        RECT 2909.770 2914.425 2911.990 2916.030 ;
        RECT 2909.770 2908.985 2910.610 2910.590 ;
        RECT 2909.770 2903.545 2910.610 2905.150 ;
        RECT 2909.770 2898.105 2910.610 2899.710 ;
        RECT 2909.770 2892.665 2910.610 2894.270 ;
        RECT 2909.770 2887.225 2910.610 2888.830 ;
        RECT 2909.770 2881.785 2910.610 2883.390 ;
        RECT 2909.770 2876.345 2910.610 2877.950 ;
        RECT 2909.770 2870.905 2910.610 2872.510 ;
        RECT 2909.770 2865.465 2910.610 2867.070 ;
        RECT 2909.770 2860.025 2910.610 2861.630 ;
        RECT 2909.770 2854.585 2910.610 2856.190 ;
        RECT 2909.770 2849.145 2910.610 2850.750 ;
        RECT 2909.770 2843.705 2910.610 2845.310 ;
        RECT 2909.770 2838.265 2910.610 2839.870 ;
        RECT 2909.770 2832.825 2910.610 2834.430 ;
        RECT 2909.770 2827.385 2910.610 2828.990 ;
        RECT 2909.770 2821.945 2910.610 2823.550 ;
        RECT 2909.770 2816.505 2910.610 2818.110 ;
        RECT 2909.770 2811.065 2910.610 2812.670 ;
        RECT 2909.770 2805.625 2910.610 2807.230 ;
        RECT 2909.770 2800.185 2910.610 2801.790 ;
        RECT 2909.770 2794.745 2910.610 2796.350 ;
        RECT 2909.770 2789.305 2910.610 2790.910 ;
        RECT 2909.770 2783.865 2910.610 2785.470 ;
        RECT 2909.770 2778.425 2910.610 2780.030 ;
        RECT 2908.850 2774.210 2910.610 2775.815 ;
        RECT 2909.770 2772.985 2910.610 2774.210 ;
        RECT 2909.770 2767.545 2910.610 2769.150 ;
        RECT 2909.770 2762.105 2910.610 2763.710 ;
        RECT 2909.770 2756.665 2910.610 2758.270 ;
        RECT 2909.770 2751.225 2910.610 2752.830 ;
        RECT 2909.770 2745.785 2910.610 2747.390 ;
        RECT 2909.770 2740.345 2910.610 2741.950 ;
        RECT 2909.770 2734.905 2910.610 2736.510 ;
        RECT 2909.770 2729.465 2910.610 2731.070 ;
        RECT 2909.770 2724.025 2910.610 2725.630 ;
        RECT 2909.770 2718.585 2910.610 2720.190 ;
        RECT 2909.770 2713.145 2910.610 2714.750 ;
        RECT 2909.770 2707.705 2910.610 2709.310 ;
        RECT 2909.770 2702.265 2910.610 2703.870 ;
        RECT 2909.770 2696.825 2910.610 2698.430 ;
        RECT 2906.300 2687.170 2906.930 2688.775 ;
        RECT 2906.300 2681.730 2906.930 2683.335 ;
        RECT 2906.300 2676.290 2906.930 2677.895 ;
        RECT 2906.300 2670.850 2906.930 2672.455 ;
        RECT 2906.300 2665.410 2906.930 2667.015 ;
        RECT 2906.300 2659.970 2906.930 2661.575 ;
        RECT 2906.300 2654.530 2906.930 2656.135 ;
        RECT 2906.300 2649.090 2906.930 2650.695 ;
        RECT 2906.300 2643.650 2906.930 2645.255 ;
        RECT 2906.300 2638.210 2906.930 2639.815 ;
        RECT 2906.300 2632.770 2906.930 2634.375 ;
        RECT 2906.300 2627.330 2906.930 2628.935 ;
        RECT 2906.300 2621.890 2906.930 2623.495 ;
        RECT 2906.300 2616.450 2906.930 2618.055 ;
        RECT 2906.300 2611.010 2906.930 2612.615 ;
        RECT 2906.300 2605.570 2906.930 2607.175 ;
        RECT 2906.300 2600.130 2906.930 2601.735 ;
        RECT 2906.300 2594.690 2906.930 2596.295 ;
        RECT 2906.300 2589.250 2906.930 2590.855 ;
        RECT 2906.300 2583.810 2906.930 2585.415 ;
        RECT 2906.300 2578.370 2906.930 2579.975 ;
        RECT 2906.300 2572.930 2906.930 2574.535 ;
        RECT 2906.300 2567.490 2906.930 2569.095 ;
        RECT 2906.300 2562.050 2906.930 2563.655 ;
        RECT 2906.300 2556.610 2906.930 2558.215 ;
        RECT 2906.300 2551.170 2906.930 2552.775 ;
        RECT 2906.300 2545.730 2906.930 2547.335 ;
        RECT 2906.300 2540.290 2906.930 2541.895 ;
        RECT 2906.300 2534.850 2906.930 2536.455 ;
        RECT 2906.300 2529.410 2906.930 2531.015 ;
        RECT 2906.300 2523.970 2906.930 2525.575 ;
        RECT 2906.300 2518.530 2906.930 2520.135 ;
        RECT 2906.300 2513.090 2906.930 2514.695 ;
        RECT 2906.300 2507.650 2906.930 2509.255 ;
        RECT 2906.300 2502.210 2906.930 2503.815 ;
        RECT 2906.300 2496.770 2906.930 2498.375 ;
        RECT 2906.300 2491.330 2906.930 2492.935 ;
        RECT 2906.300 2485.890 2906.930 2487.495 ;
        RECT 2906.300 2480.450 2906.930 2482.055 ;
        RECT 2906.300 2475.010 2906.930 2476.615 ;
        RECT 2906.300 2469.570 2906.930 2471.175 ;
        RECT 2906.300 2464.130 2906.930 2465.735 ;
        RECT 2906.300 2458.690 2906.930 2460.295 ;
        RECT 2906.300 2453.250 2906.930 2454.855 ;
        RECT 2906.300 2447.810 2906.930 2449.415 ;
        RECT 2906.300 2442.370 2906.930 2443.975 ;
        RECT 2906.300 2436.930 2906.930 2438.535 ;
        RECT 2906.300 2431.490 2906.930 2433.095 ;
        RECT 2906.300 2426.050 2906.930 2427.655 ;
        RECT 2906.300 2420.610 2906.930 2422.215 ;
        RECT 2906.300 2415.170 2906.930 2416.775 ;
        RECT 2906.300 2409.730 2906.930 2411.335 ;
        RECT 2906.300 2404.290 2906.930 2405.895 ;
        RECT 2906.300 2398.850 2906.930 2400.455 ;
        RECT 2906.300 2393.410 2906.930 2395.015 ;
        RECT 2906.300 2387.970 2906.930 2389.575 ;
        RECT 2906.300 2382.530 2906.930 2384.135 ;
        RECT 2906.300 2377.090 2906.930 2378.695 ;
        RECT 2906.300 2371.650 2906.930 2373.255 ;
        RECT 2906.300 2366.210 2906.930 2367.815 ;
        RECT 2906.300 2360.770 2906.930 2362.375 ;
        RECT 2906.300 2355.330 2906.930 2356.935 ;
        RECT 2906.300 2349.890 2906.930 2351.495 ;
        RECT 2906.300 2344.450 2906.930 2346.055 ;
        RECT 2906.300 2339.010 2906.930 2340.615 ;
        RECT 2906.300 2333.570 2906.930 2335.175 ;
        RECT 2906.300 2328.130 2906.930 2329.735 ;
        RECT 2906.300 2322.690 2906.930 2324.295 ;
        RECT 2906.300 2317.250 2906.930 2318.855 ;
        RECT 2906.300 2311.810 2906.930 2313.415 ;
        RECT 2906.300 2306.370 2906.930 2307.975 ;
        RECT 2906.300 2300.930 2906.930 2302.535 ;
        RECT 2906.300 2295.490 2906.930 2297.095 ;
        RECT 2906.300 2290.050 2906.930 2291.655 ;
        RECT 2906.300 2284.610 2906.930 2286.215 ;
        RECT 2906.300 2279.170 2906.930 2280.775 ;
        RECT 2906.300 2273.730 2906.930 2275.335 ;
        RECT 2906.300 2268.290 2906.930 2269.895 ;
        RECT 2906.300 2262.850 2906.930 2264.455 ;
        RECT 2906.300 2257.410 2906.930 2259.015 ;
        RECT 2906.300 2251.970 2906.930 2253.575 ;
        RECT 2906.300 2246.530 2906.930 2248.135 ;
        RECT 2906.300 2241.090 2906.930 2242.695 ;
        RECT 2906.300 2235.650 2906.930 2237.255 ;
        RECT 2906.300 2230.210 2906.930 2231.815 ;
        RECT 2906.300 2224.770 2906.930 2226.375 ;
        RECT 2906.300 2219.330 2906.930 2220.935 ;
        RECT 2906.300 2213.890 2906.930 2215.495 ;
        RECT 2906.300 2208.450 2906.930 2210.055 ;
        RECT 2906.300 2203.010 2906.930 2204.615 ;
        RECT 2906.300 2197.570 2906.930 2199.175 ;
        RECT 2906.300 2192.130 2906.930 2193.735 ;
        RECT 2906.300 2186.690 2906.930 2188.295 ;
        RECT 2906.300 2181.250 2906.930 2182.855 ;
        RECT 2906.300 2175.810 2906.930 2177.415 ;
        RECT 2906.300 2170.370 2906.930 2171.975 ;
        RECT 2906.300 2164.930 2906.930 2166.535 ;
        RECT 2906.300 2159.490 2906.930 2161.095 ;
        RECT 2906.300 2154.050 2906.930 2155.655 ;
        RECT 2906.300 2148.610 2906.930 2150.215 ;
        RECT 2906.300 2143.170 2906.930 2144.775 ;
        RECT 2906.300 2137.730 2906.930 2139.335 ;
        RECT 2906.300 2132.290 2906.930 2133.895 ;
        RECT 2906.300 2126.850 2906.930 2128.455 ;
        RECT 2906.300 2121.410 2906.930 2123.015 ;
        RECT 2906.300 2115.970 2906.930 2117.575 ;
        RECT 2906.300 2110.530 2906.930 2112.135 ;
        RECT 2906.300 2105.090 2906.930 2106.695 ;
        RECT 2906.300 2099.650 2906.930 2101.255 ;
        RECT 2906.300 2094.210 2906.930 2095.815 ;
        RECT 2906.300 2088.770 2906.930 2090.375 ;
        RECT 2906.300 2083.330 2906.930 2084.935 ;
        RECT 2906.300 2077.890 2906.930 2079.495 ;
        RECT 2906.300 2072.450 2906.930 2074.055 ;
        RECT 2906.300 2067.010 2906.930 2068.615 ;
        RECT 2906.300 2061.570 2906.930 2063.175 ;
        RECT 2906.300 2056.130 2906.930 2057.735 ;
        RECT 2906.300 2050.690 2906.930 2052.295 ;
        RECT 2906.300 2045.250 2906.930 2046.855 ;
        RECT 2906.300 2039.810 2906.930 2041.415 ;
        RECT 2906.300 2034.370 2906.930 2035.975 ;
        RECT 2906.300 2028.930 2906.930 2030.535 ;
        RECT 2906.300 2023.490 2906.930 2025.095 ;
        RECT 2906.300 2018.050 2906.930 2019.655 ;
        RECT 2906.300 2012.610 2906.930 2014.215 ;
        RECT 2906.300 2007.170 2906.930 2008.775 ;
        RECT 2906.300 2001.730 2906.930 2003.335 ;
        RECT 2906.300 1996.290 2906.930 1997.895 ;
        RECT 2906.300 1990.850 2906.930 1992.455 ;
        RECT 2906.300 1985.410 2906.930 1987.015 ;
        RECT 2906.300 1979.970 2906.930 1981.575 ;
        RECT 2906.300 1974.530 2906.930 1976.135 ;
        RECT 2906.300 1969.090 2906.930 1970.695 ;
        RECT 2906.300 1963.650 2906.930 1965.255 ;
        RECT 2906.300 1958.210 2906.930 1959.815 ;
        RECT 2906.300 1952.770 2906.930 1954.375 ;
        RECT 2906.300 1947.330 2906.930 1948.935 ;
        RECT 2906.300 1941.890 2906.930 1943.495 ;
        RECT 2906.300 1936.450 2906.930 1938.055 ;
        RECT 2906.300 1931.010 2906.930 1932.615 ;
        RECT 2906.300 1925.570 2906.930 1927.175 ;
        RECT 2906.300 1920.130 2906.930 1921.735 ;
        RECT 2906.300 1914.690 2906.930 1916.295 ;
        RECT 2906.300 1909.250 2906.930 1910.855 ;
        RECT 2906.300 1903.810 2906.930 1905.415 ;
        RECT 2906.300 1898.370 2906.930 1899.975 ;
        RECT 2906.300 1892.930 2906.930 1894.535 ;
        RECT 2906.300 1887.490 2906.930 1889.095 ;
        RECT 2906.300 1882.050 2906.930 1883.655 ;
        RECT 2906.300 1876.610 2906.930 1878.215 ;
        RECT 2906.300 1871.170 2906.930 1872.775 ;
        RECT 2906.300 1865.730 2906.930 1867.335 ;
        RECT 2906.300 1860.290 2906.930 1861.895 ;
        RECT 2906.300 1854.850 2906.930 1856.455 ;
        RECT 2906.300 1849.410 2906.930 1851.015 ;
        RECT 2906.300 1843.970 2906.930 1845.575 ;
        RECT 2906.300 1838.530 2906.930 1840.135 ;
        RECT 2906.300 1833.090 2906.930 1834.695 ;
        RECT 2906.300 1827.650 2906.930 1829.255 ;
        RECT 2906.300 1822.210 2906.930 1823.815 ;
        RECT 2906.300 1816.770 2906.930 1818.375 ;
        RECT 2906.300 1811.330 2906.930 1812.935 ;
        RECT 2906.300 1805.890 2906.930 1807.495 ;
        RECT 2906.300 1800.450 2906.930 1802.055 ;
        RECT 2906.300 1795.010 2906.930 1796.615 ;
        RECT 2906.300 1789.570 2906.930 1791.175 ;
        RECT 2906.300 1784.130 2906.930 1785.735 ;
        RECT 2906.300 1778.690 2906.930 1780.295 ;
        RECT 2906.300 1773.250 2906.930 1774.855 ;
        RECT 2906.300 1767.810 2906.930 1769.415 ;
        RECT 2906.300 1762.370 2906.930 1763.975 ;
        RECT 2906.300 1756.930 2906.930 1758.535 ;
        RECT 2906.300 1751.490 2906.930 1753.095 ;
        RECT 2906.300 1746.050 2906.930 1747.655 ;
        RECT 2906.300 1740.610 2906.930 1742.215 ;
        RECT 2906.300 1735.170 2906.930 1736.775 ;
        RECT 2906.300 1729.730 2906.930 1731.335 ;
        RECT 2906.300 1724.290 2906.930 1725.895 ;
        RECT 2906.300 1718.850 2906.930 1720.455 ;
        RECT 2906.300 1713.410 2906.930 1715.015 ;
        RECT 2906.300 1707.970 2906.930 1709.575 ;
        RECT 2906.300 1702.530 2906.930 1704.135 ;
        RECT 2906.300 1697.090 2906.930 1698.695 ;
        RECT 2906.300 1691.650 2906.930 1693.255 ;
        RECT 2906.300 1686.210 2906.930 1687.815 ;
        RECT 2906.300 1680.770 2906.930 1682.375 ;
        RECT 2906.300 1675.330 2906.930 1676.935 ;
        RECT 2906.300 1669.890 2906.930 1671.495 ;
        RECT 2906.300 1664.450 2906.930 1666.055 ;
        RECT 2906.300 1659.010 2906.930 1660.615 ;
        RECT 2906.300 1653.570 2906.930 1655.175 ;
        RECT 2906.300 1648.130 2906.930 1649.735 ;
        RECT 2906.300 1642.690 2906.930 1644.295 ;
        RECT 2906.300 1637.250 2906.930 1638.855 ;
        RECT 2906.300 1631.810 2906.930 1633.415 ;
        RECT 2906.300 1626.370 2906.930 1627.975 ;
        RECT 2906.300 1620.930 2906.930 1622.535 ;
        RECT 2906.300 1615.490 2906.930 1617.095 ;
        RECT 2906.300 1610.050 2906.930 1611.655 ;
        RECT 2906.300 1604.610 2906.930 1606.215 ;
        RECT 2906.300 1599.170 2906.930 1600.775 ;
        RECT 2906.300 1593.730 2906.930 1595.335 ;
        RECT 2906.300 1588.290 2906.930 1589.895 ;
        RECT 2906.300 1582.850 2906.930 1584.455 ;
        RECT 2906.300 1577.410 2906.930 1579.015 ;
        RECT 2906.300 1571.970 2906.930 1573.575 ;
        RECT 2906.300 1566.530 2906.930 1568.135 ;
        RECT 2906.300 1561.090 2906.930 1562.695 ;
        RECT 2906.300 1555.650 2906.930 1557.255 ;
        RECT 2906.300 1550.210 2906.930 1551.815 ;
        RECT 2906.300 1544.770 2906.930 1546.375 ;
        RECT 2906.300 1539.330 2906.930 1540.935 ;
        RECT 2906.300 1533.890 2906.930 1535.495 ;
        RECT 2906.300 1528.450 2906.930 1530.055 ;
        RECT 2906.300 1523.010 2906.930 1524.615 ;
        RECT 2906.300 1517.570 2906.930 1519.175 ;
        RECT 2906.300 1512.130 2906.930 1513.735 ;
        RECT 2906.300 1506.690 2906.930 1508.295 ;
        RECT 2906.300 1501.250 2906.930 1502.855 ;
        RECT 2906.300 1495.810 2906.930 1497.415 ;
        RECT 2906.300 1490.370 2906.930 1491.975 ;
        RECT 2906.300 1484.930 2906.930 1486.535 ;
        RECT 2906.300 1479.490 2906.930 1481.095 ;
        RECT 2906.300 1474.050 2906.930 1475.655 ;
        RECT 2906.300 1468.610 2906.930 1470.215 ;
        RECT 2906.300 1463.170 2906.930 1464.775 ;
        RECT 2906.300 1457.730 2906.930 1459.335 ;
        RECT 2906.300 1452.290 2906.930 1453.895 ;
        RECT 2906.300 1446.850 2906.930 1448.455 ;
        RECT 2906.300 1441.410 2906.930 1443.015 ;
        RECT 2906.300 1435.970 2906.930 1437.575 ;
        RECT 2906.300 1430.530 2906.930 1432.135 ;
        RECT 2906.300 1425.090 2906.930 1426.695 ;
        RECT 2906.300 1419.650 2906.930 1421.255 ;
        RECT 2906.300 1414.210 2906.930 1415.815 ;
        RECT 2906.300 1408.770 2906.930 1410.375 ;
        RECT 2906.300 1403.330 2906.930 1404.935 ;
        RECT 2906.300 1397.890 2906.930 1399.495 ;
        RECT 2906.300 1392.450 2906.930 1394.055 ;
        RECT 2906.300 1387.010 2906.930 1388.615 ;
        RECT 2906.300 1381.570 2906.930 1383.175 ;
        RECT 2906.300 1376.130 2906.930 1377.735 ;
        RECT 2906.300 1370.690 2906.930 1372.295 ;
        RECT 2906.300 1365.250 2906.930 1366.855 ;
        RECT 2906.300 1359.810 2906.930 1361.415 ;
        RECT 2906.300 1354.370 2906.930 1355.975 ;
        RECT 2906.300 1348.930 2906.930 1350.535 ;
        RECT 2906.300 1343.490 2906.930 1345.095 ;
        RECT 2906.300 1338.050 2906.930 1339.655 ;
        RECT 2906.300 1332.610 2906.930 1334.215 ;
        RECT 2906.300 1327.170 2906.930 1328.775 ;
        RECT 2906.300 1321.730 2906.930 1323.335 ;
        RECT 2906.300 1316.290 2906.930 1317.895 ;
        RECT 2906.300 1310.850 2906.930 1312.455 ;
        RECT 2906.300 1305.410 2906.930 1307.015 ;
        RECT 2906.300 1299.970 2906.930 1301.575 ;
        RECT 2906.300 1294.530 2906.930 1296.135 ;
        RECT 2906.300 1289.090 2906.930 1290.695 ;
        RECT 2906.300 1283.650 2906.930 1285.255 ;
        RECT 2906.300 1278.210 2906.930 1279.815 ;
        RECT 2906.300 1272.770 2906.930 1274.375 ;
        RECT 2906.300 1267.330 2906.930 1268.935 ;
        RECT 2906.300 1261.890 2906.930 1263.495 ;
        RECT 2906.300 1256.450 2906.930 1258.055 ;
        RECT 2906.300 1251.010 2906.930 1252.615 ;
        RECT 2906.300 1245.570 2906.930 1247.175 ;
        RECT 2909.770 1238.905 2910.610 1240.510 ;
        RECT 2909.770 1233.465 2910.610 1235.070 ;
        RECT 2909.770 1228.025 2910.610 1229.630 ;
        RECT 2909.770 1222.585 2910.610 1224.190 ;
        RECT 2909.770 1217.145 2910.610 1218.750 ;
        RECT 2909.770 1211.705 2910.610 1213.310 ;
        RECT 2909.770 1206.265 2910.610 1207.870 ;
        RECT 2909.770 1200.825 2910.610 1202.430 ;
        RECT 2909.770 1195.385 2910.610 1196.990 ;
        RECT 2909.770 1189.945 2910.610 1191.550 ;
        RECT 2909.770 1184.505 2910.610 1186.110 ;
        RECT 2909.770 1179.065 2910.610 1180.670 ;
        RECT 2909.770 1173.625 2910.610 1175.230 ;
        RECT 2909.770 1168.185 2910.610 1169.790 ;
        RECT 2909.770 1162.745 2910.610 1164.350 ;
        RECT 2909.770 1157.305 2910.610 1158.910 ;
        RECT 2909.770 1151.865 2910.610 1153.470 ;
        RECT 2909.770 1146.425 2910.610 1148.030 ;
        RECT 2909.770 1140.985 2910.610 1142.590 ;
        RECT 2909.770 1135.545 2910.610 1137.150 ;
        RECT 2909.770 1130.105 2910.610 1131.710 ;
        RECT 2909.770 1124.665 2910.610 1126.270 ;
        RECT 2909.770 1119.225 2910.610 1120.830 ;
        RECT 2909.770 1113.785 2910.610 1115.390 ;
        RECT 2909.770 1108.345 2910.610 1109.950 ;
        RECT 2909.770 1102.905 2910.610 1104.510 ;
        RECT 2909.770 1097.465 2910.610 1099.070 ;
        RECT 2909.770 1092.025 2910.610 1093.630 ;
        RECT 2909.770 1086.585 2910.610 1088.190 ;
        RECT 2909.770 1081.145 2910.610 1082.750 ;
        RECT 2909.770 1075.705 2910.610 1077.310 ;
        RECT 2909.770 1070.265 2910.610 1071.870 ;
        RECT 2909.770 1064.825 2910.610 1066.430 ;
        RECT 2909.770 1059.385 2910.610 1060.990 ;
        RECT 2909.770 1053.945 2910.610 1055.550 ;
        RECT 2909.770 1048.505 2910.610 1050.110 ;
        RECT 2909.770 1043.065 2910.610 1044.670 ;
        RECT 2909.770 1037.625 2910.610 1039.230 ;
        RECT 2909.770 1032.185 2910.610 1033.790 ;
        RECT 2909.770 1026.745 2910.610 1028.350 ;
        RECT 2909.770 1021.305 2910.610 1022.910 ;
        RECT 2909.770 1015.865 2910.610 1017.470 ;
        RECT 2909.770 1010.425 2910.610 1012.030 ;
        RECT 2908.850 1006.210 2910.610 1007.815 ;
        RECT 2909.770 1004.985 2910.610 1006.210 ;
        RECT 2909.770 999.545 2910.610 1001.150 ;
        RECT 2908.850 995.330 2910.610 996.935 ;
        RECT 2909.770 994.105 2910.610 995.330 ;
        RECT 2909.770 988.665 2910.610 990.270 ;
        RECT 2909.770 983.225 2910.610 984.830 ;
        RECT 2909.770 977.785 2910.610 979.390 ;
        RECT 2909.770 972.345 2910.610 973.950 ;
        RECT 2909.770 966.905 2910.610 968.510 ;
        RECT 2909.770 961.465 2910.610 963.070 ;
        RECT 2909.770 956.025 2910.610 957.630 ;
        RECT 2909.770 950.585 2910.610 952.190 ;
        RECT 2909.770 945.145 2910.610 946.750 ;
        RECT 2909.770 939.705 2910.610 941.310 ;
        RECT 2909.770 934.265 2910.610 935.870 ;
        RECT 2909.770 928.825 2910.610 930.430 ;
        RECT 2909.770 923.385 2910.610 924.990 ;
        RECT 2909.770 917.945 2910.610 919.550 ;
        RECT 2909.770 912.505 2910.610 914.110 ;
        RECT 2909.770 907.065 2910.610 908.670 ;
        RECT 2909.770 901.625 2910.610 903.230 ;
        RECT 2909.770 896.185 2910.610 897.790 ;
        RECT 2909.770 890.745 2910.610 892.350 ;
        RECT 2909.770 885.305 2910.610 886.910 ;
        RECT 2909.770 879.865 2910.610 881.470 ;
        RECT 2909.770 874.425 2910.610 876.030 ;
        RECT 2909.770 868.985 2910.610 870.590 ;
        RECT 2909.770 863.545 2910.610 865.150 ;
        RECT 2909.770 858.105 2910.610 859.710 ;
        RECT 2909.770 852.665 2910.610 854.270 ;
        RECT 2909.770 847.225 2910.610 848.830 ;
        RECT 2909.770 841.785 2910.610 843.390 ;
        RECT 2909.770 836.345 2910.610 837.950 ;
        RECT 2909.770 830.905 2910.610 832.510 ;
        RECT 2909.770 825.465 2910.610 827.070 ;
        RECT 2909.770 820.025 2910.610 821.630 ;
        RECT 2909.770 814.585 2910.610 816.190 ;
        RECT 2908.850 810.370 2910.610 811.975 ;
        RECT 2909.770 809.145 2910.610 810.370 ;
        RECT 2909.770 803.705 2910.610 805.310 ;
        RECT 2909.770 798.265 2910.610 799.870 ;
        RECT 2909.770 792.825 2910.610 794.430 ;
        RECT 2909.770 787.385 2910.610 788.990 ;
        RECT 2909.770 781.945 2910.610 783.550 ;
        RECT 2909.770 776.505 2910.610 778.110 ;
        RECT 2909.770 771.065 2910.610 772.670 ;
        RECT 2909.770 765.625 2910.610 767.230 ;
        RECT 2909.770 760.185 2910.610 761.790 ;
        RECT 2909.770 754.745 2910.610 756.350 ;
        RECT 2909.770 749.305 2910.610 750.910 ;
        RECT 2909.770 743.865 2910.610 745.470 ;
        RECT 2909.770 738.425 2910.610 740.030 ;
        RECT 2908.850 734.210 2910.610 735.815 ;
        RECT 2909.770 732.985 2910.610 734.210 ;
        RECT 2909.770 727.545 2910.610 729.150 ;
        RECT 2909.770 722.105 2910.610 723.710 ;
        RECT 2909.770 716.665 2910.610 718.270 ;
        RECT 2909.770 711.225 2910.610 712.830 ;
        RECT 2909.770 705.785 2910.610 707.390 ;
        RECT 2909.770 700.345 2910.610 701.950 ;
        RECT 2909.770 694.905 2910.610 696.510 ;
        RECT 2909.770 689.465 2910.610 691.070 ;
        RECT 2909.770 684.025 2910.610 685.630 ;
        RECT 2909.770 678.585 2910.610 680.190 ;
        RECT 2909.770 673.145 2910.610 674.750 ;
        RECT 2909.770 667.705 2910.610 669.310 ;
        RECT 2909.770 662.265 2910.610 663.870 ;
        RECT 2909.770 656.825 2910.610 658.430 ;
        RECT 2909.770 651.385 2910.610 652.990 ;
        RECT 2909.770 645.945 2910.610 647.550 ;
        RECT 2909.770 640.505 2910.610 642.110 ;
        RECT 2909.770 635.065 2910.610 636.670 ;
        RECT 2909.770 629.625 2910.610 631.230 ;
        RECT 2909.770 624.185 2910.610 625.790 ;
        RECT 2909.770 618.745 2910.610 620.350 ;
        RECT 2909.770 613.305 2910.610 614.910 ;
        RECT 2909.770 607.865 2910.610 609.470 ;
        RECT 2909.770 602.425 2910.610 604.030 ;
        RECT 2909.770 596.985 2910.610 598.590 ;
        RECT 2909.770 591.545 2910.610 593.150 ;
        RECT 2909.770 586.105 2910.610 587.710 ;
        RECT 2909.770 580.665 2910.610 582.270 ;
        RECT 2909.770 575.225 2910.610 576.830 ;
        RECT 2909.770 569.785 2910.610 571.390 ;
        RECT 2909.770 564.345 2910.610 565.950 ;
        RECT 2909.770 558.905 2910.610 560.510 ;
        RECT 2909.770 553.465 2910.610 555.070 ;
        RECT 2909.770 548.025 2910.610 549.630 ;
        RECT 2909.770 542.585 2910.610 544.190 ;
        RECT 2909.770 537.145 2910.610 538.750 ;
        RECT 2909.770 531.705 2910.610 533.310 ;
        RECT 2909.770 526.265 2910.610 527.870 ;
        RECT 2909.770 520.825 2910.610 522.430 ;
        RECT 2909.770 515.385 2910.610 516.990 ;
        RECT 2909.770 509.945 2910.610 511.550 ;
        RECT 2909.770 504.505 2910.610 506.110 ;
        RECT 2909.770 499.065 2910.610 500.670 ;
        RECT 2909.770 493.625 2910.610 495.230 ;
        RECT 2909.770 488.185 2910.610 489.790 ;
        RECT 2909.770 482.745 2910.610 484.350 ;
        RECT 2909.770 477.305 2910.610 478.910 ;
        RECT 2909.770 471.865 2910.610 473.470 ;
        RECT 2908.850 467.650 2910.610 469.255 ;
        RECT 2909.770 466.425 2910.610 467.650 ;
        RECT 2909.770 460.985 2910.610 462.590 ;
        RECT 2909.770 455.545 2910.610 457.150 ;
        RECT 2909.770 450.105 2911.990 451.710 ;
        RECT 2909.770 444.665 2910.610 446.270 ;
        RECT 2909.770 439.225 2910.610 440.830 ;
        RECT 2909.770 433.785 2910.610 435.390 ;
        RECT 2909.770 428.345 2910.610 429.950 ;
        RECT 2909.770 422.905 2910.610 424.510 ;
        RECT 2909.770 417.465 2910.610 419.070 ;
        RECT 2909.770 412.025 2910.610 413.630 ;
        RECT 2909.770 406.585 2910.610 408.190 ;
        RECT 2909.770 401.145 2910.610 402.750 ;
        RECT 2909.770 395.705 2910.610 397.310 ;
        RECT 2909.770 390.265 2910.610 391.870 ;
        RECT 2909.770 384.825 2910.610 386.430 ;
        RECT 2909.770 379.385 2910.610 380.990 ;
        RECT 2909.770 373.945 2910.610 375.550 ;
        RECT 2909.770 368.505 2910.610 370.110 ;
        RECT 2909.770 363.065 2910.610 364.670 ;
        RECT 2909.770 357.625 2910.610 359.230 ;
        RECT 2909.770 352.185 2910.610 353.790 ;
        RECT 2909.770 346.745 2910.610 348.350 ;
        RECT 2909.770 341.305 2910.610 342.910 ;
        RECT 2909.770 335.865 2910.610 337.470 ;
        RECT 2909.770 330.425 2910.610 332.030 ;
        RECT 2909.770 324.985 2910.610 326.590 ;
        RECT 2909.770 319.545 2910.610 321.150 ;
        RECT 2909.770 314.105 2910.610 315.710 ;
        RECT 2909.770 308.665 2910.610 310.270 ;
        RECT 2909.770 303.225 2910.610 304.830 ;
        RECT 2909.770 297.785 2910.610 299.390 ;
        RECT 2909.770 292.345 2910.610 293.950 ;
        RECT 2908.850 288.130 2910.610 289.735 ;
        RECT 2909.770 286.905 2910.610 288.130 ;
        RECT 2909.770 281.465 2910.610 283.070 ;
        RECT 2909.770 276.025 2910.610 277.630 ;
        RECT 2909.770 270.585 2910.610 272.190 ;
        RECT 2909.770 265.145 2910.610 266.750 ;
        RECT 2909.770 259.705 2910.610 261.310 ;
        RECT 2909.770 254.265 2910.610 255.870 ;
        RECT 2909.770 248.825 2910.610 250.430 ;
        RECT 2909.770 243.385 2910.610 244.990 ;
        RECT 2909.770 237.945 2910.610 239.550 ;
        RECT 2909.770 232.505 2911.990 234.110 ;
        RECT 2909.770 227.065 2910.610 228.670 ;
        RECT 2909.770 221.625 2910.610 223.230 ;
        RECT 2909.770 216.185 2910.610 217.790 ;
        RECT 2909.770 210.745 2910.610 212.350 ;
        RECT 2909.770 205.305 2910.610 206.910 ;
        RECT 2909.770 199.865 2910.610 201.470 ;
        RECT 2909.770 194.425 2910.610 196.030 ;
        RECT 2909.770 188.985 2910.610 190.590 ;
        RECT 2909.770 183.545 2910.610 185.150 ;
        RECT 2909.770 178.105 2910.610 179.710 ;
        RECT 2909.770 172.665 2910.610 174.270 ;
        RECT 2909.770 167.225 2910.610 168.830 ;
        RECT 2909.770 161.785 2910.610 163.390 ;
        RECT 2909.770 156.345 2910.610 157.950 ;
        RECT 2909.770 150.905 2910.610 152.510 ;
        RECT 2909.770 145.465 2910.610 147.070 ;
        RECT 2909.770 140.025 2910.610 141.630 ;
        RECT 2909.770 134.585 2910.610 136.190 ;
        RECT 2909.770 129.145 2910.610 130.750 ;
        RECT 2909.770 123.705 2910.610 125.310 ;
        RECT 2909.770 118.265 2910.610 119.870 ;
        RECT 2909.770 112.825 2910.610 114.430 ;
        RECT 2909.770 107.385 2910.610 108.990 ;
        RECT 2909.770 101.945 2910.610 103.550 ;
        RECT 2909.770 96.505 2910.610 98.110 ;
        RECT 2909.770 91.065 2910.610 92.670 ;
        RECT 2909.770 85.625 2910.610 87.230 ;
        RECT 2909.770 80.185 2910.610 81.790 ;
        RECT 2909.770 74.745 2910.610 76.350 ;
        RECT 2909.770 69.305 2910.610 70.910 ;
        RECT 2909.770 63.865 2910.610 65.470 ;
        RECT 2908.850 59.650 2910.610 61.255 ;
        RECT 2909.770 58.425 2910.610 59.650 ;
        RECT 2909.770 52.985 2910.610 54.590 ;
        RECT 2909.770 47.545 2910.610 49.150 ;
        RECT 2909.770 42.105 2910.610 43.710 ;
        RECT 2909.770 36.665 2910.610 38.270 ;
        RECT 2909.770 31.225 2910.610 32.830 ;
        RECT 2909.770 25.785 2910.610 27.390 ;
        RECT 2909.770 20.345 2910.610 21.950 ;
        RECT 2908.850 16.510 2911.990 17.735 ;
        RECT 2907.010 14.905 2911.990 16.510 ;
        RECT 19.590 10.690 20.430 12.295 ;
        RECT 33.850 10.690 34.690 12.295 ;
        RECT 48.110 10.690 48.950 12.295 ;
        RECT 62.370 10.690 63.210 12.295 ;
        RECT 76.630 10.690 77.470 12.295 ;
        RECT 90.890 10.690 91.730 12.295 ;
        RECT 105.150 10.690 105.990 12.295 ;
        RECT 119.410 10.690 120.250 12.295 ;
        RECT 133.670 10.690 134.510 12.295 ;
        RECT 147.930 10.690 148.770 12.295 ;
        RECT 162.190 10.690 163.030 12.295 ;
        RECT 176.450 10.690 177.290 12.295 ;
        RECT 190.710 10.690 191.550 12.295 ;
        RECT 204.970 10.690 213.170 12.295 ;
        RECT 219.230 10.690 220.070 12.295 ;
        RECT 233.490 10.690 234.330 12.295 ;
        RECT 247.750 10.690 248.590 12.295 ;
        RECT 262.010 10.690 269.290 12.295 ;
        RECT 276.270 10.690 277.110 12.295 ;
        RECT 290.530 10.690 291.370 12.295 ;
        RECT 304.790 10.690 305.630 12.295 ;
        RECT 319.050 10.690 319.890 12.295 ;
        RECT 333.310 10.690 334.150 12.295 ;
        RECT 347.570 10.690 348.410 12.295 ;
        RECT 361.830 10.690 362.670 12.295 ;
        RECT 376.090 10.690 376.930 12.295 ;
        RECT 390.350 10.690 401.310 12.295 ;
        RECT 404.610 10.690 405.450 12.295 ;
        RECT 418.870 10.690 419.710 12.295 ;
        RECT 433.130 10.690 433.970 12.295 ;
        RECT 447.390 10.690 448.230 12.295 ;
        RECT 461.650 10.690 462.490 12.295 ;
        RECT 475.910 10.690 476.750 12.295 ;
        RECT 490.170 10.690 491.010 12.295 ;
        RECT 504.430 10.690 505.270 12.295 ;
        RECT 518.690 10.690 519.530 12.295 ;
        RECT 532.950 10.690 533.790 12.295 ;
        RECT 547.210 10.690 548.050 12.295 ;
        RECT 561.470 10.690 562.310 12.295 ;
        RECT 575.730 10.690 576.570 12.295 ;
        RECT 589.990 10.690 590.830 12.295 ;
        RECT 604.250 10.690 605.090 12.295 ;
        RECT 618.510 10.690 619.350 12.295 ;
        RECT 632.770 10.690 633.610 12.295 ;
        RECT 647.030 10.690 647.870 12.295 ;
        RECT 661.290 10.690 662.130 12.295 ;
        RECT 675.550 10.690 676.390 12.295 ;
        RECT 689.810 10.690 690.650 12.295 ;
        RECT 704.070 10.690 704.910 12.295 ;
        RECT 718.330 10.690 719.170 12.295 ;
        RECT 732.590 10.690 733.430 12.295 ;
        RECT 746.850 10.690 747.690 12.295 ;
        RECT 761.110 10.690 761.950 12.295 ;
        RECT 775.370 10.690 776.210 12.295 ;
        RECT 789.630 10.690 790.470 12.295 ;
        RECT 803.890 10.690 804.730 12.295 ;
        RECT 818.150 10.690 818.990 12.295 ;
        RECT 832.410 10.690 833.250 12.295 ;
        RECT 846.670 10.690 847.510 12.295 ;
        RECT 860.930 10.690 861.770 12.295 ;
        RECT 875.190 10.690 876.030 12.295 ;
        RECT 889.450 10.690 890.290 12.295 ;
        RECT 903.710 10.690 904.550 12.295 ;
        RECT 917.970 10.690 918.810 12.295 ;
        RECT 932.230 10.690 933.070 12.295 ;
        RECT 946.490 10.690 947.330 12.295 ;
        RECT 960.750 10.690 961.590 12.295 ;
        RECT 975.010 10.690 975.850 12.295 ;
        RECT 989.270 10.690 990.110 12.295 ;
        RECT 1003.530 10.690 1004.370 12.295 ;
        RECT 1017.790 10.690 1018.630 12.295 ;
        RECT 1032.050 10.690 1032.890 12.295 ;
        RECT 1046.310 10.690 1047.150 12.295 ;
        RECT 1060.570 10.690 1061.410 12.295 ;
        RECT 1074.830 10.690 1075.670 12.295 ;
        RECT 1089.090 10.690 1089.930 12.295 ;
        RECT 1103.350 10.690 1104.190 12.295 ;
        RECT 1117.610 10.690 1118.450 12.295 ;
        RECT 1131.870 10.690 1132.710 12.295 ;
        RECT 1146.130 10.690 1146.970 12.295 ;
        RECT 1160.390 10.690 1161.230 12.295 ;
        RECT 1174.650 10.690 1175.490 12.295 ;
        RECT 1188.910 10.690 1189.750 12.295 ;
        RECT 1203.170 10.690 1204.010 12.295 ;
        RECT 1217.430 10.690 1218.270 12.295 ;
        RECT 1231.690 10.690 1232.530 12.295 ;
        RECT 1245.950 10.690 1246.790 12.295 ;
        RECT 1260.210 10.690 1261.050 12.295 ;
        RECT 1274.470 10.690 1275.310 12.295 ;
        RECT 1288.730 10.690 1289.570 12.295 ;
        RECT 1302.990 10.690 1303.830 12.295 ;
        RECT 1317.250 10.690 1318.090 12.295 ;
        RECT 1331.510 10.690 1332.350 12.295 ;
        RECT 1345.770 10.690 1346.610 12.295 ;
        RECT 1360.030 10.690 1360.870 12.295 ;
        RECT 1374.290 10.690 1375.130 12.295 ;
        RECT 1388.550 10.690 1389.390 12.295 ;
        RECT 1402.810 10.690 1403.650 12.295 ;
        RECT 1417.070 10.690 1417.910 12.295 ;
        RECT 1431.330 10.690 1432.170 12.295 ;
        RECT 1445.590 10.690 1446.430 12.295 ;
        RECT 1459.850 10.690 1460.690 12.295 ;
        RECT 1474.110 10.690 1474.950 12.295 ;
        RECT 1488.370 10.690 1489.210 12.295 ;
        RECT 1502.630 10.690 1503.470 12.295 ;
        RECT 1516.890 10.690 1517.730 12.295 ;
        RECT 1531.150 10.690 1531.990 12.295 ;
        RECT 1545.410 10.690 1546.250 12.295 ;
        RECT 1559.670 10.690 1560.510 12.295 ;
        RECT 1573.930 10.690 1574.770 12.295 ;
        RECT 1588.190 10.690 1589.030 12.295 ;
        RECT 1602.450 10.690 1603.290 12.295 ;
        RECT 1616.710 10.690 1617.550 12.295 ;
        RECT 1630.970 10.690 1631.810 12.295 ;
        RECT 1645.230 10.690 1646.070 12.295 ;
        RECT 1659.490 10.690 1660.330 12.295 ;
        RECT 1673.750 10.690 1674.590 12.295 ;
        RECT 1688.010 10.690 1688.850 12.295 ;
        RECT 1702.270 10.690 1703.110 12.295 ;
        RECT 1716.530 10.690 1717.370 12.295 ;
        RECT 1730.790 10.690 1731.630 12.295 ;
        RECT 1745.050 10.690 1745.890 12.295 ;
        RECT 1759.310 10.690 1760.150 12.295 ;
        RECT 1773.570 10.690 1774.410 12.295 ;
        RECT 1787.830 10.690 1788.670 12.295 ;
        RECT 1802.090 10.690 1802.930 12.295 ;
        RECT 1816.350 10.690 1817.190 12.295 ;
        RECT 1830.610 10.690 1831.450 12.295 ;
        RECT 1844.870 10.690 1845.710 12.295 ;
        RECT 1859.130 10.690 1859.970 12.295 ;
        RECT 1873.390 10.690 1874.230 12.295 ;
        RECT 1887.650 10.690 1888.490 12.295 ;
        RECT 1901.910 10.690 1902.750 12.295 ;
        RECT 1916.170 10.690 1917.010 12.295 ;
        RECT 1930.430 10.690 1931.270 12.295 ;
        RECT 1944.690 10.690 1945.530 12.295 ;
        RECT 1958.950 10.690 1959.790 12.295 ;
        RECT 1973.210 10.690 1974.050 12.295 ;
        RECT 1987.470 10.690 1988.310 12.295 ;
        RECT 2001.730 10.690 2002.570 12.295 ;
        RECT 2015.990 10.690 2016.830 12.295 ;
        RECT 2030.250 10.690 2031.090 12.295 ;
        RECT 2044.510 10.690 2045.350 12.295 ;
        RECT 2058.770 10.690 2059.610 12.295 ;
        RECT 2073.030 10.690 2073.870 12.295 ;
        RECT 2087.290 10.690 2088.130 12.295 ;
        RECT 2101.550 10.690 2102.390 12.295 ;
        RECT 2115.810 10.690 2116.650 12.295 ;
        RECT 2130.070 10.690 2130.910 12.295 ;
        RECT 2144.330 10.690 2145.170 12.295 ;
        RECT 2158.590 10.690 2159.430 12.295 ;
        RECT 2172.850 10.690 2173.690 12.295 ;
        RECT 2187.110 10.690 2187.950 12.295 ;
        RECT 2201.370 10.690 2202.210 12.295 ;
        RECT 2215.630 10.690 2216.470 12.295 ;
        RECT 2229.890 10.690 2230.730 12.295 ;
        RECT 2244.150 10.690 2244.990 12.295 ;
        RECT 2258.410 10.690 2259.250 12.295 ;
        RECT 2272.670 10.690 2273.510 12.295 ;
        RECT 2286.930 10.690 2287.770 12.295 ;
        RECT 2301.190 10.690 2302.030 12.295 ;
        RECT 2315.450 10.690 2316.290 12.295 ;
        RECT 2329.710 10.690 2330.550 12.295 ;
        RECT 2343.970 10.690 2344.810 12.295 ;
        RECT 2358.230 10.690 2359.070 12.295 ;
        RECT 2372.490 10.690 2373.330 12.295 ;
        RECT 2386.750 10.690 2387.590 12.295 ;
        RECT 2401.010 10.690 2401.850 12.295 ;
        RECT 2415.270 10.690 2416.110 12.295 ;
        RECT 2429.530 10.690 2430.370 12.295 ;
        RECT 2443.790 10.690 2444.630 12.295 ;
        RECT 2458.050 10.690 2458.890 12.295 ;
        RECT 2472.310 10.690 2473.150 12.295 ;
        RECT 2486.570 10.690 2487.410 12.295 ;
        RECT 2500.830 10.690 2501.670 12.295 ;
        RECT 2515.090 10.690 2515.930 12.295 ;
        RECT 2529.350 10.690 2530.190 12.295 ;
        RECT 2543.610 10.690 2544.450 12.295 ;
        RECT 2557.870 10.690 2558.710 12.295 ;
        RECT 2572.130 10.690 2572.970 12.295 ;
        RECT 2586.390 10.690 2587.230 12.295 ;
        RECT 2600.650 10.690 2601.490 12.295 ;
        RECT 2614.910 10.690 2615.750 12.295 ;
        RECT 2629.170 10.690 2630.010 12.295 ;
        RECT 2643.430 10.690 2644.270 12.295 ;
        RECT 2657.690 10.690 2658.530 12.295 ;
        RECT 2671.950 10.690 2672.790 12.295 ;
        RECT 2686.210 10.690 2687.050 12.295 ;
        RECT 2700.470 10.690 2701.310 12.295 ;
        RECT 2714.730 10.690 2715.570 12.295 ;
        RECT 2728.990 10.690 2729.830 12.295 ;
        RECT 2743.250 10.690 2744.090 12.295 ;
        RECT 2757.510 10.690 2758.350 12.295 ;
        RECT 2771.770 10.690 2772.610 12.295 ;
        RECT 2786.030 10.690 2786.870 12.295 ;
        RECT 2800.290 10.690 2801.130 12.295 ;
        RECT 2814.550 10.690 2815.390 12.295 ;
        RECT 2828.810 10.690 2829.650 12.295 ;
        RECT 2843.070 10.690 2843.910 12.295 ;
        RECT 2857.330 10.690 2858.170 12.295 ;
        RECT 2871.590 10.690 2872.430 12.295 ;
        RECT 2885.850 10.690 2886.690 12.295 ;
        RECT 2900.110 10.690 2900.950 12.295 ;
      LAYER li1 ;
        RECT 5.520 3508.715 6.900 3508.885 ;
        RECT 19.780 3508.715 20.240 3508.885 ;
        RECT 34.040 3508.715 34.500 3508.885 ;
        RECT 48.300 3508.715 48.760 3508.885 ;
        RECT 62.560 3508.715 63.020 3508.885 ;
        RECT 76.820 3508.715 77.280 3508.885 ;
        RECT 91.080 3508.715 91.540 3508.885 ;
        RECT 105.340 3508.715 105.800 3508.885 ;
        RECT 119.600 3508.715 120.060 3508.885 ;
        RECT 133.860 3508.715 134.320 3508.885 ;
        RECT 148.120 3508.715 148.580 3508.885 ;
        RECT 162.380 3508.715 162.840 3508.885 ;
        RECT 176.640 3508.715 177.100 3508.885 ;
        RECT 190.900 3508.715 191.360 3508.885 ;
        RECT 205.160 3508.715 205.620 3508.885 ;
        RECT 219.420 3508.715 219.880 3508.885 ;
        RECT 233.680 3508.715 234.140 3508.885 ;
        RECT 247.940 3508.715 248.400 3508.885 ;
        RECT 262.200 3508.715 262.660 3508.885 ;
        RECT 276.460 3508.715 276.920 3508.885 ;
        RECT 290.720 3508.715 291.180 3508.885 ;
        RECT 304.980 3508.715 305.440 3508.885 ;
        RECT 319.240 3508.715 319.700 3508.885 ;
        RECT 333.500 3508.715 333.960 3508.885 ;
        RECT 347.760 3508.715 348.220 3508.885 ;
        RECT 362.020 3508.715 362.480 3508.885 ;
        RECT 376.280 3508.715 376.740 3508.885 ;
        RECT 390.540 3508.715 391.000 3508.885 ;
        RECT 404.800 3508.715 405.260 3508.885 ;
        RECT 419.060 3508.715 419.520 3508.885 ;
        RECT 433.320 3508.715 433.780 3508.885 ;
        RECT 447.580 3508.715 448.040 3508.885 ;
        RECT 461.840 3508.715 462.300 3508.885 ;
        RECT 476.100 3508.715 476.560 3508.885 ;
        RECT 490.360 3508.715 490.820 3508.885 ;
        RECT 504.620 3508.715 505.080 3508.885 ;
        RECT 518.880 3508.715 519.340 3508.885 ;
        RECT 533.140 3508.715 533.600 3508.885 ;
        RECT 547.400 3508.715 547.860 3508.885 ;
        RECT 561.660 3508.715 562.120 3508.885 ;
        RECT 575.920 3508.715 576.380 3508.885 ;
        RECT 590.180 3508.715 590.640 3508.885 ;
        RECT 604.440 3508.715 604.900 3508.885 ;
        RECT 618.700 3508.715 619.160 3508.885 ;
        RECT 632.960 3508.715 633.420 3508.885 ;
        RECT 647.220 3508.715 647.680 3508.885 ;
        RECT 661.480 3508.715 661.940 3508.885 ;
        RECT 675.740 3508.715 676.200 3508.885 ;
        RECT 690.000 3508.715 690.460 3508.885 ;
        RECT 704.260 3508.715 704.720 3508.885 ;
        RECT 718.520 3508.715 718.980 3508.885 ;
        RECT 732.780 3508.715 733.240 3508.885 ;
        RECT 747.040 3508.715 747.500 3508.885 ;
        RECT 761.300 3508.715 761.760 3508.885 ;
        RECT 775.560 3508.715 776.020 3508.885 ;
        RECT 789.820 3508.715 790.280 3508.885 ;
        RECT 804.080 3508.715 804.540 3508.885 ;
        RECT 818.340 3508.715 818.800 3508.885 ;
        RECT 832.600 3508.715 833.060 3508.885 ;
        RECT 846.860 3508.715 847.320 3508.885 ;
        RECT 861.120 3508.715 861.580 3508.885 ;
        RECT 875.380 3508.715 875.840 3508.885 ;
        RECT 889.640 3508.715 890.100 3508.885 ;
        RECT 903.900 3508.715 904.360 3508.885 ;
        RECT 918.160 3508.715 918.620 3508.885 ;
        RECT 932.420 3508.715 932.880 3508.885 ;
        RECT 946.680 3508.715 947.140 3508.885 ;
        RECT 960.940 3508.715 961.400 3508.885 ;
        RECT 975.200 3508.715 975.660 3508.885 ;
        RECT 989.460 3508.715 989.920 3508.885 ;
        RECT 1003.720 3508.715 1004.180 3508.885 ;
        RECT 1017.980 3508.715 1018.440 3508.885 ;
        RECT 1032.240 3508.715 1032.700 3508.885 ;
        RECT 1046.500 3508.715 1046.960 3508.885 ;
        RECT 1060.760 3508.715 1061.220 3508.885 ;
        RECT 1075.020 3508.715 1075.480 3508.885 ;
        RECT 1089.280 3508.715 1089.740 3508.885 ;
        RECT 1103.540 3508.715 1104.000 3508.885 ;
        RECT 1117.800 3508.715 1118.260 3508.885 ;
        RECT 1132.060 3508.715 1132.520 3508.885 ;
        RECT 1146.320 3508.715 1146.780 3508.885 ;
        RECT 1160.580 3508.715 1161.040 3508.885 ;
        RECT 1174.840 3508.715 1175.300 3508.885 ;
        RECT 1189.100 3508.715 1189.560 3508.885 ;
        RECT 1203.360 3508.715 1203.820 3508.885 ;
        RECT 1217.620 3508.715 1218.080 3508.885 ;
        RECT 1231.880 3508.715 1232.340 3508.885 ;
        RECT 1246.140 3508.715 1246.600 3508.885 ;
        RECT 1260.400 3508.715 1260.860 3508.885 ;
        RECT 1274.660 3508.715 1275.120 3508.885 ;
        RECT 1288.920 3508.715 1289.380 3508.885 ;
        RECT 1303.180 3508.715 1303.640 3508.885 ;
        RECT 1317.440 3508.715 1317.900 3508.885 ;
        RECT 1331.700 3508.715 1332.160 3508.885 ;
        RECT 1345.960 3508.715 1346.420 3508.885 ;
        RECT 1360.220 3508.715 1360.680 3508.885 ;
        RECT 1374.480 3508.715 1374.940 3508.885 ;
        RECT 1388.740 3508.715 1389.200 3508.885 ;
        RECT 1403.000 3508.715 1403.460 3508.885 ;
        RECT 1417.260 3508.715 1417.720 3508.885 ;
        RECT 1431.520 3508.715 1431.980 3508.885 ;
        RECT 1445.780 3508.715 1446.240 3508.885 ;
        RECT 1460.040 3508.715 1460.500 3508.885 ;
        RECT 1474.300 3508.715 1474.760 3508.885 ;
        RECT 1488.560 3508.715 1489.020 3508.885 ;
        RECT 1502.820 3508.715 1503.280 3508.885 ;
        RECT 1517.080 3508.715 1517.540 3508.885 ;
        RECT 1531.340 3508.715 1531.800 3508.885 ;
        RECT 1545.600 3508.715 1546.060 3508.885 ;
        RECT 1559.860 3508.715 1560.320 3508.885 ;
        RECT 1574.120 3508.715 1574.580 3508.885 ;
        RECT 1588.380 3508.715 1588.840 3508.885 ;
        RECT 1602.640 3508.715 1603.100 3508.885 ;
        RECT 1616.900 3508.715 1617.360 3508.885 ;
        RECT 1631.160 3508.715 1631.620 3508.885 ;
        RECT 1645.420 3508.715 1645.880 3508.885 ;
        RECT 1659.680 3508.715 1660.140 3508.885 ;
        RECT 1673.940 3508.715 1674.400 3508.885 ;
        RECT 1688.200 3508.715 1688.660 3508.885 ;
        RECT 1702.460 3508.715 1702.920 3508.885 ;
        RECT 1716.720 3508.715 1717.180 3508.885 ;
        RECT 1730.980 3508.715 1731.440 3508.885 ;
        RECT 1745.240 3508.715 1745.700 3508.885 ;
        RECT 1759.500 3508.715 1759.960 3508.885 ;
        RECT 1773.760 3508.715 1774.220 3508.885 ;
        RECT 1788.020 3508.715 1788.480 3508.885 ;
        RECT 1802.280 3508.715 1802.740 3508.885 ;
        RECT 1816.540 3508.715 1817.000 3508.885 ;
        RECT 1830.800 3508.715 1831.260 3508.885 ;
        RECT 1845.060 3508.715 1845.520 3508.885 ;
        RECT 1859.320 3508.715 1859.780 3508.885 ;
        RECT 1873.580 3508.715 1874.040 3508.885 ;
        RECT 1887.840 3508.715 1888.300 3508.885 ;
        RECT 1902.100 3508.715 1902.560 3508.885 ;
        RECT 1916.360 3508.715 1916.820 3508.885 ;
        RECT 1930.620 3508.715 1931.080 3508.885 ;
        RECT 1944.880 3508.715 1945.340 3508.885 ;
        RECT 1959.140 3508.715 1959.600 3508.885 ;
        RECT 1973.400 3508.715 1973.860 3508.885 ;
        RECT 1987.660 3508.715 1988.120 3508.885 ;
        RECT 2001.920 3508.715 2002.380 3508.885 ;
        RECT 2016.180 3508.715 2016.640 3508.885 ;
        RECT 2030.440 3508.715 2030.900 3508.885 ;
        RECT 2044.700 3508.715 2045.160 3508.885 ;
        RECT 2058.960 3508.715 2059.420 3508.885 ;
        RECT 2073.220 3508.715 2073.680 3508.885 ;
        RECT 2087.480 3508.715 2087.940 3508.885 ;
        RECT 2101.740 3508.715 2102.200 3508.885 ;
        RECT 2116.000 3508.715 2116.460 3508.885 ;
        RECT 2130.260 3508.715 2130.720 3508.885 ;
        RECT 2144.520 3508.715 2144.980 3508.885 ;
        RECT 2158.780 3508.715 2159.240 3508.885 ;
        RECT 2173.040 3508.715 2173.500 3508.885 ;
        RECT 2187.300 3508.715 2187.760 3508.885 ;
        RECT 2201.560 3508.715 2202.020 3508.885 ;
        RECT 2215.820 3508.715 2216.280 3508.885 ;
        RECT 2230.080 3508.715 2230.540 3508.885 ;
        RECT 2244.340 3508.715 2244.800 3508.885 ;
        RECT 2258.600 3508.715 2259.060 3508.885 ;
        RECT 2272.860 3508.715 2273.320 3508.885 ;
        RECT 2287.120 3508.715 2287.580 3508.885 ;
        RECT 2301.380 3508.715 2301.840 3508.885 ;
        RECT 2315.640 3508.715 2316.100 3508.885 ;
        RECT 2329.900 3508.715 2330.360 3508.885 ;
        RECT 2344.160 3508.715 2344.620 3508.885 ;
        RECT 2358.420 3508.715 2358.880 3508.885 ;
        RECT 2372.680 3508.715 2373.140 3508.885 ;
        RECT 2386.940 3508.715 2387.400 3508.885 ;
        RECT 2401.200 3508.715 2401.660 3508.885 ;
        RECT 2415.460 3508.715 2415.920 3508.885 ;
        RECT 2429.720 3508.715 2430.180 3508.885 ;
        RECT 2443.980 3508.715 2444.440 3508.885 ;
        RECT 2458.240 3508.715 2458.700 3508.885 ;
        RECT 2472.500 3508.715 2472.960 3508.885 ;
        RECT 2486.760 3508.715 2487.220 3508.885 ;
        RECT 2501.020 3508.715 2501.480 3508.885 ;
        RECT 2515.280 3508.715 2515.740 3508.885 ;
        RECT 2529.540 3508.715 2530.000 3508.885 ;
        RECT 2543.800 3508.715 2544.260 3508.885 ;
        RECT 2558.060 3508.715 2558.520 3508.885 ;
        RECT 2572.320 3508.715 2572.780 3508.885 ;
        RECT 2586.580 3508.715 2587.040 3508.885 ;
        RECT 2600.840 3508.715 2601.300 3508.885 ;
        RECT 2615.100 3508.715 2615.560 3508.885 ;
        RECT 2629.360 3508.715 2629.820 3508.885 ;
        RECT 2643.620 3508.715 2644.080 3508.885 ;
        RECT 2657.880 3508.715 2658.340 3508.885 ;
        RECT 2672.140 3508.715 2672.600 3508.885 ;
        RECT 2686.400 3508.715 2686.860 3508.885 ;
        RECT 2700.660 3508.715 2701.120 3508.885 ;
        RECT 2714.920 3508.715 2715.380 3508.885 ;
        RECT 2729.180 3508.715 2729.640 3508.885 ;
        RECT 2743.440 3508.715 2743.900 3508.885 ;
        RECT 2757.700 3508.715 2758.160 3508.885 ;
        RECT 2771.960 3508.715 2772.420 3508.885 ;
        RECT 2786.220 3508.715 2786.680 3508.885 ;
        RECT 2800.480 3508.715 2800.940 3508.885 ;
        RECT 2814.740 3508.715 2815.200 3508.885 ;
        RECT 2829.000 3508.715 2829.460 3508.885 ;
        RECT 2843.260 3508.715 2843.720 3508.885 ;
        RECT 2857.520 3508.715 2857.980 3508.885 ;
        RECT 2871.780 3508.715 2872.240 3508.885 ;
        RECT 2886.040 3508.715 2886.500 3508.885 ;
        RECT 2900.300 3508.715 2900.760 3508.885 ;
        RECT 2912.720 3508.715 2914.100 3508.885 ;
        RECT 5.605 3507.625 6.815 3508.715 ;
        RECT 6.295 3507.085 6.815 3507.625 ;
        RECT 19.865 3507.550 20.155 3508.715 ;
        RECT 34.125 3507.550 34.415 3508.715 ;
        RECT 48.385 3507.550 48.675 3508.715 ;
        RECT 62.645 3507.550 62.935 3508.715 ;
        RECT 76.905 3507.550 77.195 3508.715 ;
        RECT 91.165 3507.550 91.455 3508.715 ;
        RECT 105.425 3507.550 105.715 3508.715 ;
        RECT 119.685 3507.550 119.975 3508.715 ;
        RECT 133.945 3507.550 134.235 3508.715 ;
        RECT 148.205 3507.550 148.495 3508.715 ;
        RECT 162.465 3507.550 162.755 3508.715 ;
        RECT 176.725 3507.550 177.015 3508.715 ;
        RECT 190.985 3507.550 191.275 3508.715 ;
        RECT 205.245 3507.550 205.535 3508.715 ;
        RECT 219.505 3507.550 219.795 3508.715 ;
        RECT 233.765 3507.550 234.055 3508.715 ;
        RECT 248.025 3507.550 248.315 3508.715 ;
        RECT 262.285 3507.550 262.575 3508.715 ;
        RECT 276.545 3507.550 276.835 3508.715 ;
        RECT 290.805 3507.550 291.095 3508.715 ;
        RECT 305.065 3507.550 305.355 3508.715 ;
        RECT 319.325 3507.550 319.615 3508.715 ;
        RECT 333.585 3507.550 333.875 3508.715 ;
        RECT 347.845 3507.550 348.135 3508.715 ;
        RECT 362.105 3507.550 362.395 3508.715 ;
        RECT 376.365 3507.550 376.655 3508.715 ;
        RECT 390.625 3507.550 390.915 3508.715 ;
        RECT 404.885 3507.550 405.175 3508.715 ;
        RECT 419.145 3507.550 419.435 3508.715 ;
        RECT 433.405 3507.550 433.695 3508.715 ;
        RECT 447.665 3507.550 447.955 3508.715 ;
        RECT 461.925 3507.550 462.215 3508.715 ;
        RECT 476.185 3507.550 476.475 3508.715 ;
        RECT 490.445 3507.550 490.735 3508.715 ;
        RECT 504.705 3507.550 504.995 3508.715 ;
        RECT 518.965 3507.550 519.255 3508.715 ;
        RECT 533.225 3507.550 533.515 3508.715 ;
        RECT 547.485 3507.550 547.775 3508.715 ;
        RECT 561.745 3507.550 562.035 3508.715 ;
        RECT 576.005 3507.550 576.295 3508.715 ;
        RECT 590.265 3507.550 590.555 3508.715 ;
        RECT 604.525 3507.550 604.815 3508.715 ;
        RECT 618.785 3507.550 619.075 3508.715 ;
        RECT 633.045 3507.550 633.335 3508.715 ;
        RECT 647.305 3507.550 647.595 3508.715 ;
        RECT 661.565 3507.550 661.855 3508.715 ;
        RECT 675.825 3507.550 676.115 3508.715 ;
        RECT 690.085 3507.550 690.375 3508.715 ;
        RECT 704.345 3507.550 704.635 3508.715 ;
        RECT 718.605 3507.550 718.895 3508.715 ;
        RECT 732.865 3507.550 733.155 3508.715 ;
        RECT 747.125 3507.550 747.415 3508.715 ;
        RECT 761.385 3507.550 761.675 3508.715 ;
        RECT 775.645 3507.550 775.935 3508.715 ;
        RECT 789.905 3507.550 790.195 3508.715 ;
        RECT 804.165 3507.550 804.455 3508.715 ;
        RECT 818.425 3507.550 818.715 3508.715 ;
        RECT 832.685 3507.550 832.975 3508.715 ;
        RECT 846.945 3507.550 847.235 3508.715 ;
        RECT 861.205 3507.550 861.495 3508.715 ;
        RECT 875.465 3507.550 875.755 3508.715 ;
        RECT 889.725 3507.550 890.015 3508.715 ;
        RECT 903.985 3507.550 904.275 3508.715 ;
        RECT 918.245 3507.550 918.535 3508.715 ;
        RECT 932.505 3507.550 932.795 3508.715 ;
        RECT 946.765 3507.550 947.055 3508.715 ;
        RECT 961.025 3507.550 961.315 3508.715 ;
        RECT 975.285 3507.550 975.575 3508.715 ;
        RECT 989.545 3507.550 989.835 3508.715 ;
        RECT 1003.805 3507.550 1004.095 3508.715 ;
        RECT 1018.065 3507.550 1018.355 3508.715 ;
        RECT 1032.325 3507.550 1032.615 3508.715 ;
        RECT 1046.585 3507.550 1046.875 3508.715 ;
        RECT 1060.845 3507.550 1061.135 3508.715 ;
        RECT 1075.105 3507.550 1075.395 3508.715 ;
        RECT 1089.365 3507.550 1089.655 3508.715 ;
        RECT 1103.625 3507.550 1103.915 3508.715 ;
        RECT 1117.885 3507.550 1118.175 3508.715 ;
        RECT 1132.145 3507.550 1132.435 3508.715 ;
        RECT 1146.405 3507.550 1146.695 3508.715 ;
        RECT 1160.665 3507.550 1160.955 3508.715 ;
        RECT 1174.925 3507.550 1175.215 3508.715 ;
        RECT 1189.185 3507.550 1189.475 3508.715 ;
        RECT 1203.445 3507.550 1203.735 3508.715 ;
        RECT 1217.705 3507.550 1217.995 3508.715 ;
        RECT 1231.965 3507.550 1232.255 3508.715 ;
        RECT 1246.225 3507.550 1246.515 3508.715 ;
        RECT 1260.485 3507.550 1260.775 3508.715 ;
        RECT 1274.745 3507.550 1275.035 3508.715 ;
        RECT 1289.005 3507.550 1289.295 3508.715 ;
        RECT 1303.265 3507.550 1303.555 3508.715 ;
        RECT 1317.525 3507.550 1317.815 3508.715 ;
        RECT 1331.785 3507.550 1332.075 3508.715 ;
        RECT 1346.045 3507.550 1346.335 3508.715 ;
        RECT 1360.305 3507.550 1360.595 3508.715 ;
        RECT 1374.565 3507.550 1374.855 3508.715 ;
        RECT 1388.825 3507.550 1389.115 3508.715 ;
        RECT 1403.085 3507.550 1403.375 3508.715 ;
        RECT 1417.345 3507.550 1417.635 3508.715 ;
        RECT 1431.605 3507.550 1431.895 3508.715 ;
        RECT 1445.865 3507.550 1446.155 3508.715 ;
        RECT 1460.125 3507.550 1460.415 3508.715 ;
        RECT 1474.385 3507.550 1474.675 3508.715 ;
        RECT 1488.645 3507.550 1488.935 3508.715 ;
        RECT 1502.905 3507.550 1503.195 3508.715 ;
        RECT 1517.165 3507.550 1517.455 3508.715 ;
        RECT 1531.425 3507.550 1531.715 3508.715 ;
        RECT 1545.685 3507.550 1545.975 3508.715 ;
        RECT 1559.945 3507.550 1560.235 3508.715 ;
        RECT 1574.205 3507.550 1574.495 3508.715 ;
        RECT 1588.465 3507.550 1588.755 3508.715 ;
        RECT 1602.725 3507.550 1603.015 3508.715 ;
        RECT 1616.985 3507.550 1617.275 3508.715 ;
        RECT 1631.245 3507.550 1631.535 3508.715 ;
        RECT 1645.505 3507.550 1645.795 3508.715 ;
        RECT 1659.765 3507.550 1660.055 3508.715 ;
        RECT 1674.025 3507.550 1674.315 3508.715 ;
        RECT 1688.285 3507.550 1688.575 3508.715 ;
        RECT 1702.545 3507.550 1702.835 3508.715 ;
        RECT 1716.805 3507.550 1717.095 3508.715 ;
        RECT 1731.065 3507.550 1731.355 3508.715 ;
        RECT 1745.325 3507.550 1745.615 3508.715 ;
        RECT 1759.585 3507.550 1759.875 3508.715 ;
        RECT 1773.845 3507.550 1774.135 3508.715 ;
        RECT 1788.105 3507.550 1788.395 3508.715 ;
        RECT 1802.365 3507.550 1802.655 3508.715 ;
        RECT 1816.625 3507.550 1816.915 3508.715 ;
        RECT 1830.885 3507.550 1831.175 3508.715 ;
        RECT 1845.145 3507.550 1845.435 3508.715 ;
        RECT 1859.405 3507.550 1859.695 3508.715 ;
        RECT 1873.665 3507.550 1873.955 3508.715 ;
        RECT 1887.925 3507.550 1888.215 3508.715 ;
        RECT 1902.185 3507.550 1902.475 3508.715 ;
        RECT 1916.445 3507.550 1916.735 3508.715 ;
        RECT 1930.705 3507.550 1930.995 3508.715 ;
        RECT 1944.965 3507.550 1945.255 3508.715 ;
        RECT 1959.225 3507.550 1959.515 3508.715 ;
        RECT 1973.485 3507.550 1973.775 3508.715 ;
        RECT 1987.745 3507.550 1988.035 3508.715 ;
        RECT 2002.005 3507.550 2002.295 3508.715 ;
        RECT 2016.265 3507.550 2016.555 3508.715 ;
        RECT 2030.525 3507.550 2030.815 3508.715 ;
        RECT 2044.785 3507.550 2045.075 3508.715 ;
        RECT 2059.045 3507.550 2059.335 3508.715 ;
        RECT 2073.305 3507.550 2073.595 3508.715 ;
        RECT 2087.565 3507.550 2087.855 3508.715 ;
        RECT 2101.825 3507.550 2102.115 3508.715 ;
        RECT 2116.085 3507.550 2116.375 3508.715 ;
        RECT 2130.345 3507.550 2130.635 3508.715 ;
        RECT 2144.605 3507.550 2144.895 3508.715 ;
        RECT 2158.865 3507.550 2159.155 3508.715 ;
        RECT 2173.125 3507.550 2173.415 3508.715 ;
        RECT 2187.385 3507.550 2187.675 3508.715 ;
        RECT 2201.645 3507.550 2201.935 3508.715 ;
        RECT 2215.905 3507.550 2216.195 3508.715 ;
        RECT 2230.165 3507.550 2230.455 3508.715 ;
        RECT 2244.425 3507.550 2244.715 3508.715 ;
        RECT 2258.685 3507.550 2258.975 3508.715 ;
        RECT 2272.945 3507.550 2273.235 3508.715 ;
        RECT 2287.205 3507.550 2287.495 3508.715 ;
        RECT 2301.465 3507.550 2301.755 3508.715 ;
        RECT 2315.725 3507.550 2316.015 3508.715 ;
        RECT 2329.985 3507.550 2330.275 3508.715 ;
        RECT 2344.245 3507.550 2344.535 3508.715 ;
        RECT 2358.505 3507.550 2358.795 3508.715 ;
        RECT 2372.765 3507.550 2373.055 3508.715 ;
        RECT 2387.025 3507.550 2387.315 3508.715 ;
        RECT 2401.285 3507.550 2401.575 3508.715 ;
        RECT 2415.545 3507.550 2415.835 3508.715 ;
        RECT 2429.805 3507.550 2430.095 3508.715 ;
        RECT 2444.065 3507.550 2444.355 3508.715 ;
        RECT 2458.325 3507.550 2458.615 3508.715 ;
        RECT 2472.585 3507.550 2472.875 3508.715 ;
        RECT 2486.845 3507.550 2487.135 3508.715 ;
        RECT 2501.105 3507.550 2501.395 3508.715 ;
        RECT 2515.365 3507.550 2515.655 3508.715 ;
        RECT 2529.625 3507.550 2529.915 3508.715 ;
        RECT 2543.885 3507.550 2544.175 3508.715 ;
        RECT 2558.145 3507.550 2558.435 3508.715 ;
        RECT 2572.405 3507.550 2572.695 3508.715 ;
        RECT 2586.665 3507.550 2586.955 3508.715 ;
        RECT 2600.925 3507.550 2601.215 3508.715 ;
        RECT 2615.185 3507.550 2615.475 3508.715 ;
        RECT 2629.445 3507.550 2629.735 3508.715 ;
        RECT 2643.705 3507.550 2643.995 3508.715 ;
        RECT 2657.965 3507.550 2658.255 3508.715 ;
        RECT 2672.225 3507.550 2672.515 3508.715 ;
        RECT 2686.485 3507.550 2686.775 3508.715 ;
        RECT 2700.745 3507.550 2701.035 3508.715 ;
        RECT 2715.005 3507.550 2715.295 3508.715 ;
        RECT 2729.265 3507.550 2729.555 3508.715 ;
        RECT 2743.525 3507.550 2743.815 3508.715 ;
        RECT 2757.785 3507.550 2758.075 3508.715 ;
        RECT 2772.045 3507.550 2772.335 3508.715 ;
        RECT 2786.305 3507.550 2786.595 3508.715 ;
        RECT 2800.565 3507.550 2800.855 3508.715 ;
        RECT 2814.825 3507.550 2815.115 3508.715 ;
        RECT 2829.085 3507.550 2829.375 3508.715 ;
        RECT 2843.345 3507.550 2843.635 3508.715 ;
        RECT 2857.605 3507.550 2857.895 3508.715 ;
        RECT 2871.865 3507.550 2872.155 3508.715 ;
        RECT 2886.125 3507.550 2886.415 3508.715 ;
        RECT 2900.385 3507.550 2900.675 3508.715 ;
        RECT 2912.805 3507.625 2914.015 3508.715 ;
        RECT 2912.805 3507.085 2913.325 3507.625 ;
        RECT 6.295 3504.535 6.815 3505.075 ;
        RECT 5.605 3503.445 6.815 3504.535 ;
        RECT 2912.805 3504.535 2913.325 3505.075 ;
        RECT 9.935 3503.445 10.265 3504.170 ;
        RECT 11.315 3503.445 11.645 3504.170 ;
        RECT 2909.315 3503.445 2909.645 3504.170 ;
        RECT 2910.695 3503.445 2911.025 3504.170 ;
        RECT 2912.805 3503.445 2914.015 3504.535 ;
        RECT 5.520 3503.275 6.900 3503.445 ;
        RECT 9.660 3503.275 12.420 3503.445 ;
        RECT 2909.040 3503.275 2911.800 3503.445 ;
        RECT 2912.720 3503.275 2914.100 3503.445 ;
        RECT 5.605 3502.185 6.815 3503.275 ;
        RECT 6.295 3501.645 6.815 3502.185 ;
        RECT 2910.045 3502.110 2910.335 3503.275 ;
        RECT 2912.805 3502.185 2914.015 3503.275 ;
        RECT 2912.805 3501.645 2913.325 3502.185 ;
        RECT 6.295 3499.095 6.815 3499.635 ;
        RECT 5.605 3498.005 6.815 3499.095 ;
        RECT 2912.805 3499.095 2913.325 3499.635 ;
        RECT 2912.805 3498.005 2914.015 3499.095 ;
        RECT 5.520 3497.835 6.900 3498.005 ;
        RECT 2909.960 3497.835 2910.420 3498.005 ;
        RECT 2912.720 3497.835 2914.100 3498.005 ;
        RECT 5.605 3496.745 6.815 3497.835 ;
        RECT 6.295 3496.205 6.815 3496.745 ;
        RECT 2910.045 3496.670 2910.335 3497.835 ;
        RECT 2912.805 3496.745 2914.015 3497.835 ;
        RECT 2912.805 3496.205 2913.325 3496.745 ;
        RECT 6.295 3493.655 6.815 3494.195 ;
        RECT 5.605 3492.565 6.815 3493.655 ;
        RECT 2912.805 3493.655 2913.325 3494.195 ;
        RECT 2912.805 3492.565 2914.015 3493.655 ;
        RECT 5.520 3492.395 6.900 3492.565 ;
        RECT 2909.960 3492.395 2910.420 3492.565 ;
        RECT 2912.720 3492.395 2914.100 3492.565 ;
        RECT 5.605 3491.305 6.815 3492.395 ;
        RECT 6.295 3490.765 6.815 3491.305 ;
        RECT 2910.045 3491.230 2910.335 3492.395 ;
        RECT 2912.805 3491.305 2914.015 3492.395 ;
        RECT 2912.805 3490.765 2913.325 3491.305 ;
        RECT 6.295 3488.215 6.815 3488.755 ;
        RECT 5.605 3487.125 6.815 3488.215 ;
        RECT 2912.805 3488.215 2913.325 3488.755 ;
        RECT 2912.805 3487.125 2914.015 3488.215 ;
        RECT 5.520 3486.955 6.900 3487.125 ;
        RECT 2909.960 3486.955 2910.420 3487.125 ;
        RECT 2912.720 3486.955 2914.100 3487.125 ;
        RECT 5.605 3485.865 6.815 3486.955 ;
        RECT 6.295 3485.325 6.815 3485.865 ;
        RECT 2910.045 3485.790 2910.335 3486.955 ;
        RECT 2912.805 3485.865 2914.015 3486.955 ;
        RECT 2912.805 3485.325 2913.325 3485.865 ;
        RECT 6.295 3482.775 6.815 3483.315 ;
        RECT 5.605 3481.685 6.815 3482.775 ;
        RECT 2912.805 3482.775 2913.325 3483.315 ;
        RECT 2912.805 3481.685 2914.015 3482.775 ;
        RECT 5.520 3481.515 6.900 3481.685 ;
        RECT 2909.960 3481.515 2910.420 3481.685 ;
        RECT 2912.720 3481.515 2914.100 3481.685 ;
        RECT 5.605 3480.425 6.815 3481.515 ;
        RECT 6.295 3479.885 6.815 3480.425 ;
        RECT 2910.045 3480.350 2910.335 3481.515 ;
        RECT 2912.805 3480.425 2914.015 3481.515 ;
        RECT 2912.805 3479.885 2913.325 3480.425 ;
        RECT 6.295 3477.335 6.815 3477.875 ;
        RECT 5.605 3476.245 6.815 3477.335 ;
        RECT 2912.805 3477.335 2913.325 3477.875 ;
        RECT 2912.805 3476.245 2914.015 3477.335 ;
        RECT 5.520 3476.075 6.900 3476.245 ;
        RECT 2909.960 3476.075 2910.420 3476.245 ;
        RECT 2912.720 3476.075 2914.100 3476.245 ;
        RECT 5.605 3474.985 6.815 3476.075 ;
        RECT 6.295 3474.445 6.815 3474.985 ;
        RECT 2910.045 3474.910 2910.335 3476.075 ;
        RECT 2912.805 3474.985 2914.015 3476.075 ;
        RECT 2912.805 3474.445 2913.325 3474.985 ;
        RECT 6.295 3471.895 6.815 3472.435 ;
        RECT 5.605 3470.805 6.815 3471.895 ;
        RECT 2912.805 3471.895 2913.325 3472.435 ;
        RECT 2912.805 3470.805 2914.015 3471.895 ;
        RECT 5.520 3470.635 6.900 3470.805 ;
        RECT 2909.960 3470.635 2910.420 3470.805 ;
        RECT 2912.720 3470.635 2914.100 3470.805 ;
        RECT 5.605 3469.545 6.815 3470.635 ;
        RECT 6.295 3469.005 6.815 3469.545 ;
        RECT 2910.045 3469.470 2910.335 3470.635 ;
        RECT 2912.805 3469.545 2914.015 3470.635 ;
        RECT 2912.805 3469.005 2913.325 3469.545 ;
        RECT 6.295 3466.455 6.815 3466.995 ;
        RECT 5.605 3465.365 6.815 3466.455 ;
        RECT 2912.805 3466.455 2913.325 3466.995 ;
        RECT 2912.805 3465.365 2914.015 3466.455 ;
        RECT 5.520 3465.195 6.900 3465.365 ;
        RECT 2909.960 3465.195 2910.420 3465.365 ;
        RECT 2912.720 3465.195 2914.100 3465.365 ;
        RECT 5.605 3464.105 6.815 3465.195 ;
        RECT 6.295 3463.565 6.815 3464.105 ;
        RECT 2910.045 3464.030 2910.335 3465.195 ;
        RECT 2912.805 3464.105 2914.015 3465.195 ;
        RECT 2912.805 3463.565 2913.325 3464.105 ;
        RECT 6.295 3461.015 6.815 3461.555 ;
        RECT 5.605 3459.925 6.815 3461.015 ;
        RECT 2912.805 3461.015 2913.325 3461.555 ;
        RECT 2912.805 3459.925 2914.015 3461.015 ;
        RECT 5.520 3459.755 6.900 3459.925 ;
        RECT 2909.960 3459.755 2910.420 3459.925 ;
        RECT 2912.720 3459.755 2914.100 3459.925 ;
        RECT 5.605 3458.665 6.815 3459.755 ;
        RECT 6.295 3458.125 6.815 3458.665 ;
        RECT 2910.045 3458.590 2910.335 3459.755 ;
        RECT 2912.805 3458.665 2914.015 3459.755 ;
        RECT 2912.805 3458.125 2913.325 3458.665 ;
        RECT 6.295 3455.575 6.815 3456.115 ;
        RECT 5.605 3454.485 6.815 3455.575 ;
        RECT 2912.805 3455.575 2913.325 3456.115 ;
        RECT 2912.805 3454.485 2914.015 3455.575 ;
        RECT 5.520 3454.315 6.900 3454.485 ;
        RECT 2909.960 3454.315 2910.420 3454.485 ;
        RECT 2912.720 3454.315 2914.100 3454.485 ;
        RECT 5.605 3453.225 6.815 3454.315 ;
        RECT 6.295 3452.685 6.815 3453.225 ;
        RECT 2910.045 3453.150 2910.335 3454.315 ;
        RECT 2912.805 3453.225 2914.015 3454.315 ;
        RECT 2912.805 3452.685 2913.325 3453.225 ;
        RECT 6.295 3450.135 6.815 3450.675 ;
        RECT 5.605 3449.045 6.815 3450.135 ;
        RECT 2912.805 3450.135 2913.325 3450.675 ;
        RECT 2912.805 3449.045 2914.015 3450.135 ;
        RECT 5.520 3448.875 6.900 3449.045 ;
        RECT 2909.960 3448.875 2910.420 3449.045 ;
        RECT 2912.720 3448.875 2914.100 3449.045 ;
        RECT 5.605 3447.785 6.815 3448.875 ;
        RECT 6.295 3447.245 6.815 3447.785 ;
        RECT 2910.045 3447.710 2910.335 3448.875 ;
        RECT 2912.805 3447.785 2914.015 3448.875 ;
        RECT 2912.805 3447.245 2913.325 3447.785 ;
        RECT 6.295 3444.695 6.815 3445.235 ;
        RECT 5.605 3443.605 6.815 3444.695 ;
        RECT 2912.805 3444.695 2913.325 3445.235 ;
        RECT 2912.805 3443.605 2914.015 3444.695 ;
        RECT 5.520 3443.435 6.900 3443.605 ;
        RECT 2909.960 3443.435 2910.420 3443.605 ;
        RECT 2912.720 3443.435 2914.100 3443.605 ;
        RECT 5.605 3442.345 6.815 3443.435 ;
        RECT 6.295 3441.805 6.815 3442.345 ;
        RECT 2910.045 3442.270 2910.335 3443.435 ;
        RECT 2912.805 3442.345 2914.015 3443.435 ;
        RECT 2912.805 3441.805 2913.325 3442.345 ;
        RECT 6.295 3439.255 6.815 3439.795 ;
        RECT 5.605 3438.165 6.815 3439.255 ;
        RECT 2912.805 3439.255 2913.325 3439.795 ;
        RECT 2912.805 3438.165 2914.015 3439.255 ;
        RECT 5.520 3437.995 6.900 3438.165 ;
        RECT 2909.960 3437.995 2910.420 3438.165 ;
        RECT 2912.720 3437.995 2914.100 3438.165 ;
        RECT 5.605 3436.905 6.815 3437.995 ;
        RECT 6.295 3436.365 6.815 3436.905 ;
        RECT 2910.045 3436.830 2910.335 3437.995 ;
        RECT 2912.805 3436.905 2914.015 3437.995 ;
        RECT 2912.805 3436.365 2913.325 3436.905 ;
        RECT 6.295 3433.815 6.815 3434.355 ;
        RECT 5.605 3432.725 6.815 3433.815 ;
        RECT 2912.805 3433.815 2913.325 3434.355 ;
        RECT 2912.805 3432.725 2914.015 3433.815 ;
        RECT 5.520 3432.555 6.900 3432.725 ;
        RECT 2909.960 3432.555 2910.420 3432.725 ;
        RECT 2912.720 3432.555 2914.100 3432.725 ;
        RECT 5.605 3431.465 6.815 3432.555 ;
        RECT 6.295 3430.925 6.815 3431.465 ;
        RECT 2910.045 3431.390 2910.335 3432.555 ;
        RECT 2912.805 3431.465 2914.015 3432.555 ;
        RECT 2912.805 3430.925 2913.325 3431.465 ;
        RECT 6.295 3428.375 6.815 3428.915 ;
        RECT 5.605 3427.285 6.815 3428.375 ;
        RECT 2912.805 3428.375 2913.325 3428.915 ;
        RECT 2912.805 3427.285 2914.015 3428.375 ;
        RECT 5.520 3427.115 6.900 3427.285 ;
        RECT 2909.960 3427.115 2910.420 3427.285 ;
        RECT 2912.720 3427.115 2914.100 3427.285 ;
        RECT 5.605 3426.025 6.815 3427.115 ;
        RECT 6.295 3425.485 6.815 3426.025 ;
        RECT 2910.045 3425.950 2910.335 3427.115 ;
        RECT 2912.805 3426.025 2914.015 3427.115 ;
        RECT 2912.805 3425.485 2913.325 3426.025 ;
        RECT 6.295 3422.935 6.815 3423.475 ;
        RECT 5.605 3421.845 6.815 3422.935 ;
        RECT 2912.805 3422.935 2913.325 3423.475 ;
        RECT 2912.805 3421.845 2914.015 3422.935 ;
        RECT 5.520 3421.675 6.900 3421.845 ;
        RECT 2909.960 3421.675 2910.420 3421.845 ;
        RECT 2912.720 3421.675 2914.100 3421.845 ;
        RECT 5.605 3420.585 6.815 3421.675 ;
        RECT 6.295 3420.045 6.815 3420.585 ;
        RECT 2910.045 3420.510 2910.335 3421.675 ;
        RECT 2912.805 3420.585 2914.015 3421.675 ;
        RECT 2912.805 3420.045 2913.325 3420.585 ;
        RECT 6.295 3417.495 6.815 3418.035 ;
        RECT 5.605 3416.405 6.815 3417.495 ;
        RECT 2912.805 3417.495 2913.325 3418.035 ;
        RECT 2912.805 3416.405 2914.015 3417.495 ;
        RECT 5.520 3416.235 6.900 3416.405 ;
        RECT 2909.960 3416.235 2910.420 3416.405 ;
        RECT 2912.720 3416.235 2914.100 3416.405 ;
        RECT 5.605 3415.145 6.815 3416.235 ;
        RECT 6.295 3414.605 6.815 3415.145 ;
        RECT 2910.045 3415.070 2910.335 3416.235 ;
        RECT 2912.805 3415.145 2914.015 3416.235 ;
        RECT 2912.805 3414.605 2913.325 3415.145 ;
        RECT 6.295 3412.055 6.815 3412.595 ;
        RECT 5.605 3410.965 6.815 3412.055 ;
        RECT 2912.805 3412.055 2913.325 3412.595 ;
        RECT 2912.805 3410.965 2914.015 3412.055 ;
        RECT 5.520 3410.795 6.900 3410.965 ;
        RECT 2909.960 3410.795 2910.420 3410.965 ;
        RECT 2912.720 3410.795 2914.100 3410.965 ;
        RECT 5.605 3409.705 6.815 3410.795 ;
        RECT 6.295 3409.165 6.815 3409.705 ;
        RECT 2910.045 3409.630 2910.335 3410.795 ;
        RECT 2912.805 3409.705 2914.015 3410.795 ;
        RECT 2912.805 3409.165 2913.325 3409.705 ;
        RECT 6.295 3406.615 6.815 3407.155 ;
        RECT 5.605 3405.525 6.815 3406.615 ;
        RECT 2912.805 3406.615 2913.325 3407.155 ;
        RECT 2912.805 3405.525 2914.015 3406.615 ;
        RECT 5.520 3405.355 6.900 3405.525 ;
        RECT 2909.960 3405.355 2910.420 3405.525 ;
        RECT 2912.720 3405.355 2914.100 3405.525 ;
        RECT 5.605 3404.265 6.815 3405.355 ;
        RECT 6.295 3403.725 6.815 3404.265 ;
        RECT 2910.045 3404.190 2910.335 3405.355 ;
        RECT 2912.805 3404.265 2914.015 3405.355 ;
        RECT 2912.805 3403.725 2913.325 3404.265 ;
        RECT 6.295 3401.175 6.815 3401.715 ;
        RECT 5.605 3400.085 6.815 3401.175 ;
        RECT 2912.805 3401.175 2913.325 3401.715 ;
        RECT 2909.315 3400.085 2909.645 3400.810 ;
        RECT 2912.805 3400.085 2914.015 3401.175 ;
        RECT 5.520 3399.915 6.900 3400.085 ;
        RECT 2909.040 3399.915 2910.420 3400.085 ;
        RECT 2912.720 3399.915 2914.100 3400.085 ;
        RECT 5.605 3398.825 6.815 3399.915 ;
        RECT 6.295 3398.285 6.815 3398.825 ;
        RECT 2910.045 3398.750 2910.335 3399.915 ;
        RECT 2912.805 3398.825 2914.015 3399.915 ;
        RECT 2912.805 3398.285 2913.325 3398.825 ;
        RECT 6.295 3395.735 6.815 3396.275 ;
        RECT 5.605 3394.645 6.815 3395.735 ;
        RECT 2912.805 3395.735 2913.325 3396.275 ;
        RECT 2912.805 3394.645 2914.015 3395.735 ;
        RECT 5.520 3394.475 6.900 3394.645 ;
        RECT 2909.960 3394.475 2910.420 3394.645 ;
        RECT 2912.720 3394.475 2914.100 3394.645 ;
        RECT 5.605 3393.385 6.815 3394.475 ;
        RECT 6.295 3392.845 6.815 3393.385 ;
        RECT 2910.045 3393.310 2910.335 3394.475 ;
        RECT 2912.805 3393.385 2914.015 3394.475 ;
        RECT 2912.805 3392.845 2913.325 3393.385 ;
        RECT 6.295 3390.295 6.815 3390.835 ;
        RECT 5.605 3389.205 6.815 3390.295 ;
        RECT 2912.805 3390.295 2913.325 3390.835 ;
        RECT 2912.805 3389.205 2914.015 3390.295 ;
        RECT 5.520 3389.035 6.900 3389.205 ;
        RECT 2909.960 3389.035 2910.420 3389.205 ;
        RECT 2912.720 3389.035 2914.100 3389.205 ;
        RECT 5.605 3387.945 6.815 3389.035 ;
        RECT 6.295 3387.405 6.815 3387.945 ;
        RECT 2910.045 3387.870 2910.335 3389.035 ;
        RECT 2912.805 3387.945 2914.015 3389.035 ;
        RECT 2912.805 3387.405 2913.325 3387.945 ;
        RECT 6.295 3384.855 6.815 3385.395 ;
        RECT 5.605 3383.765 6.815 3384.855 ;
        RECT 2912.805 3384.855 2913.325 3385.395 ;
        RECT 2912.805 3383.765 2914.015 3384.855 ;
        RECT 5.520 3383.595 6.900 3383.765 ;
        RECT 2909.960 3383.595 2910.420 3383.765 ;
        RECT 2912.720 3383.595 2914.100 3383.765 ;
        RECT 5.605 3382.505 6.815 3383.595 ;
        RECT 6.295 3381.965 6.815 3382.505 ;
        RECT 2910.045 3382.430 2910.335 3383.595 ;
        RECT 2912.805 3382.505 2914.015 3383.595 ;
        RECT 2912.805 3381.965 2913.325 3382.505 ;
        RECT 6.295 3379.415 6.815 3379.955 ;
        RECT 5.605 3378.325 6.815 3379.415 ;
        RECT 2912.805 3379.415 2913.325 3379.955 ;
        RECT 2912.805 3378.325 2914.015 3379.415 ;
        RECT 5.520 3378.155 6.900 3378.325 ;
        RECT 2909.960 3378.155 2910.420 3378.325 ;
        RECT 2912.720 3378.155 2914.100 3378.325 ;
        RECT 5.605 3377.065 6.815 3378.155 ;
        RECT 6.295 3376.525 6.815 3377.065 ;
        RECT 2910.045 3376.990 2910.335 3378.155 ;
        RECT 2912.805 3377.065 2914.015 3378.155 ;
        RECT 2912.805 3376.525 2913.325 3377.065 ;
        RECT 6.295 3373.975 6.815 3374.515 ;
        RECT 5.605 3372.885 6.815 3373.975 ;
        RECT 2912.805 3373.975 2913.325 3374.515 ;
        RECT 2912.805 3372.885 2914.015 3373.975 ;
        RECT 5.520 3372.715 6.900 3372.885 ;
        RECT 2909.960 3372.715 2910.420 3372.885 ;
        RECT 2912.720 3372.715 2914.100 3372.885 ;
        RECT 5.605 3371.625 6.815 3372.715 ;
        RECT 6.295 3371.085 6.815 3371.625 ;
        RECT 2910.045 3371.550 2910.335 3372.715 ;
        RECT 2912.805 3371.625 2914.015 3372.715 ;
        RECT 2912.805 3371.085 2913.325 3371.625 ;
        RECT 6.295 3368.535 6.815 3369.075 ;
        RECT 5.605 3367.445 6.815 3368.535 ;
        RECT 2912.805 3368.535 2913.325 3369.075 ;
        RECT 2912.805 3367.445 2914.015 3368.535 ;
        RECT 5.520 3367.275 6.900 3367.445 ;
        RECT 2909.960 3367.275 2911.800 3367.445 ;
        RECT 2912.720 3367.275 2914.100 3367.445 ;
        RECT 5.605 3366.185 6.815 3367.275 ;
        RECT 6.295 3365.645 6.815 3366.185 ;
        RECT 2910.045 3366.110 2910.335 3367.275 ;
        RECT 2910.695 3366.550 2911.025 3367.275 ;
        RECT 2912.805 3366.185 2914.015 3367.275 ;
        RECT 2912.805 3365.645 2913.325 3366.185 ;
        RECT 6.295 3363.095 6.815 3363.635 ;
        RECT 5.605 3362.005 6.815 3363.095 ;
        RECT 2912.805 3363.095 2913.325 3363.635 ;
        RECT 2912.805 3362.005 2914.015 3363.095 ;
        RECT 5.520 3361.835 6.900 3362.005 ;
        RECT 2909.960 3361.835 2910.420 3362.005 ;
        RECT 2912.720 3361.835 2914.100 3362.005 ;
        RECT 5.605 3360.745 6.815 3361.835 ;
        RECT 6.295 3360.205 6.815 3360.745 ;
        RECT 2910.045 3360.670 2910.335 3361.835 ;
        RECT 2912.805 3360.745 2914.015 3361.835 ;
        RECT 2912.805 3360.205 2913.325 3360.745 ;
        RECT 6.295 3357.655 6.815 3358.195 ;
        RECT 5.605 3356.565 6.815 3357.655 ;
        RECT 2912.805 3357.655 2913.325 3358.195 ;
        RECT 2912.805 3356.565 2914.015 3357.655 ;
        RECT 5.520 3356.395 6.900 3356.565 ;
        RECT 2909.960 3356.395 2910.420 3356.565 ;
        RECT 2912.720 3356.395 2914.100 3356.565 ;
        RECT 5.605 3355.305 6.815 3356.395 ;
        RECT 6.295 3354.765 6.815 3355.305 ;
        RECT 2910.045 3355.230 2910.335 3356.395 ;
        RECT 2912.805 3355.305 2914.015 3356.395 ;
        RECT 2912.805 3354.765 2913.325 3355.305 ;
        RECT 6.295 3352.215 6.815 3352.755 ;
        RECT 5.605 3351.125 6.815 3352.215 ;
        RECT 2912.805 3352.215 2913.325 3352.755 ;
        RECT 2912.805 3351.125 2914.015 3352.215 ;
        RECT 5.520 3350.955 6.900 3351.125 ;
        RECT 2909.960 3350.955 2910.420 3351.125 ;
        RECT 2912.720 3350.955 2914.100 3351.125 ;
        RECT 5.605 3349.865 6.815 3350.955 ;
        RECT 6.295 3349.325 6.815 3349.865 ;
        RECT 2910.045 3349.790 2910.335 3350.955 ;
        RECT 2912.805 3349.865 2914.015 3350.955 ;
        RECT 2912.805 3349.325 2913.325 3349.865 ;
        RECT 6.295 3346.775 6.815 3347.315 ;
        RECT 5.605 3345.685 6.815 3346.775 ;
        RECT 2912.805 3346.775 2913.325 3347.315 ;
        RECT 2912.805 3345.685 2914.015 3346.775 ;
        RECT 5.520 3345.515 6.900 3345.685 ;
        RECT 2909.960 3345.515 2910.420 3345.685 ;
        RECT 2912.720 3345.515 2914.100 3345.685 ;
        RECT 5.605 3344.425 6.815 3345.515 ;
        RECT 6.295 3343.885 6.815 3344.425 ;
        RECT 2910.045 3344.350 2910.335 3345.515 ;
        RECT 2912.805 3344.425 2914.015 3345.515 ;
        RECT 2912.805 3343.885 2913.325 3344.425 ;
        RECT 6.295 3341.335 6.815 3341.875 ;
        RECT 5.605 3340.245 6.815 3341.335 ;
        RECT 2912.805 3341.335 2913.325 3341.875 ;
        RECT 2912.805 3340.245 2914.015 3341.335 ;
        RECT 5.520 3340.075 6.900 3340.245 ;
        RECT 2909.960 3340.075 2910.420 3340.245 ;
        RECT 2912.720 3340.075 2914.100 3340.245 ;
        RECT 5.605 3338.985 6.815 3340.075 ;
        RECT 6.295 3338.445 6.815 3338.985 ;
        RECT 2910.045 3338.910 2910.335 3340.075 ;
        RECT 2912.805 3338.985 2914.015 3340.075 ;
        RECT 2912.805 3338.445 2913.325 3338.985 ;
        RECT 6.295 3335.895 6.815 3336.435 ;
        RECT 5.605 3334.805 6.815 3335.895 ;
        RECT 2912.805 3335.895 2913.325 3336.435 ;
        RECT 2912.805 3334.805 2914.015 3335.895 ;
        RECT 5.520 3334.635 6.900 3334.805 ;
        RECT 2909.960 3334.635 2910.420 3334.805 ;
        RECT 2912.720 3334.635 2914.100 3334.805 ;
        RECT 5.605 3333.545 6.815 3334.635 ;
        RECT 6.295 3333.005 6.815 3333.545 ;
        RECT 2910.045 3333.470 2910.335 3334.635 ;
        RECT 2912.805 3333.545 2914.015 3334.635 ;
        RECT 2912.805 3333.005 2913.325 3333.545 ;
        RECT 6.295 3330.455 6.815 3330.995 ;
        RECT 5.605 3329.365 6.815 3330.455 ;
        RECT 2912.805 3330.455 2913.325 3330.995 ;
        RECT 2912.805 3329.365 2914.015 3330.455 ;
        RECT 5.520 3329.195 6.900 3329.365 ;
        RECT 2909.960 3329.195 2910.420 3329.365 ;
        RECT 2912.720 3329.195 2914.100 3329.365 ;
        RECT 5.605 3328.105 6.815 3329.195 ;
        RECT 6.295 3327.565 6.815 3328.105 ;
        RECT 2910.045 3328.030 2910.335 3329.195 ;
        RECT 2912.805 3328.105 2914.015 3329.195 ;
        RECT 2912.805 3327.565 2913.325 3328.105 ;
        RECT 6.295 3325.015 6.815 3325.555 ;
        RECT 5.605 3323.925 6.815 3325.015 ;
        RECT 2912.805 3325.015 2913.325 3325.555 ;
        RECT 2912.805 3323.925 2914.015 3325.015 ;
        RECT 5.520 3323.755 6.900 3323.925 ;
        RECT 2909.960 3323.755 2910.420 3323.925 ;
        RECT 2912.720 3323.755 2914.100 3323.925 ;
        RECT 5.605 3322.665 6.815 3323.755 ;
        RECT 6.295 3322.125 6.815 3322.665 ;
        RECT 2910.045 3322.590 2910.335 3323.755 ;
        RECT 2912.805 3322.665 2914.015 3323.755 ;
        RECT 2912.805 3322.125 2913.325 3322.665 ;
        RECT 6.295 3319.575 6.815 3320.115 ;
        RECT 5.605 3318.485 6.815 3319.575 ;
        RECT 2912.805 3319.575 2913.325 3320.115 ;
        RECT 2912.805 3318.485 2914.015 3319.575 ;
        RECT 5.520 3318.315 6.900 3318.485 ;
        RECT 2909.960 3318.315 2910.420 3318.485 ;
        RECT 2912.720 3318.315 2914.100 3318.485 ;
        RECT 5.605 3317.225 6.815 3318.315 ;
        RECT 6.295 3316.685 6.815 3317.225 ;
        RECT 2910.045 3317.150 2910.335 3318.315 ;
        RECT 2912.805 3317.225 2914.015 3318.315 ;
        RECT 2912.805 3316.685 2913.325 3317.225 ;
        RECT 6.295 3314.135 6.815 3314.675 ;
        RECT 5.605 3313.045 6.815 3314.135 ;
        RECT 2912.805 3314.135 2913.325 3314.675 ;
        RECT 2912.805 3313.045 2914.015 3314.135 ;
        RECT 5.520 3312.875 6.900 3313.045 ;
        RECT 2909.960 3312.875 2910.420 3313.045 ;
        RECT 2912.720 3312.875 2914.100 3313.045 ;
        RECT 5.605 3311.785 6.815 3312.875 ;
        RECT 6.295 3311.245 6.815 3311.785 ;
        RECT 2910.045 3311.710 2910.335 3312.875 ;
        RECT 2912.805 3311.785 2914.015 3312.875 ;
        RECT 2912.805 3311.245 2913.325 3311.785 ;
        RECT 6.295 3308.695 6.815 3309.235 ;
        RECT 5.605 3307.605 6.815 3308.695 ;
        RECT 2912.805 3308.695 2913.325 3309.235 ;
        RECT 2912.805 3307.605 2914.015 3308.695 ;
        RECT 5.520 3307.435 6.900 3307.605 ;
        RECT 2909.960 3307.435 2910.420 3307.605 ;
        RECT 2912.720 3307.435 2914.100 3307.605 ;
        RECT 5.605 3306.345 6.815 3307.435 ;
        RECT 6.295 3305.805 6.815 3306.345 ;
        RECT 2910.045 3306.270 2910.335 3307.435 ;
        RECT 2912.805 3306.345 2914.015 3307.435 ;
        RECT 2912.805 3305.805 2913.325 3306.345 ;
        RECT 6.295 3303.255 6.815 3303.795 ;
        RECT 5.605 3302.165 6.815 3303.255 ;
        RECT 2912.805 3303.255 2913.325 3303.795 ;
        RECT 2912.805 3302.165 2914.015 3303.255 ;
        RECT 5.520 3301.995 6.900 3302.165 ;
        RECT 2909.960 3301.995 2910.420 3302.165 ;
        RECT 2912.720 3301.995 2914.100 3302.165 ;
        RECT 5.605 3300.905 6.815 3301.995 ;
        RECT 6.295 3300.365 6.815 3300.905 ;
        RECT 2910.045 3300.830 2910.335 3301.995 ;
        RECT 2912.805 3300.905 2914.015 3301.995 ;
        RECT 2912.805 3300.365 2913.325 3300.905 ;
        RECT 6.295 3297.815 6.815 3298.355 ;
        RECT 5.605 3296.725 6.815 3297.815 ;
        RECT 2912.805 3297.815 2913.325 3298.355 ;
        RECT 2912.805 3296.725 2914.015 3297.815 ;
        RECT 5.520 3296.555 6.900 3296.725 ;
        RECT 2909.960 3296.555 2910.420 3296.725 ;
        RECT 2912.720 3296.555 2914.100 3296.725 ;
        RECT 5.605 3295.465 6.815 3296.555 ;
        RECT 6.295 3294.925 6.815 3295.465 ;
        RECT 2910.045 3295.390 2910.335 3296.555 ;
        RECT 2912.805 3295.465 2914.015 3296.555 ;
        RECT 2912.805 3294.925 2913.325 3295.465 ;
        RECT 6.295 3292.375 6.815 3292.915 ;
        RECT 5.605 3291.285 6.815 3292.375 ;
        RECT 2912.805 3292.375 2913.325 3292.915 ;
        RECT 2912.805 3291.285 2914.015 3292.375 ;
        RECT 5.520 3291.115 6.900 3291.285 ;
        RECT 2909.960 3291.115 2910.420 3291.285 ;
        RECT 2912.720 3291.115 2914.100 3291.285 ;
        RECT 5.605 3290.025 6.815 3291.115 ;
        RECT 6.295 3289.485 6.815 3290.025 ;
        RECT 2910.045 3289.950 2910.335 3291.115 ;
        RECT 2912.805 3290.025 2914.015 3291.115 ;
        RECT 2912.805 3289.485 2913.325 3290.025 ;
        RECT 6.295 3286.935 6.815 3287.475 ;
        RECT 5.605 3285.845 6.815 3286.935 ;
        RECT 2912.805 3286.935 2913.325 3287.475 ;
        RECT 2912.805 3285.845 2914.015 3286.935 ;
        RECT 5.520 3285.675 6.900 3285.845 ;
        RECT 2909.960 3285.675 2910.420 3285.845 ;
        RECT 2912.720 3285.675 2914.100 3285.845 ;
        RECT 5.605 3284.585 6.815 3285.675 ;
        RECT 6.295 3284.045 6.815 3284.585 ;
        RECT 2910.045 3284.510 2910.335 3285.675 ;
        RECT 2912.805 3284.585 2914.015 3285.675 ;
        RECT 2912.805 3284.045 2913.325 3284.585 ;
        RECT 6.295 3281.495 6.815 3282.035 ;
        RECT 5.605 3280.405 6.815 3281.495 ;
        RECT 2912.805 3281.495 2913.325 3282.035 ;
        RECT 2912.805 3280.405 2914.015 3281.495 ;
        RECT 5.520 3280.235 6.900 3280.405 ;
        RECT 2909.960 3280.235 2910.420 3280.405 ;
        RECT 2912.720 3280.235 2914.100 3280.405 ;
        RECT 5.605 3279.145 6.815 3280.235 ;
        RECT 6.295 3278.605 6.815 3279.145 ;
        RECT 2910.045 3279.070 2910.335 3280.235 ;
        RECT 2912.805 3279.145 2914.015 3280.235 ;
        RECT 2912.805 3278.605 2913.325 3279.145 ;
        RECT 6.295 3276.055 6.815 3276.595 ;
        RECT 5.605 3274.965 6.815 3276.055 ;
        RECT 2912.805 3276.055 2913.325 3276.595 ;
        RECT 2912.805 3274.965 2914.015 3276.055 ;
        RECT 5.520 3274.795 6.900 3274.965 ;
        RECT 2909.960 3274.795 2910.420 3274.965 ;
        RECT 2912.720 3274.795 2914.100 3274.965 ;
        RECT 5.605 3273.705 6.815 3274.795 ;
        RECT 6.295 3273.165 6.815 3273.705 ;
        RECT 2910.045 3273.630 2910.335 3274.795 ;
        RECT 2912.805 3273.705 2914.015 3274.795 ;
        RECT 2912.805 3273.165 2913.325 3273.705 ;
        RECT 6.295 3270.615 6.815 3271.155 ;
        RECT 5.605 3269.525 6.815 3270.615 ;
        RECT 2912.805 3270.615 2913.325 3271.155 ;
        RECT 2912.805 3269.525 2914.015 3270.615 ;
        RECT 5.520 3269.355 6.900 3269.525 ;
        RECT 2909.960 3269.355 2910.420 3269.525 ;
        RECT 2912.720 3269.355 2914.100 3269.525 ;
        RECT 5.605 3268.265 6.815 3269.355 ;
        RECT 6.295 3267.725 6.815 3268.265 ;
        RECT 2910.045 3268.190 2910.335 3269.355 ;
        RECT 2912.805 3268.265 2914.015 3269.355 ;
        RECT 2912.805 3267.725 2913.325 3268.265 ;
        RECT 6.295 3265.175 6.815 3265.715 ;
        RECT 5.605 3264.085 6.815 3265.175 ;
        RECT 2912.805 3265.175 2913.325 3265.715 ;
        RECT 2912.805 3264.085 2914.015 3265.175 ;
        RECT 5.520 3263.915 6.900 3264.085 ;
        RECT 2909.960 3263.915 2910.420 3264.085 ;
        RECT 2912.720 3263.915 2914.100 3264.085 ;
        RECT 5.605 3262.825 6.815 3263.915 ;
        RECT 6.295 3262.285 6.815 3262.825 ;
        RECT 2910.045 3262.750 2910.335 3263.915 ;
        RECT 2912.805 3262.825 2914.015 3263.915 ;
        RECT 2912.805 3262.285 2913.325 3262.825 ;
        RECT 6.295 3259.735 6.815 3260.275 ;
        RECT 5.605 3258.645 6.815 3259.735 ;
        RECT 2912.805 3259.735 2913.325 3260.275 ;
        RECT 2912.805 3258.645 2914.015 3259.735 ;
        RECT 5.520 3258.475 6.900 3258.645 ;
        RECT 2909.960 3258.475 2910.420 3258.645 ;
        RECT 2912.720 3258.475 2914.100 3258.645 ;
        RECT 5.605 3257.385 6.815 3258.475 ;
        RECT 6.295 3256.845 6.815 3257.385 ;
        RECT 2910.045 3257.310 2910.335 3258.475 ;
        RECT 2912.805 3257.385 2914.015 3258.475 ;
        RECT 2912.805 3256.845 2913.325 3257.385 ;
        RECT 6.295 3254.295 6.815 3254.835 ;
        RECT 5.605 3253.205 6.815 3254.295 ;
        RECT 2912.805 3254.295 2913.325 3254.835 ;
        RECT 2912.805 3253.205 2914.015 3254.295 ;
        RECT 5.520 3253.035 6.900 3253.205 ;
        RECT 2909.960 3253.035 2910.420 3253.205 ;
        RECT 2912.720 3253.035 2914.100 3253.205 ;
        RECT 5.605 3251.945 6.815 3253.035 ;
        RECT 6.295 3251.405 6.815 3251.945 ;
        RECT 2910.045 3251.870 2910.335 3253.035 ;
        RECT 2912.805 3251.945 2914.015 3253.035 ;
        RECT 2912.805 3251.405 2913.325 3251.945 ;
        RECT 6.295 3248.855 6.815 3249.395 ;
        RECT 5.605 3247.765 6.815 3248.855 ;
        RECT 2912.805 3248.855 2913.325 3249.395 ;
        RECT 2912.805 3247.765 2914.015 3248.855 ;
        RECT 5.520 3247.595 6.900 3247.765 ;
        RECT 2909.960 3247.595 2910.420 3247.765 ;
        RECT 2912.720 3247.595 2914.100 3247.765 ;
        RECT 5.605 3246.505 6.815 3247.595 ;
        RECT 6.295 3245.965 6.815 3246.505 ;
        RECT 2910.045 3246.430 2910.335 3247.595 ;
        RECT 2912.805 3246.505 2914.015 3247.595 ;
        RECT 2912.805 3245.965 2913.325 3246.505 ;
        RECT 6.295 3243.415 6.815 3243.955 ;
        RECT 5.605 3242.325 6.815 3243.415 ;
        RECT 2912.805 3243.415 2913.325 3243.955 ;
        RECT 2912.805 3242.325 2914.015 3243.415 ;
        RECT 5.520 3242.155 6.900 3242.325 ;
        RECT 2909.960 3242.155 2910.420 3242.325 ;
        RECT 2912.720 3242.155 2914.100 3242.325 ;
        RECT 5.605 3241.065 6.815 3242.155 ;
        RECT 6.295 3240.525 6.815 3241.065 ;
        RECT 2910.045 3240.990 2910.335 3242.155 ;
        RECT 2912.805 3241.065 2914.015 3242.155 ;
        RECT 2912.805 3240.525 2913.325 3241.065 ;
        RECT 6.295 3237.975 6.815 3238.515 ;
        RECT 5.605 3236.885 6.815 3237.975 ;
        RECT 2912.805 3237.975 2913.325 3238.515 ;
        RECT 2912.805 3236.885 2914.015 3237.975 ;
        RECT 5.520 3236.715 6.900 3236.885 ;
        RECT 2909.960 3236.715 2910.420 3236.885 ;
        RECT 2912.720 3236.715 2914.100 3236.885 ;
        RECT 5.605 3235.625 6.815 3236.715 ;
        RECT 6.295 3235.085 6.815 3235.625 ;
        RECT 2910.045 3235.550 2910.335 3236.715 ;
        RECT 2912.805 3235.625 2914.015 3236.715 ;
        RECT 2912.805 3235.085 2913.325 3235.625 ;
        RECT 6.295 3232.535 6.815 3233.075 ;
        RECT 5.605 3231.445 6.815 3232.535 ;
        RECT 2912.805 3232.535 2913.325 3233.075 ;
        RECT 2912.805 3231.445 2914.015 3232.535 ;
        RECT 5.520 3231.275 6.900 3231.445 ;
        RECT 2909.960 3231.275 2910.420 3231.445 ;
        RECT 2912.720 3231.275 2914.100 3231.445 ;
        RECT 5.605 3230.185 6.815 3231.275 ;
        RECT 6.295 3229.645 6.815 3230.185 ;
        RECT 2910.045 3230.110 2910.335 3231.275 ;
        RECT 2912.805 3230.185 2914.015 3231.275 ;
        RECT 2912.805 3229.645 2913.325 3230.185 ;
        RECT 6.295 3227.095 6.815 3227.635 ;
        RECT 5.605 3226.005 6.815 3227.095 ;
        RECT 2912.805 3227.095 2913.325 3227.635 ;
        RECT 2912.805 3226.005 2914.015 3227.095 ;
        RECT 5.520 3225.835 6.900 3226.005 ;
        RECT 8.740 3225.835 10.120 3226.005 ;
        RECT 2909.960 3225.835 2910.420 3226.005 ;
        RECT 2912.720 3225.835 2914.100 3226.005 ;
        RECT 5.605 3224.745 6.815 3225.835 ;
        RECT 9.015 3225.110 9.345 3225.835 ;
        RECT 6.295 3224.205 6.815 3224.745 ;
        RECT 2910.045 3224.670 2910.335 3225.835 ;
        RECT 2912.805 3224.745 2914.015 3225.835 ;
        RECT 2912.805 3224.205 2913.325 3224.745 ;
        RECT 6.295 3221.655 6.815 3222.195 ;
        RECT 5.605 3220.565 6.815 3221.655 ;
        RECT 2912.805 3221.655 2913.325 3222.195 ;
        RECT 2912.805 3220.565 2914.015 3221.655 ;
        RECT 5.520 3220.395 6.900 3220.565 ;
        RECT 2909.960 3220.395 2910.420 3220.565 ;
        RECT 2912.720 3220.395 2914.100 3220.565 ;
        RECT 5.605 3219.305 6.815 3220.395 ;
        RECT 6.295 3218.765 6.815 3219.305 ;
        RECT 2910.045 3219.230 2910.335 3220.395 ;
        RECT 2912.805 3219.305 2914.015 3220.395 ;
        RECT 2912.805 3218.765 2913.325 3219.305 ;
        RECT 6.295 3216.215 6.815 3216.755 ;
        RECT 5.605 3215.125 6.815 3216.215 ;
        RECT 2912.805 3216.215 2913.325 3216.755 ;
        RECT 2912.805 3215.125 2914.015 3216.215 ;
        RECT 5.520 3214.955 6.900 3215.125 ;
        RECT 2909.960 3214.955 2910.420 3215.125 ;
        RECT 2912.720 3214.955 2914.100 3215.125 ;
        RECT 5.605 3213.865 6.815 3214.955 ;
        RECT 6.295 3213.325 6.815 3213.865 ;
        RECT 2910.045 3213.790 2910.335 3214.955 ;
        RECT 2912.805 3213.865 2914.015 3214.955 ;
        RECT 2912.805 3213.325 2913.325 3213.865 ;
        RECT 6.295 3210.775 6.815 3211.315 ;
        RECT 5.605 3209.685 6.815 3210.775 ;
        RECT 2912.805 3210.775 2913.325 3211.315 ;
        RECT 2912.805 3209.685 2914.015 3210.775 ;
        RECT 5.520 3209.515 6.900 3209.685 ;
        RECT 2909.960 3209.515 2910.420 3209.685 ;
        RECT 2912.720 3209.515 2914.100 3209.685 ;
        RECT 5.605 3208.425 6.815 3209.515 ;
        RECT 6.295 3207.885 6.815 3208.425 ;
        RECT 2910.045 3208.350 2910.335 3209.515 ;
        RECT 2912.805 3208.425 2914.015 3209.515 ;
        RECT 2912.805 3207.885 2913.325 3208.425 ;
        RECT 6.295 3205.335 6.815 3205.875 ;
        RECT 5.605 3204.245 6.815 3205.335 ;
        RECT 2912.805 3205.335 2913.325 3205.875 ;
        RECT 2912.805 3204.245 2914.015 3205.335 ;
        RECT 5.520 3204.075 6.900 3204.245 ;
        RECT 2909.960 3204.075 2911.800 3204.245 ;
        RECT 2912.720 3204.075 2914.100 3204.245 ;
        RECT 5.605 3202.985 6.815 3204.075 ;
        RECT 6.295 3202.445 6.815 3202.985 ;
        RECT 2910.045 3202.910 2910.335 3204.075 ;
        RECT 2910.695 3203.350 2911.025 3204.075 ;
        RECT 2912.805 3202.985 2914.015 3204.075 ;
        RECT 2912.805 3202.445 2913.325 3202.985 ;
        RECT 6.295 3199.895 6.815 3200.435 ;
        RECT 5.605 3198.805 6.815 3199.895 ;
        RECT 2912.805 3199.895 2913.325 3200.435 ;
        RECT 2912.805 3198.805 2914.015 3199.895 ;
        RECT 5.520 3198.635 6.900 3198.805 ;
        RECT 2909.960 3198.635 2910.420 3198.805 ;
        RECT 2912.720 3198.635 2914.100 3198.805 ;
        RECT 5.605 3197.545 6.815 3198.635 ;
        RECT 6.295 3197.005 6.815 3197.545 ;
        RECT 2910.045 3197.470 2910.335 3198.635 ;
        RECT 2912.805 3197.545 2914.015 3198.635 ;
        RECT 2912.805 3197.005 2913.325 3197.545 ;
        RECT 6.295 3194.455 6.815 3194.995 ;
        RECT 5.605 3193.365 6.815 3194.455 ;
        RECT 2912.805 3194.455 2913.325 3194.995 ;
        RECT 2912.805 3193.365 2914.015 3194.455 ;
        RECT 5.520 3193.195 6.900 3193.365 ;
        RECT 2909.960 3193.195 2910.420 3193.365 ;
        RECT 2912.720 3193.195 2914.100 3193.365 ;
        RECT 5.605 3192.105 6.815 3193.195 ;
        RECT 6.295 3191.565 6.815 3192.105 ;
        RECT 2910.045 3192.030 2910.335 3193.195 ;
        RECT 2912.805 3192.105 2914.015 3193.195 ;
        RECT 2912.805 3191.565 2913.325 3192.105 ;
        RECT 6.295 3189.015 6.815 3189.555 ;
        RECT 5.605 3187.925 6.815 3189.015 ;
        RECT 2912.805 3189.015 2913.325 3189.555 ;
        RECT 2912.805 3187.925 2914.015 3189.015 ;
        RECT 5.520 3187.755 6.900 3187.925 ;
        RECT 2909.960 3187.755 2910.420 3187.925 ;
        RECT 2912.720 3187.755 2914.100 3187.925 ;
        RECT 5.605 3186.665 6.815 3187.755 ;
        RECT 6.295 3186.125 6.815 3186.665 ;
        RECT 2910.045 3186.590 2910.335 3187.755 ;
        RECT 2912.805 3186.665 2914.015 3187.755 ;
        RECT 2912.805 3186.125 2913.325 3186.665 ;
        RECT 6.295 3183.575 6.815 3184.115 ;
        RECT 5.605 3182.485 6.815 3183.575 ;
        RECT 2912.805 3183.575 2913.325 3184.115 ;
        RECT 2912.805 3182.485 2914.015 3183.575 ;
        RECT 5.520 3182.315 6.900 3182.485 ;
        RECT 2909.960 3182.315 2910.420 3182.485 ;
        RECT 2912.720 3182.315 2914.100 3182.485 ;
        RECT 5.605 3181.225 6.815 3182.315 ;
        RECT 6.295 3180.685 6.815 3181.225 ;
        RECT 2910.045 3181.150 2910.335 3182.315 ;
        RECT 2912.805 3181.225 2914.015 3182.315 ;
        RECT 2912.805 3180.685 2913.325 3181.225 ;
        RECT 6.295 3178.135 6.815 3178.675 ;
        RECT 5.605 3177.045 6.815 3178.135 ;
        RECT 2912.805 3178.135 2913.325 3178.675 ;
        RECT 2912.805 3177.045 2914.015 3178.135 ;
        RECT 5.520 3176.875 6.900 3177.045 ;
        RECT 2909.960 3176.875 2910.420 3177.045 ;
        RECT 2912.720 3176.875 2914.100 3177.045 ;
        RECT 5.605 3175.785 6.815 3176.875 ;
        RECT 6.295 3175.245 6.815 3175.785 ;
        RECT 2910.045 3175.710 2910.335 3176.875 ;
        RECT 2912.805 3175.785 2914.015 3176.875 ;
        RECT 2912.805 3175.245 2913.325 3175.785 ;
        RECT 6.295 3172.695 6.815 3173.235 ;
        RECT 5.605 3171.605 6.815 3172.695 ;
        RECT 2912.805 3172.695 2913.325 3173.235 ;
        RECT 2912.805 3171.605 2914.015 3172.695 ;
        RECT 5.520 3171.435 6.900 3171.605 ;
        RECT 2909.960 3171.435 2910.420 3171.605 ;
        RECT 2912.720 3171.435 2914.100 3171.605 ;
        RECT 5.605 3170.345 6.815 3171.435 ;
        RECT 6.295 3169.805 6.815 3170.345 ;
        RECT 2910.045 3170.270 2910.335 3171.435 ;
        RECT 2912.805 3170.345 2914.015 3171.435 ;
        RECT 2912.805 3169.805 2913.325 3170.345 ;
        RECT 6.295 3167.255 6.815 3167.795 ;
        RECT 5.605 3166.165 6.815 3167.255 ;
        RECT 2912.805 3167.255 2913.325 3167.795 ;
        RECT 2912.805 3166.165 2914.015 3167.255 ;
        RECT 5.520 3165.995 6.900 3166.165 ;
        RECT 2909.960 3165.995 2910.420 3166.165 ;
        RECT 2912.720 3165.995 2914.100 3166.165 ;
        RECT 5.605 3164.905 6.815 3165.995 ;
        RECT 6.295 3164.365 6.815 3164.905 ;
        RECT 2910.045 3164.830 2910.335 3165.995 ;
        RECT 2912.805 3164.905 2914.015 3165.995 ;
        RECT 2912.805 3164.365 2913.325 3164.905 ;
        RECT 6.295 3161.815 6.815 3162.355 ;
        RECT 5.605 3160.725 6.815 3161.815 ;
        RECT 2912.805 3161.815 2913.325 3162.355 ;
        RECT 2912.805 3160.725 2914.015 3161.815 ;
        RECT 5.520 3160.555 6.900 3160.725 ;
        RECT 2909.960 3160.555 2910.420 3160.725 ;
        RECT 2912.720 3160.555 2914.100 3160.725 ;
        RECT 5.605 3159.465 6.815 3160.555 ;
        RECT 6.295 3158.925 6.815 3159.465 ;
        RECT 2910.045 3159.390 2910.335 3160.555 ;
        RECT 2912.805 3159.465 2914.015 3160.555 ;
        RECT 2912.805 3158.925 2913.325 3159.465 ;
        RECT 6.295 3156.375 6.815 3156.915 ;
        RECT 5.605 3155.285 6.815 3156.375 ;
        RECT 2912.805 3156.375 2913.325 3156.915 ;
        RECT 2912.805 3155.285 2914.015 3156.375 ;
        RECT 5.520 3155.115 6.900 3155.285 ;
        RECT 2909.960 3155.115 2910.420 3155.285 ;
        RECT 2912.720 3155.115 2914.100 3155.285 ;
        RECT 5.605 3154.025 6.815 3155.115 ;
        RECT 6.295 3153.485 6.815 3154.025 ;
        RECT 2910.045 3153.950 2910.335 3155.115 ;
        RECT 2912.805 3154.025 2914.015 3155.115 ;
        RECT 2912.805 3153.485 2913.325 3154.025 ;
        RECT 6.295 3150.935 6.815 3151.475 ;
        RECT 5.605 3149.845 6.815 3150.935 ;
        RECT 2912.805 3150.935 2913.325 3151.475 ;
        RECT 2912.805 3149.845 2914.015 3150.935 ;
        RECT 5.520 3149.675 6.900 3149.845 ;
        RECT 2909.960 3149.675 2910.420 3149.845 ;
        RECT 2912.720 3149.675 2914.100 3149.845 ;
        RECT 5.605 3148.585 6.815 3149.675 ;
        RECT 6.295 3148.045 6.815 3148.585 ;
        RECT 2910.045 3148.510 2910.335 3149.675 ;
        RECT 2912.805 3148.585 2914.015 3149.675 ;
        RECT 2912.805 3148.045 2913.325 3148.585 ;
        RECT 6.295 3145.495 6.815 3146.035 ;
        RECT 5.605 3144.405 6.815 3145.495 ;
        RECT 2912.805 3145.495 2913.325 3146.035 ;
        RECT 2912.805 3144.405 2914.015 3145.495 ;
        RECT 5.520 3144.235 6.900 3144.405 ;
        RECT 2909.960 3144.235 2910.420 3144.405 ;
        RECT 2912.720 3144.235 2914.100 3144.405 ;
        RECT 5.605 3143.145 6.815 3144.235 ;
        RECT 6.295 3142.605 6.815 3143.145 ;
        RECT 2910.045 3143.070 2910.335 3144.235 ;
        RECT 2912.805 3143.145 2914.015 3144.235 ;
        RECT 2912.805 3142.605 2913.325 3143.145 ;
        RECT 6.295 3140.055 6.815 3140.595 ;
        RECT 5.605 3138.965 6.815 3140.055 ;
        RECT 2912.805 3140.055 2913.325 3140.595 ;
        RECT 2912.805 3138.965 2914.015 3140.055 ;
        RECT 5.520 3138.795 6.900 3138.965 ;
        RECT 2909.960 3138.795 2910.420 3138.965 ;
        RECT 2912.720 3138.795 2914.100 3138.965 ;
        RECT 5.605 3137.705 6.815 3138.795 ;
        RECT 6.295 3137.165 6.815 3137.705 ;
        RECT 2910.045 3137.630 2910.335 3138.795 ;
        RECT 2912.805 3137.705 2914.015 3138.795 ;
        RECT 2912.805 3137.165 2913.325 3137.705 ;
        RECT 6.295 3134.615 6.815 3135.155 ;
        RECT 5.605 3133.525 6.815 3134.615 ;
        RECT 2912.805 3134.615 2913.325 3135.155 ;
        RECT 2912.805 3133.525 2914.015 3134.615 ;
        RECT 5.520 3133.355 6.900 3133.525 ;
        RECT 2909.960 3133.355 2910.420 3133.525 ;
        RECT 2912.720 3133.355 2914.100 3133.525 ;
        RECT 5.605 3132.265 6.815 3133.355 ;
        RECT 6.295 3131.725 6.815 3132.265 ;
        RECT 2910.045 3132.190 2910.335 3133.355 ;
        RECT 2912.805 3132.265 2914.015 3133.355 ;
        RECT 2912.805 3131.725 2913.325 3132.265 ;
        RECT 6.295 3129.175 6.815 3129.715 ;
        RECT 5.605 3128.085 6.815 3129.175 ;
        RECT 2912.805 3129.175 2913.325 3129.715 ;
        RECT 2912.805 3128.085 2914.015 3129.175 ;
        RECT 5.520 3127.915 6.900 3128.085 ;
        RECT 2909.960 3127.915 2910.420 3128.085 ;
        RECT 2912.720 3127.915 2914.100 3128.085 ;
        RECT 5.605 3126.825 6.815 3127.915 ;
        RECT 6.295 3126.285 6.815 3126.825 ;
        RECT 2910.045 3126.750 2910.335 3127.915 ;
        RECT 2912.805 3126.825 2914.015 3127.915 ;
        RECT 2912.805 3126.285 2913.325 3126.825 ;
        RECT 6.295 3123.735 6.815 3124.275 ;
        RECT 5.605 3122.645 6.815 3123.735 ;
        RECT 2912.805 3123.735 2913.325 3124.275 ;
        RECT 2912.805 3122.645 2914.015 3123.735 ;
        RECT 5.520 3122.475 6.900 3122.645 ;
        RECT 2909.960 3122.475 2910.420 3122.645 ;
        RECT 2912.720 3122.475 2914.100 3122.645 ;
        RECT 5.605 3121.385 6.815 3122.475 ;
        RECT 6.295 3120.845 6.815 3121.385 ;
        RECT 2910.045 3121.310 2910.335 3122.475 ;
        RECT 2912.805 3121.385 2914.015 3122.475 ;
        RECT 2912.805 3120.845 2913.325 3121.385 ;
        RECT 6.295 3118.295 6.815 3118.835 ;
        RECT 5.605 3117.205 6.815 3118.295 ;
        RECT 2912.805 3118.295 2913.325 3118.835 ;
        RECT 2912.805 3117.205 2914.015 3118.295 ;
        RECT 5.520 3117.035 6.900 3117.205 ;
        RECT 2909.960 3117.035 2910.420 3117.205 ;
        RECT 2912.720 3117.035 2914.100 3117.205 ;
        RECT 5.605 3115.945 6.815 3117.035 ;
        RECT 6.295 3115.405 6.815 3115.945 ;
        RECT 2910.045 3115.870 2910.335 3117.035 ;
        RECT 2912.805 3115.945 2914.015 3117.035 ;
        RECT 2912.805 3115.405 2913.325 3115.945 ;
        RECT 6.295 3112.855 6.815 3113.395 ;
        RECT 5.605 3111.765 6.815 3112.855 ;
        RECT 2912.805 3112.855 2913.325 3113.395 ;
        RECT 2912.805 3111.765 2914.015 3112.855 ;
        RECT 5.520 3111.595 6.900 3111.765 ;
        RECT 2909.960 3111.595 2910.420 3111.765 ;
        RECT 2912.720 3111.595 2914.100 3111.765 ;
        RECT 5.605 3110.505 6.815 3111.595 ;
        RECT 6.295 3109.965 6.815 3110.505 ;
        RECT 2910.045 3110.430 2910.335 3111.595 ;
        RECT 2912.805 3110.505 2914.015 3111.595 ;
        RECT 2912.805 3109.965 2913.325 3110.505 ;
        RECT 6.295 3107.415 6.815 3107.955 ;
        RECT 5.605 3106.325 6.815 3107.415 ;
        RECT 2912.805 3107.415 2913.325 3107.955 ;
        RECT 2912.805 3106.325 2914.015 3107.415 ;
        RECT 5.520 3106.155 6.900 3106.325 ;
        RECT 2909.960 3106.155 2910.420 3106.325 ;
        RECT 2912.720 3106.155 2914.100 3106.325 ;
        RECT 5.605 3105.065 6.815 3106.155 ;
        RECT 6.295 3104.525 6.815 3105.065 ;
        RECT 2910.045 3104.990 2910.335 3106.155 ;
        RECT 2912.805 3105.065 2914.015 3106.155 ;
        RECT 2912.805 3104.525 2913.325 3105.065 ;
        RECT 6.295 3101.975 6.815 3102.515 ;
        RECT 5.605 3100.885 6.815 3101.975 ;
        RECT 2912.805 3101.975 2913.325 3102.515 ;
        RECT 2912.805 3100.885 2914.015 3101.975 ;
        RECT 5.520 3100.715 6.900 3100.885 ;
        RECT 2909.960 3100.715 2910.420 3100.885 ;
        RECT 2912.720 3100.715 2914.100 3100.885 ;
        RECT 5.605 3099.625 6.815 3100.715 ;
        RECT 6.295 3099.085 6.815 3099.625 ;
        RECT 2910.045 3099.550 2910.335 3100.715 ;
        RECT 2912.805 3099.625 2914.015 3100.715 ;
        RECT 2912.805 3099.085 2913.325 3099.625 ;
        RECT 6.295 3096.535 6.815 3097.075 ;
        RECT 5.605 3095.445 6.815 3096.535 ;
        RECT 2912.805 3096.535 2913.325 3097.075 ;
        RECT 2909.315 3095.445 2909.645 3096.170 ;
        RECT 2912.805 3095.445 2914.015 3096.535 ;
        RECT 5.520 3095.275 6.900 3095.445 ;
        RECT 2909.040 3095.275 2910.420 3095.445 ;
        RECT 2912.720 3095.275 2914.100 3095.445 ;
        RECT 5.605 3094.185 6.815 3095.275 ;
        RECT 6.295 3093.645 6.815 3094.185 ;
        RECT 2910.045 3094.110 2910.335 3095.275 ;
        RECT 2912.805 3094.185 2914.015 3095.275 ;
        RECT 2912.805 3093.645 2913.325 3094.185 ;
        RECT 6.295 3091.095 6.815 3091.635 ;
        RECT 5.605 3090.005 6.815 3091.095 ;
        RECT 2912.805 3091.095 2913.325 3091.635 ;
        RECT 2912.805 3090.005 2914.015 3091.095 ;
        RECT 5.520 3089.835 6.900 3090.005 ;
        RECT 2909.960 3089.835 2910.420 3090.005 ;
        RECT 2912.720 3089.835 2914.100 3090.005 ;
        RECT 5.605 3088.745 6.815 3089.835 ;
        RECT 6.295 3088.205 6.815 3088.745 ;
        RECT 2910.045 3088.670 2910.335 3089.835 ;
        RECT 2912.805 3088.745 2914.015 3089.835 ;
        RECT 2912.805 3088.205 2913.325 3088.745 ;
        RECT 6.295 3085.655 6.815 3086.195 ;
        RECT 5.605 3084.565 6.815 3085.655 ;
        RECT 2912.805 3085.655 2913.325 3086.195 ;
        RECT 2912.805 3084.565 2914.015 3085.655 ;
        RECT 5.520 3084.395 6.900 3084.565 ;
        RECT 2909.960 3084.395 2910.420 3084.565 ;
        RECT 2912.720 3084.395 2914.100 3084.565 ;
        RECT 5.605 3083.305 6.815 3084.395 ;
        RECT 6.295 3082.765 6.815 3083.305 ;
        RECT 2910.045 3083.230 2910.335 3084.395 ;
        RECT 2912.805 3083.305 2914.015 3084.395 ;
        RECT 2912.805 3082.765 2913.325 3083.305 ;
        RECT 6.295 3080.215 6.815 3080.755 ;
        RECT 5.605 3079.125 6.815 3080.215 ;
        RECT 2912.805 3080.215 2913.325 3080.755 ;
        RECT 2912.805 3079.125 2914.015 3080.215 ;
        RECT 5.520 3078.955 6.900 3079.125 ;
        RECT 2909.960 3078.955 2910.420 3079.125 ;
        RECT 2912.720 3078.955 2914.100 3079.125 ;
        RECT 5.605 3077.865 6.815 3078.955 ;
        RECT 6.295 3077.325 6.815 3077.865 ;
        RECT 2910.045 3077.790 2910.335 3078.955 ;
        RECT 2912.805 3077.865 2914.015 3078.955 ;
        RECT 2912.805 3077.325 2913.325 3077.865 ;
        RECT 6.295 3074.775 6.815 3075.315 ;
        RECT 5.605 3073.685 6.815 3074.775 ;
        RECT 2912.805 3074.775 2913.325 3075.315 ;
        RECT 2912.805 3073.685 2914.015 3074.775 ;
        RECT 5.520 3073.515 6.900 3073.685 ;
        RECT 2909.960 3073.515 2910.420 3073.685 ;
        RECT 2912.720 3073.515 2914.100 3073.685 ;
        RECT 5.605 3072.425 6.815 3073.515 ;
        RECT 6.295 3071.885 6.815 3072.425 ;
        RECT 2910.045 3072.350 2910.335 3073.515 ;
        RECT 2912.805 3072.425 2914.015 3073.515 ;
        RECT 2912.805 3071.885 2913.325 3072.425 ;
        RECT 6.295 3069.335 6.815 3069.875 ;
        RECT 5.605 3068.245 6.815 3069.335 ;
        RECT 2912.805 3069.335 2913.325 3069.875 ;
        RECT 2912.805 3068.245 2914.015 3069.335 ;
        RECT 5.520 3068.075 6.900 3068.245 ;
        RECT 2909.960 3068.075 2910.420 3068.245 ;
        RECT 2912.720 3068.075 2914.100 3068.245 ;
        RECT 5.605 3066.985 6.815 3068.075 ;
        RECT 6.295 3066.445 6.815 3066.985 ;
        RECT 2910.045 3066.910 2910.335 3068.075 ;
        RECT 2912.805 3066.985 2914.015 3068.075 ;
        RECT 2912.805 3066.445 2913.325 3066.985 ;
        RECT 6.295 3063.895 6.815 3064.435 ;
        RECT 5.605 3062.805 6.815 3063.895 ;
        RECT 2912.805 3063.895 2913.325 3064.435 ;
        RECT 2912.805 3062.805 2914.015 3063.895 ;
        RECT 5.520 3062.635 6.900 3062.805 ;
        RECT 2909.960 3062.635 2910.420 3062.805 ;
        RECT 2912.720 3062.635 2914.100 3062.805 ;
        RECT 5.605 3061.545 6.815 3062.635 ;
        RECT 6.295 3061.005 6.815 3061.545 ;
        RECT 2910.045 3061.470 2910.335 3062.635 ;
        RECT 2912.805 3061.545 2914.015 3062.635 ;
        RECT 2912.805 3061.005 2913.325 3061.545 ;
        RECT 6.295 3058.455 6.815 3058.995 ;
        RECT 5.605 3057.365 6.815 3058.455 ;
        RECT 2912.805 3058.455 2913.325 3058.995 ;
        RECT 2912.805 3057.365 2914.015 3058.455 ;
        RECT 5.520 3057.195 6.900 3057.365 ;
        RECT 2909.960 3057.195 2910.420 3057.365 ;
        RECT 2912.720 3057.195 2914.100 3057.365 ;
        RECT 5.605 3056.105 6.815 3057.195 ;
        RECT 6.295 3055.565 6.815 3056.105 ;
        RECT 2910.045 3056.030 2910.335 3057.195 ;
        RECT 2912.805 3056.105 2914.015 3057.195 ;
        RECT 2912.805 3055.565 2913.325 3056.105 ;
        RECT 6.295 3053.015 6.815 3053.555 ;
        RECT 5.605 3051.925 6.815 3053.015 ;
        RECT 2912.805 3053.015 2913.325 3053.555 ;
        RECT 2912.805 3051.925 2914.015 3053.015 ;
        RECT 5.520 3051.755 6.900 3051.925 ;
        RECT 2909.960 3051.755 2910.420 3051.925 ;
        RECT 2912.720 3051.755 2914.100 3051.925 ;
        RECT 5.605 3050.665 6.815 3051.755 ;
        RECT 6.295 3050.125 6.815 3050.665 ;
        RECT 2910.045 3050.590 2910.335 3051.755 ;
        RECT 2912.805 3050.665 2914.015 3051.755 ;
        RECT 2912.805 3050.125 2913.325 3050.665 ;
        RECT 6.295 3047.575 6.815 3048.115 ;
        RECT 5.605 3046.485 6.815 3047.575 ;
        RECT 2912.805 3047.575 2913.325 3048.115 ;
        RECT 2912.805 3046.485 2914.015 3047.575 ;
        RECT 5.520 3046.315 6.900 3046.485 ;
        RECT 2909.960 3046.315 2910.420 3046.485 ;
        RECT 2912.720 3046.315 2914.100 3046.485 ;
        RECT 5.605 3045.225 6.815 3046.315 ;
        RECT 6.295 3044.685 6.815 3045.225 ;
        RECT 2910.045 3045.150 2910.335 3046.315 ;
        RECT 2912.805 3045.225 2914.015 3046.315 ;
        RECT 2912.805 3044.685 2913.325 3045.225 ;
        RECT 6.295 3042.135 6.815 3042.675 ;
        RECT 5.605 3041.045 6.815 3042.135 ;
        RECT 2912.805 3042.135 2913.325 3042.675 ;
        RECT 2912.805 3041.045 2914.015 3042.135 ;
        RECT 5.520 3040.875 6.900 3041.045 ;
        RECT 2909.960 3040.875 2910.420 3041.045 ;
        RECT 2912.720 3040.875 2914.100 3041.045 ;
        RECT 5.605 3039.785 6.815 3040.875 ;
        RECT 6.295 3039.245 6.815 3039.785 ;
        RECT 2910.045 3039.710 2910.335 3040.875 ;
        RECT 2912.805 3039.785 2914.015 3040.875 ;
        RECT 2912.805 3039.245 2913.325 3039.785 ;
        RECT 6.295 3036.695 6.815 3037.235 ;
        RECT 5.605 3035.605 6.815 3036.695 ;
        RECT 2912.805 3036.695 2913.325 3037.235 ;
        RECT 2912.805 3035.605 2914.015 3036.695 ;
        RECT 5.520 3035.435 6.900 3035.605 ;
        RECT 2909.960 3035.435 2910.420 3035.605 ;
        RECT 2912.720 3035.435 2914.100 3035.605 ;
        RECT 5.605 3034.345 6.815 3035.435 ;
        RECT 6.295 3033.805 6.815 3034.345 ;
        RECT 2910.045 3034.270 2910.335 3035.435 ;
        RECT 2912.805 3034.345 2914.015 3035.435 ;
        RECT 2912.805 3033.805 2913.325 3034.345 ;
        RECT 6.295 3031.255 6.815 3031.795 ;
        RECT 5.605 3030.165 6.815 3031.255 ;
        RECT 2912.805 3031.255 2913.325 3031.795 ;
        RECT 2912.805 3030.165 2914.015 3031.255 ;
        RECT 5.520 3029.995 6.900 3030.165 ;
        RECT 2909.960 3029.995 2910.420 3030.165 ;
        RECT 2912.720 3029.995 2914.100 3030.165 ;
        RECT 5.605 3028.905 6.815 3029.995 ;
        RECT 6.295 3028.365 6.815 3028.905 ;
        RECT 2910.045 3028.830 2910.335 3029.995 ;
        RECT 2912.805 3028.905 2914.015 3029.995 ;
        RECT 2912.805 3028.365 2913.325 3028.905 ;
        RECT 6.295 3025.815 6.815 3026.355 ;
        RECT 5.605 3024.725 6.815 3025.815 ;
        RECT 2912.805 3025.815 2913.325 3026.355 ;
        RECT 2912.805 3024.725 2914.015 3025.815 ;
        RECT 5.520 3024.555 6.900 3024.725 ;
        RECT 2909.960 3024.555 2910.420 3024.725 ;
        RECT 2912.720 3024.555 2914.100 3024.725 ;
        RECT 5.605 3023.465 6.815 3024.555 ;
        RECT 6.295 3022.925 6.815 3023.465 ;
        RECT 2910.045 3023.390 2910.335 3024.555 ;
        RECT 2912.805 3023.465 2914.015 3024.555 ;
        RECT 2912.805 3022.925 2913.325 3023.465 ;
        RECT 6.295 3020.375 6.815 3020.915 ;
        RECT 5.605 3019.285 6.815 3020.375 ;
        RECT 2912.805 3020.375 2913.325 3020.915 ;
        RECT 2912.805 3019.285 2914.015 3020.375 ;
        RECT 5.520 3019.115 6.900 3019.285 ;
        RECT 2909.960 3019.115 2910.420 3019.285 ;
        RECT 2912.720 3019.115 2914.100 3019.285 ;
        RECT 5.605 3018.025 6.815 3019.115 ;
        RECT 6.295 3017.485 6.815 3018.025 ;
        RECT 2910.045 3017.950 2910.335 3019.115 ;
        RECT 2912.805 3018.025 2914.015 3019.115 ;
        RECT 2912.805 3017.485 2913.325 3018.025 ;
        RECT 6.295 3014.935 6.815 3015.475 ;
        RECT 5.605 3013.845 6.815 3014.935 ;
        RECT 2912.805 3014.935 2913.325 3015.475 ;
        RECT 2912.805 3013.845 2914.015 3014.935 ;
        RECT 5.520 3013.675 6.900 3013.845 ;
        RECT 8.740 3013.675 10.120 3013.845 ;
        RECT 2909.960 3013.675 2910.420 3013.845 ;
        RECT 2912.720 3013.675 2914.100 3013.845 ;
        RECT 5.605 3012.585 6.815 3013.675 ;
        RECT 9.015 3012.950 9.345 3013.675 ;
        RECT 6.295 3012.045 6.815 3012.585 ;
        RECT 2910.045 3012.510 2910.335 3013.675 ;
        RECT 2912.805 3012.585 2914.015 3013.675 ;
        RECT 2912.805 3012.045 2913.325 3012.585 ;
        RECT 6.295 3009.495 6.815 3010.035 ;
        RECT 5.605 3008.405 6.815 3009.495 ;
        RECT 2912.805 3009.495 2913.325 3010.035 ;
        RECT 2912.805 3008.405 2914.015 3009.495 ;
        RECT 5.520 3008.235 6.900 3008.405 ;
        RECT 2909.960 3008.235 2910.420 3008.405 ;
        RECT 2912.720 3008.235 2914.100 3008.405 ;
        RECT 5.605 3007.145 6.815 3008.235 ;
        RECT 6.295 3006.605 6.815 3007.145 ;
        RECT 2910.045 3007.070 2910.335 3008.235 ;
        RECT 2912.805 3007.145 2914.015 3008.235 ;
        RECT 2912.805 3006.605 2913.325 3007.145 ;
        RECT 6.295 3004.055 6.815 3004.595 ;
        RECT 5.605 3002.965 6.815 3004.055 ;
        RECT 2912.805 3004.055 2913.325 3004.595 ;
        RECT 2912.805 3002.965 2914.015 3004.055 ;
        RECT 5.520 3002.795 6.900 3002.965 ;
        RECT 2909.960 3002.795 2910.420 3002.965 ;
        RECT 2912.720 3002.795 2914.100 3002.965 ;
        RECT 5.605 3001.705 6.815 3002.795 ;
        RECT 6.295 3001.165 6.815 3001.705 ;
        RECT 2910.045 3001.630 2910.335 3002.795 ;
        RECT 2912.805 3001.705 2914.015 3002.795 ;
        RECT 2912.805 3001.165 2913.325 3001.705 ;
        RECT 6.295 2998.615 6.815 2999.155 ;
        RECT 5.605 2997.525 6.815 2998.615 ;
        RECT 2912.805 2998.615 2913.325 2999.155 ;
        RECT 2912.805 2997.525 2914.015 2998.615 ;
        RECT 5.520 2997.355 6.900 2997.525 ;
        RECT 2909.960 2997.355 2910.420 2997.525 ;
        RECT 2912.720 2997.355 2914.100 2997.525 ;
        RECT 5.605 2996.265 6.815 2997.355 ;
        RECT 6.295 2995.725 6.815 2996.265 ;
        RECT 2910.045 2996.190 2910.335 2997.355 ;
        RECT 2912.805 2996.265 2914.015 2997.355 ;
        RECT 2912.805 2995.725 2913.325 2996.265 ;
        RECT 6.295 2993.175 6.815 2993.715 ;
        RECT 5.605 2992.085 6.815 2993.175 ;
        RECT 2912.805 2993.175 2913.325 2993.715 ;
        RECT 2912.805 2992.085 2914.015 2993.175 ;
        RECT 5.520 2991.915 6.900 2992.085 ;
        RECT 2909.960 2991.915 2910.420 2992.085 ;
        RECT 2912.720 2991.915 2914.100 2992.085 ;
        RECT 5.605 2990.825 6.815 2991.915 ;
        RECT 6.295 2990.285 6.815 2990.825 ;
        RECT 2910.045 2990.750 2910.335 2991.915 ;
        RECT 2912.805 2990.825 2914.015 2991.915 ;
        RECT 2912.805 2990.285 2913.325 2990.825 ;
        RECT 6.295 2987.735 6.815 2988.275 ;
        RECT 5.605 2986.645 6.815 2987.735 ;
        RECT 2912.805 2987.735 2913.325 2988.275 ;
        RECT 2912.805 2986.645 2914.015 2987.735 ;
        RECT 5.520 2986.475 6.900 2986.645 ;
        RECT 2909.960 2986.475 2910.420 2986.645 ;
        RECT 2912.720 2986.475 2914.100 2986.645 ;
        RECT 5.605 2985.385 6.815 2986.475 ;
        RECT 6.295 2984.845 6.815 2985.385 ;
        RECT 2910.045 2985.310 2910.335 2986.475 ;
        RECT 2912.805 2985.385 2914.015 2986.475 ;
        RECT 2912.805 2984.845 2913.325 2985.385 ;
        RECT 6.295 2982.295 6.815 2982.835 ;
        RECT 5.605 2981.205 6.815 2982.295 ;
        RECT 2912.805 2982.295 2913.325 2982.835 ;
        RECT 2912.805 2981.205 2914.015 2982.295 ;
        RECT 5.520 2981.035 6.900 2981.205 ;
        RECT 2909.960 2981.035 2910.420 2981.205 ;
        RECT 2912.720 2981.035 2914.100 2981.205 ;
        RECT 5.605 2979.945 6.815 2981.035 ;
        RECT 6.295 2979.405 6.815 2979.945 ;
        RECT 2910.045 2979.870 2910.335 2981.035 ;
        RECT 2912.805 2979.945 2914.015 2981.035 ;
        RECT 2912.805 2979.405 2913.325 2979.945 ;
        RECT 6.295 2976.855 6.815 2977.395 ;
        RECT 5.605 2975.765 6.815 2976.855 ;
        RECT 2912.805 2976.855 2913.325 2977.395 ;
        RECT 2912.805 2975.765 2914.015 2976.855 ;
        RECT 5.520 2975.595 6.900 2975.765 ;
        RECT 2909.960 2975.595 2910.420 2975.765 ;
        RECT 2912.720 2975.595 2914.100 2975.765 ;
        RECT 5.605 2974.505 6.815 2975.595 ;
        RECT 6.295 2973.965 6.815 2974.505 ;
        RECT 2910.045 2974.430 2910.335 2975.595 ;
        RECT 2912.805 2974.505 2914.015 2975.595 ;
        RECT 2912.805 2973.965 2913.325 2974.505 ;
        RECT 6.295 2971.415 6.815 2971.955 ;
        RECT 5.605 2970.325 6.815 2971.415 ;
        RECT 2912.805 2971.415 2913.325 2971.955 ;
        RECT 9.015 2970.325 9.345 2971.050 ;
        RECT 2912.805 2970.325 2914.015 2971.415 ;
        RECT 5.520 2970.155 6.900 2970.325 ;
        RECT 8.740 2970.155 10.120 2970.325 ;
        RECT 2909.960 2970.155 2910.420 2970.325 ;
        RECT 2912.720 2970.155 2914.100 2970.325 ;
        RECT 5.605 2969.065 6.815 2970.155 ;
        RECT 6.295 2968.525 6.815 2969.065 ;
        RECT 2910.045 2968.990 2910.335 2970.155 ;
        RECT 2912.805 2969.065 2914.015 2970.155 ;
        RECT 2912.805 2968.525 2913.325 2969.065 ;
        RECT 6.295 2965.975 6.815 2966.515 ;
        RECT 5.605 2964.885 6.815 2965.975 ;
        RECT 2912.805 2965.975 2913.325 2966.515 ;
        RECT 2912.805 2964.885 2914.015 2965.975 ;
        RECT 5.520 2964.715 6.900 2964.885 ;
        RECT 2909.960 2964.715 2910.420 2964.885 ;
        RECT 2912.720 2964.715 2914.100 2964.885 ;
        RECT 5.605 2963.625 6.815 2964.715 ;
        RECT 6.295 2963.085 6.815 2963.625 ;
        RECT 2910.045 2963.550 2910.335 2964.715 ;
        RECT 2912.805 2963.625 2914.015 2964.715 ;
        RECT 2912.805 2963.085 2913.325 2963.625 ;
        RECT 6.295 2960.535 6.815 2961.075 ;
        RECT 5.605 2959.445 6.815 2960.535 ;
        RECT 2912.805 2960.535 2913.325 2961.075 ;
        RECT 2912.805 2959.445 2914.015 2960.535 ;
        RECT 5.520 2959.275 6.900 2959.445 ;
        RECT 2909.960 2959.275 2910.420 2959.445 ;
        RECT 2912.720 2959.275 2914.100 2959.445 ;
        RECT 5.605 2958.185 6.815 2959.275 ;
        RECT 6.295 2957.645 6.815 2958.185 ;
        RECT 2910.045 2958.110 2910.335 2959.275 ;
        RECT 2912.805 2958.185 2914.015 2959.275 ;
        RECT 2912.805 2957.645 2913.325 2958.185 ;
        RECT 6.295 2955.095 6.815 2955.635 ;
        RECT 5.605 2954.005 6.815 2955.095 ;
        RECT 2912.805 2955.095 2913.325 2955.635 ;
        RECT 9.015 2954.005 9.345 2954.730 ;
        RECT 2912.805 2954.005 2914.015 2955.095 ;
        RECT 5.520 2953.835 6.900 2954.005 ;
        RECT 8.740 2953.835 10.120 2954.005 ;
        RECT 2909.960 2953.835 2910.420 2954.005 ;
        RECT 2912.720 2953.835 2914.100 2954.005 ;
        RECT 5.605 2952.745 6.815 2953.835 ;
        RECT 6.295 2952.205 6.815 2952.745 ;
        RECT 2910.045 2952.670 2910.335 2953.835 ;
        RECT 2912.805 2952.745 2914.015 2953.835 ;
        RECT 2912.805 2952.205 2913.325 2952.745 ;
        RECT 6.295 2949.655 6.815 2950.195 ;
        RECT 5.605 2948.565 6.815 2949.655 ;
        RECT 2912.805 2949.655 2913.325 2950.195 ;
        RECT 2912.805 2948.565 2914.015 2949.655 ;
        RECT 5.520 2948.395 6.900 2948.565 ;
        RECT 2909.960 2948.395 2910.420 2948.565 ;
        RECT 2912.720 2948.395 2914.100 2948.565 ;
        RECT 5.605 2947.305 6.815 2948.395 ;
        RECT 6.295 2946.765 6.815 2947.305 ;
        RECT 2910.045 2947.230 2910.335 2948.395 ;
        RECT 2912.805 2947.305 2914.015 2948.395 ;
        RECT 2912.805 2946.765 2913.325 2947.305 ;
        RECT 6.295 2944.215 6.815 2944.755 ;
        RECT 5.605 2943.125 6.815 2944.215 ;
        RECT 2912.805 2944.215 2913.325 2944.755 ;
        RECT 2912.805 2943.125 2914.015 2944.215 ;
        RECT 5.520 2942.955 6.900 2943.125 ;
        RECT 2909.960 2942.955 2910.420 2943.125 ;
        RECT 2912.720 2942.955 2914.100 2943.125 ;
        RECT 5.605 2941.865 6.815 2942.955 ;
        RECT 6.295 2941.325 6.815 2941.865 ;
        RECT 2910.045 2941.790 2910.335 2942.955 ;
        RECT 2912.805 2941.865 2914.015 2942.955 ;
        RECT 2912.805 2941.325 2913.325 2941.865 ;
        RECT 6.295 2938.775 6.815 2939.315 ;
        RECT 5.605 2937.685 6.815 2938.775 ;
        RECT 2912.805 2938.775 2913.325 2939.315 ;
        RECT 2912.805 2937.685 2914.015 2938.775 ;
        RECT 5.520 2937.515 6.900 2937.685 ;
        RECT 2909.960 2937.515 2910.420 2937.685 ;
        RECT 2912.720 2937.515 2914.100 2937.685 ;
        RECT 5.605 2936.425 6.815 2937.515 ;
        RECT 6.295 2935.885 6.815 2936.425 ;
        RECT 2910.045 2936.350 2910.335 2937.515 ;
        RECT 2912.805 2936.425 2914.015 2937.515 ;
        RECT 2912.805 2935.885 2913.325 2936.425 ;
        RECT 6.295 2933.335 6.815 2933.875 ;
        RECT 5.605 2932.245 6.815 2933.335 ;
        RECT 2912.805 2933.335 2913.325 2933.875 ;
        RECT 2912.805 2932.245 2914.015 2933.335 ;
        RECT 5.520 2932.075 6.900 2932.245 ;
        RECT 2909.960 2932.075 2910.420 2932.245 ;
        RECT 2912.720 2932.075 2914.100 2932.245 ;
        RECT 5.605 2930.985 6.815 2932.075 ;
        RECT 6.295 2930.445 6.815 2930.985 ;
        RECT 2910.045 2930.910 2910.335 2932.075 ;
        RECT 2912.805 2930.985 2914.015 2932.075 ;
        RECT 2912.805 2930.445 2913.325 2930.985 ;
        RECT 6.295 2927.895 6.815 2928.435 ;
        RECT 5.605 2926.805 6.815 2927.895 ;
        RECT 2912.805 2927.895 2913.325 2928.435 ;
        RECT 2912.805 2926.805 2914.015 2927.895 ;
        RECT 5.520 2926.635 6.900 2926.805 ;
        RECT 2909.960 2926.635 2910.420 2926.805 ;
        RECT 2912.720 2926.635 2914.100 2926.805 ;
        RECT 5.605 2925.545 6.815 2926.635 ;
        RECT 6.295 2925.005 6.815 2925.545 ;
        RECT 2910.045 2925.470 2910.335 2926.635 ;
        RECT 2912.805 2925.545 2914.015 2926.635 ;
        RECT 2912.805 2925.005 2913.325 2925.545 ;
        RECT 6.295 2922.455 6.815 2922.995 ;
        RECT 5.605 2921.365 6.815 2922.455 ;
        RECT 2912.805 2922.455 2913.325 2922.995 ;
        RECT 2912.805 2921.365 2914.015 2922.455 ;
        RECT 5.520 2921.195 6.900 2921.365 ;
        RECT 2909.960 2921.195 2910.420 2921.365 ;
        RECT 2912.720 2921.195 2914.100 2921.365 ;
        RECT 5.605 2920.105 6.815 2921.195 ;
        RECT 6.295 2919.565 6.815 2920.105 ;
        RECT 2910.045 2920.030 2910.335 2921.195 ;
        RECT 2912.805 2920.105 2914.015 2921.195 ;
        RECT 2912.805 2919.565 2913.325 2920.105 ;
        RECT 6.295 2917.015 6.815 2917.555 ;
        RECT 5.605 2915.925 6.815 2917.015 ;
        RECT 2912.805 2917.015 2913.325 2917.555 ;
        RECT 2912.805 2915.925 2914.015 2917.015 ;
        RECT 5.520 2915.755 6.900 2915.925 ;
        RECT 2909.960 2915.755 2911.800 2915.925 ;
        RECT 2912.720 2915.755 2914.100 2915.925 ;
        RECT 5.605 2914.665 6.815 2915.755 ;
        RECT 6.295 2914.125 6.815 2914.665 ;
        RECT 2910.045 2914.590 2910.335 2915.755 ;
        RECT 2910.695 2915.030 2911.025 2915.755 ;
        RECT 2912.805 2914.665 2914.015 2915.755 ;
        RECT 2912.805 2914.125 2913.325 2914.665 ;
        RECT 6.295 2911.575 6.815 2912.115 ;
        RECT 5.605 2910.485 6.815 2911.575 ;
        RECT 2912.805 2911.575 2913.325 2912.115 ;
        RECT 2912.805 2910.485 2914.015 2911.575 ;
        RECT 5.520 2910.315 6.900 2910.485 ;
        RECT 2909.960 2910.315 2910.420 2910.485 ;
        RECT 2912.720 2910.315 2914.100 2910.485 ;
        RECT 5.605 2909.225 6.815 2910.315 ;
        RECT 6.295 2908.685 6.815 2909.225 ;
        RECT 2910.045 2909.150 2910.335 2910.315 ;
        RECT 2912.805 2909.225 2914.015 2910.315 ;
        RECT 2912.805 2908.685 2913.325 2909.225 ;
        RECT 6.295 2906.135 6.815 2906.675 ;
        RECT 5.605 2905.045 6.815 2906.135 ;
        RECT 2912.805 2906.135 2913.325 2906.675 ;
        RECT 2912.805 2905.045 2914.015 2906.135 ;
        RECT 5.520 2904.875 6.900 2905.045 ;
        RECT 2909.960 2904.875 2910.420 2905.045 ;
        RECT 2912.720 2904.875 2914.100 2905.045 ;
        RECT 5.605 2903.785 6.815 2904.875 ;
        RECT 6.295 2903.245 6.815 2903.785 ;
        RECT 2910.045 2903.710 2910.335 2904.875 ;
        RECT 2912.805 2903.785 2914.015 2904.875 ;
        RECT 2912.805 2903.245 2913.325 2903.785 ;
        RECT 6.295 2900.695 6.815 2901.235 ;
        RECT 5.605 2899.605 6.815 2900.695 ;
        RECT 2912.805 2900.695 2913.325 2901.235 ;
        RECT 2912.805 2899.605 2914.015 2900.695 ;
        RECT 5.520 2899.435 6.900 2899.605 ;
        RECT 2909.960 2899.435 2910.420 2899.605 ;
        RECT 2912.720 2899.435 2914.100 2899.605 ;
        RECT 5.605 2898.345 6.815 2899.435 ;
        RECT 6.295 2897.805 6.815 2898.345 ;
        RECT 2910.045 2898.270 2910.335 2899.435 ;
        RECT 2912.805 2898.345 2914.015 2899.435 ;
        RECT 2912.805 2897.805 2913.325 2898.345 ;
        RECT 6.295 2895.255 6.815 2895.795 ;
        RECT 5.605 2894.165 6.815 2895.255 ;
        RECT 2912.805 2895.255 2913.325 2895.795 ;
        RECT 2912.805 2894.165 2914.015 2895.255 ;
        RECT 5.520 2893.995 6.900 2894.165 ;
        RECT 2909.960 2893.995 2910.420 2894.165 ;
        RECT 2912.720 2893.995 2914.100 2894.165 ;
        RECT 5.605 2892.905 6.815 2893.995 ;
        RECT 6.295 2892.365 6.815 2892.905 ;
        RECT 2910.045 2892.830 2910.335 2893.995 ;
        RECT 2912.805 2892.905 2914.015 2893.995 ;
        RECT 2912.805 2892.365 2913.325 2892.905 ;
        RECT 6.295 2889.815 6.815 2890.355 ;
        RECT 5.605 2888.725 6.815 2889.815 ;
        RECT 2912.805 2889.815 2913.325 2890.355 ;
        RECT 2912.805 2888.725 2914.015 2889.815 ;
        RECT 5.520 2888.555 6.900 2888.725 ;
        RECT 2909.960 2888.555 2910.420 2888.725 ;
        RECT 2912.720 2888.555 2914.100 2888.725 ;
        RECT 5.605 2887.465 6.815 2888.555 ;
        RECT 6.295 2886.925 6.815 2887.465 ;
        RECT 2910.045 2887.390 2910.335 2888.555 ;
        RECT 2912.805 2887.465 2914.015 2888.555 ;
        RECT 2912.805 2886.925 2913.325 2887.465 ;
        RECT 6.295 2884.375 6.815 2884.915 ;
        RECT 5.605 2883.285 6.815 2884.375 ;
        RECT 2912.805 2884.375 2913.325 2884.915 ;
        RECT 9.015 2883.285 9.345 2884.010 ;
        RECT 2912.805 2883.285 2914.015 2884.375 ;
        RECT 5.520 2883.115 6.900 2883.285 ;
        RECT 8.740 2883.115 10.120 2883.285 ;
        RECT 2909.960 2883.115 2910.420 2883.285 ;
        RECT 2912.720 2883.115 2914.100 2883.285 ;
        RECT 5.605 2882.025 6.815 2883.115 ;
        RECT 6.295 2881.485 6.815 2882.025 ;
        RECT 2910.045 2881.950 2910.335 2883.115 ;
        RECT 2912.805 2882.025 2914.015 2883.115 ;
        RECT 2912.805 2881.485 2913.325 2882.025 ;
        RECT 6.295 2878.935 6.815 2879.475 ;
        RECT 5.605 2877.845 6.815 2878.935 ;
        RECT 2912.805 2878.935 2913.325 2879.475 ;
        RECT 2912.805 2877.845 2914.015 2878.935 ;
        RECT 5.520 2877.675 6.900 2877.845 ;
        RECT 2909.960 2877.675 2910.420 2877.845 ;
        RECT 2912.720 2877.675 2914.100 2877.845 ;
        RECT 5.605 2876.585 6.815 2877.675 ;
        RECT 6.295 2876.045 6.815 2876.585 ;
        RECT 2910.045 2876.510 2910.335 2877.675 ;
        RECT 2912.805 2876.585 2914.015 2877.675 ;
        RECT 2912.805 2876.045 2913.325 2876.585 ;
        RECT 6.295 2873.495 6.815 2874.035 ;
        RECT 5.605 2872.405 6.815 2873.495 ;
        RECT 2912.805 2873.495 2913.325 2874.035 ;
        RECT 2912.805 2872.405 2914.015 2873.495 ;
        RECT 5.520 2872.235 6.900 2872.405 ;
        RECT 8.740 2872.235 10.120 2872.405 ;
        RECT 2909.960 2872.235 2910.420 2872.405 ;
        RECT 2912.720 2872.235 2914.100 2872.405 ;
        RECT 5.605 2871.145 6.815 2872.235 ;
        RECT 9.015 2871.510 9.345 2872.235 ;
        RECT 6.295 2870.605 6.815 2871.145 ;
        RECT 2910.045 2871.070 2910.335 2872.235 ;
        RECT 2912.805 2871.145 2914.015 2872.235 ;
        RECT 2912.805 2870.605 2913.325 2871.145 ;
        RECT 6.295 2868.055 6.815 2868.595 ;
        RECT 5.605 2866.965 6.815 2868.055 ;
        RECT 2912.805 2868.055 2913.325 2868.595 ;
        RECT 2912.805 2866.965 2914.015 2868.055 ;
        RECT 5.520 2866.795 6.900 2866.965 ;
        RECT 2909.960 2866.795 2910.420 2866.965 ;
        RECT 2912.720 2866.795 2914.100 2866.965 ;
        RECT 5.605 2865.705 6.815 2866.795 ;
        RECT 6.295 2865.165 6.815 2865.705 ;
        RECT 2910.045 2865.630 2910.335 2866.795 ;
        RECT 2912.805 2865.705 2914.015 2866.795 ;
        RECT 2912.805 2865.165 2913.325 2865.705 ;
        RECT 6.295 2862.615 6.815 2863.155 ;
        RECT 5.605 2861.525 6.815 2862.615 ;
        RECT 2912.805 2862.615 2913.325 2863.155 ;
        RECT 2912.805 2861.525 2914.015 2862.615 ;
        RECT 5.520 2861.355 6.900 2861.525 ;
        RECT 2909.960 2861.355 2910.420 2861.525 ;
        RECT 2912.720 2861.355 2914.100 2861.525 ;
        RECT 5.605 2860.265 6.815 2861.355 ;
        RECT 6.295 2859.725 6.815 2860.265 ;
        RECT 2910.045 2860.190 2910.335 2861.355 ;
        RECT 2912.805 2860.265 2914.015 2861.355 ;
        RECT 2912.805 2859.725 2913.325 2860.265 ;
        RECT 6.295 2857.175 6.815 2857.715 ;
        RECT 5.605 2856.085 6.815 2857.175 ;
        RECT 2912.805 2857.175 2913.325 2857.715 ;
        RECT 2912.805 2856.085 2914.015 2857.175 ;
        RECT 5.520 2855.915 6.900 2856.085 ;
        RECT 2909.960 2855.915 2910.420 2856.085 ;
        RECT 2912.720 2855.915 2914.100 2856.085 ;
        RECT 5.605 2854.825 6.815 2855.915 ;
        RECT 6.295 2854.285 6.815 2854.825 ;
        RECT 2910.045 2854.750 2910.335 2855.915 ;
        RECT 2912.805 2854.825 2914.015 2855.915 ;
        RECT 2912.805 2854.285 2913.325 2854.825 ;
        RECT 6.295 2851.735 6.815 2852.275 ;
        RECT 5.605 2850.645 6.815 2851.735 ;
        RECT 2912.805 2851.735 2913.325 2852.275 ;
        RECT 2912.805 2850.645 2914.015 2851.735 ;
        RECT 5.520 2850.475 6.900 2850.645 ;
        RECT 2909.960 2850.475 2910.420 2850.645 ;
        RECT 2912.720 2850.475 2914.100 2850.645 ;
        RECT 5.605 2849.385 6.815 2850.475 ;
        RECT 6.295 2848.845 6.815 2849.385 ;
        RECT 2910.045 2849.310 2910.335 2850.475 ;
        RECT 2912.805 2849.385 2914.015 2850.475 ;
        RECT 2912.805 2848.845 2913.325 2849.385 ;
        RECT 6.295 2846.295 6.815 2846.835 ;
        RECT 5.605 2845.205 6.815 2846.295 ;
        RECT 2912.805 2846.295 2913.325 2846.835 ;
        RECT 2912.805 2845.205 2914.015 2846.295 ;
        RECT 5.520 2845.035 6.900 2845.205 ;
        RECT 2909.960 2845.035 2910.420 2845.205 ;
        RECT 2912.720 2845.035 2914.100 2845.205 ;
        RECT 5.605 2843.945 6.815 2845.035 ;
        RECT 6.295 2843.405 6.815 2843.945 ;
        RECT 2910.045 2843.870 2910.335 2845.035 ;
        RECT 2912.805 2843.945 2914.015 2845.035 ;
        RECT 2912.805 2843.405 2913.325 2843.945 ;
        RECT 6.295 2840.855 6.815 2841.395 ;
        RECT 5.605 2839.765 6.815 2840.855 ;
        RECT 2912.805 2840.855 2913.325 2841.395 ;
        RECT 2912.805 2839.765 2914.015 2840.855 ;
        RECT 5.520 2839.595 6.900 2839.765 ;
        RECT 2909.960 2839.595 2910.420 2839.765 ;
        RECT 2912.720 2839.595 2914.100 2839.765 ;
        RECT 5.605 2838.505 6.815 2839.595 ;
        RECT 6.295 2837.965 6.815 2838.505 ;
        RECT 2910.045 2838.430 2910.335 2839.595 ;
        RECT 2912.805 2838.505 2914.015 2839.595 ;
        RECT 2912.805 2837.965 2913.325 2838.505 ;
        RECT 6.295 2835.415 6.815 2835.955 ;
        RECT 5.605 2834.325 6.815 2835.415 ;
        RECT 2912.805 2835.415 2913.325 2835.955 ;
        RECT 2912.805 2834.325 2914.015 2835.415 ;
        RECT 5.520 2834.155 6.900 2834.325 ;
        RECT 2909.960 2834.155 2910.420 2834.325 ;
        RECT 2912.720 2834.155 2914.100 2834.325 ;
        RECT 5.605 2833.065 6.815 2834.155 ;
        RECT 6.295 2832.525 6.815 2833.065 ;
        RECT 2910.045 2832.990 2910.335 2834.155 ;
        RECT 2912.805 2833.065 2914.015 2834.155 ;
        RECT 2912.805 2832.525 2913.325 2833.065 ;
        RECT 6.295 2829.975 6.815 2830.515 ;
        RECT 5.605 2828.885 6.815 2829.975 ;
        RECT 2912.805 2829.975 2913.325 2830.515 ;
        RECT 2912.805 2828.885 2914.015 2829.975 ;
        RECT 5.520 2828.715 6.900 2828.885 ;
        RECT 2909.960 2828.715 2910.420 2828.885 ;
        RECT 2912.720 2828.715 2914.100 2828.885 ;
        RECT 5.605 2827.625 6.815 2828.715 ;
        RECT 6.295 2827.085 6.815 2827.625 ;
        RECT 2910.045 2827.550 2910.335 2828.715 ;
        RECT 2912.805 2827.625 2914.015 2828.715 ;
        RECT 2912.805 2827.085 2913.325 2827.625 ;
        RECT 6.295 2824.535 6.815 2825.075 ;
        RECT 5.605 2823.445 6.815 2824.535 ;
        RECT 2912.805 2824.535 2913.325 2825.075 ;
        RECT 2912.805 2823.445 2914.015 2824.535 ;
        RECT 5.520 2823.275 6.900 2823.445 ;
        RECT 2909.960 2823.275 2910.420 2823.445 ;
        RECT 2912.720 2823.275 2914.100 2823.445 ;
        RECT 5.605 2822.185 6.815 2823.275 ;
        RECT 6.295 2821.645 6.815 2822.185 ;
        RECT 2910.045 2822.110 2910.335 2823.275 ;
        RECT 2912.805 2822.185 2914.015 2823.275 ;
        RECT 2912.805 2821.645 2913.325 2822.185 ;
        RECT 6.295 2819.095 6.815 2819.635 ;
        RECT 5.605 2818.005 6.815 2819.095 ;
        RECT 2912.805 2819.095 2913.325 2819.635 ;
        RECT 2912.805 2818.005 2914.015 2819.095 ;
        RECT 5.520 2817.835 6.900 2818.005 ;
        RECT 2909.960 2817.835 2910.420 2818.005 ;
        RECT 2912.720 2817.835 2914.100 2818.005 ;
        RECT 5.605 2816.745 6.815 2817.835 ;
        RECT 6.295 2816.205 6.815 2816.745 ;
        RECT 2910.045 2816.670 2910.335 2817.835 ;
        RECT 2912.805 2816.745 2914.015 2817.835 ;
        RECT 2912.805 2816.205 2913.325 2816.745 ;
        RECT 6.295 2813.655 6.815 2814.195 ;
        RECT 5.605 2812.565 6.815 2813.655 ;
        RECT 2912.805 2813.655 2913.325 2814.195 ;
        RECT 2912.805 2812.565 2914.015 2813.655 ;
        RECT 5.520 2812.395 6.900 2812.565 ;
        RECT 2909.960 2812.395 2910.420 2812.565 ;
        RECT 2912.720 2812.395 2914.100 2812.565 ;
        RECT 5.605 2811.305 6.815 2812.395 ;
        RECT 6.295 2810.765 6.815 2811.305 ;
        RECT 2910.045 2811.230 2910.335 2812.395 ;
        RECT 2912.805 2811.305 2914.015 2812.395 ;
        RECT 2912.805 2810.765 2913.325 2811.305 ;
        RECT 6.295 2808.215 6.815 2808.755 ;
        RECT 5.605 2807.125 6.815 2808.215 ;
        RECT 2912.805 2808.215 2913.325 2808.755 ;
        RECT 2912.805 2807.125 2914.015 2808.215 ;
        RECT 5.520 2806.955 6.900 2807.125 ;
        RECT 2909.960 2806.955 2910.420 2807.125 ;
        RECT 2912.720 2806.955 2914.100 2807.125 ;
        RECT 5.605 2805.865 6.815 2806.955 ;
        RECT 6.295 2805.325 6.815 2805.865 ;
        RECT 2910.045 2805.790 2910.335 2806.955 ;
        RECT 2912.805 2805.865 2914.015 2806.955 ;
        RECT 2912.805 2805.325 2913.325 2805.865 ;
        RECT 6.295 2802.775 6.815 2803.315 ;
        RECT 5.605 2801.685 6.815 2802.775 ;
        RECT 2912.805 2802.775 2913.325 2803.315 ;
        RECT 2912.805 2801.685 2914.015 2802.775 ;
        RECT 5.520 2801.515 6.900 2801.685 ;
        RECT 2909.960 2801.515 2910.420 2801.685 ;
        RECT 2912.720 2801.515 2914.100 2801.685 ;
        RECT 5.605 2800.425 6.815 2801.515 ;
        RECT 6.295 2799.885 6.815 2800.425 ;
        RECT 2910.045 2800.350 2910.335 2801.515 ;
        RECT 2912.805 2800.425 2914.015 2801.515 ;
        RECT 2912.805 2799.885 2913.325 2800.425 ;
        RECT 6.295 2797.335 6.815 2797.875 ;
        RECT 5.605 2796.245 6.815 2797.335 ;
        RECT 2912.805 2797.335 2913.325 2797.875 ;
        RECT 2912.805 2796.245 2914.015 2797.335 ;
        RECT 5.520 2796.075 6.900 2796.245 ;
        RECT 2909.960 2796.075 2910.420 2796.245 ;
        RECT 2912.720 2796.075 2914.100 2796.245 ;
        RECT 5.605 2794.985 6.815 2796.075 ;
        RECT 6.295 2794.445 6.815 2794.985 ;
        RECT 2910.045 2794.910 2910.335 2796.075 ;
        RECT 2912.805 2794.985 2914.015 2796.075 ;
        RECT 2912.805 2794.445 2913.325 2794.985 ;
        RECT 6.295 2791.895 6.815 2792.435 ;
        RECT 5.605 2790.805 6.815 2791.895 ;
        RECT 2912.805 2791.895 2913.325 2792.435 ;
        RECT 2912.805 2790.805 2914.015 2791.895 ;
        RECT 5.520 2790.635 6.900 2790.805 ;
        RECT 2909.960 2790.635 2910.420 2790.805 ;
        RECT 2912.720 2790.635 2914.100 2790.805 ;
        RECT 5.605 2789.545 6.815 2790.635 ;
        RECT 6.295 2789.005 6.815 2789.545 ;
        RECT 2910.045 2789.470 2910.335 2790.635 ;
        RECT 2912.805 2789.545 2914.015 2790.635 ;
        RECT 2912.805 2789.005 2913.325 2789.545 ;
        RECT 6.295 2786.455 6.815 2786.995 ;
        RECT 5.605 2785.365 6.815 2786.455 ;
        RECT 2912.805 2786.455 2913.325 2786.995 ;
        RECT 2912.805 2785.365 2914.015 2786.455 ;
        RECT 5.520 2785.195 6.900 2785.365 ;
        RECT 2909.960 2785.195 2910.420 2785.365 ;
        RECT 2912.720 2785.195 2914.100 2785.365 ;
        RECT 5.605 2784.105 6.815 2785.195 ;
        RECT 6.295 2783.565 6.815 2784.105 ;
        RECT 2910.045 2784.030 2910.335 2785.195 ;
        RECT 2912.805 2784.105 2914.015 2785.195 ;
        RECT 2912.805 2783.565 2913.325 2784.105 ;
        RECT 6.295 2781.015 6.815 2781.555 ;
        RECT 5.605 2779.925 6.815 2781.015 ;
        RECT 2912.805 2781.015 2913.325 2781.555 ;
        RECT 2912.805 2779.925 2914.015 2781.015 ;
        RECT 5.520 2779.755 6.900 2779.925 ;
        RECT 2909.960 2779.755 2910.420 2779.925 ;
        RECT 2912.720 2779.755 2914.100 2779.925 ;
        RECT 5.605 2778.665 6.815 2779.755 ;
        RECT 6.295 2778.125 6.815 2778.665 ;
        RECT 2910.045 2778.590 2910.335 2779.755 ;
        RECT 2912.805 2778.665 2914.015 2779.755 ;
        RECT 2912.805 2778.125 2913.325 2778.665 ;
        RECT 6.295 2775.575 6.815 2776.115 ;
        RECT 5.605 2774.485 6.815 2775.575 ;
        RECT 2912.805 2775.575 2913.325 2776.115 ;
        RECT 2909.315 2774.485 2909.645 2775.210 ;
        RECT 2912.805 2774.485 2914.015 2775.575 ;
        RECT 5.520 2774.315 6.900 2774.485 ;
        RECT 2909.040 2774.315 2910.420 2774.485 ;
        RECT 2912.720 2774.315 2914.100 2774.485 ;
        RECT 5.605 2773.225 6.815 2774.315 ;
        RECT 6.295 2772.685 6.815 2773.225 ;
        RECT 2910.045 2773.150 2910.335 2774.315 ;
        RECT 2912.805 2773.225 2914.015 2774.315 ;
        RECT 2912.805 2772.685 2913.325 2773.225 ;
        RECT 6.295 2770.135 6.815 2770.675 ;
        RECT 5.605 2769.045 6.815 2770.135 ;
        RECT 2912.805 2770.135 2913.325 2770.675 ;
        RECT 2912.805 2769.045 2914.015 2770.135 ;
        RECT 5.520 2768.875 6.900 2769.045 ;
        RECT 2909.960 2768.875 2910.420 2769.045 ;
        RECT 2912.720 2768.875 2914.100 2769.045 ;
        RECT 5.605 2767.785 6.815 2768.875 ;
        RECT 6.295 2767.245 6.815 2767.785 ;
        RECT 2910.045 2767.710 2910.335 2768.875 ;
        RECT 2912.805 2767.785 2914.015 2768.875 ;
        RECT 2912.805 2767.245 2913.325 2767.785 ;
        RECT 6.295 2764.695 6.815 2765.235 ;
        RECT 5.605 2763.605 6.815 2764.695 ;
        RECT 2912.805 2764.695 2913.325 2765.235 ;
        RECT 2912.805 2763.605 2914.015 2764.695 ;
        RECT 5.520 2763.435 6.900 2763.605 ;
        RECT 2909.960 2763.435 2910.420 2763.605 ;
        RECT 2912.720 2763.435 2914.100 2763.605 ;
        RECT 5.605 2762.345 6.815 2763.435 ;
        RECT 6.295 2761.805 6.815 2762.345 ;
        RECT 2910.045 2762.270 2910.335 2763.435 ;
        RECT 2912.805 2762.345 2914.015 2763.435 ;
        RECT 2912.805 2761.805 2913.325 2762.345 ;
        RECT 6.295 2759.255 6.815 2759.795 ;
        RECT 5.605 2758.165 6.815 2759.255 ;
        RECT 2912.805 2759.255 2913.325 2759.795 ;
        RECT 2912.805 2758.165 2914.015 2759.255 ;
        RECT 5.520 2757.995 6.900 2758.165 ;
        RECT 2909.960 2757.995 2910.420 2758.165 ;
        RECT 2912.720 2757.995 2914.100 2758.165 ;
        RECT 5.605 2756.905 6.815 2757.995 ;
        RECT 6.295 2756.365 6.815 2756.905 ;
        RECT 2910.045 2756.830 2910.335 2757.995 ;
        RECT 2912.805 2756.905 2914.015 2757.995 ;
        RECT 2912.805 2756.365 2913.325 2756.905 ;
        RECT 6.295 2753.815 6.815 2754.355 ;
        RECT 5.605 2752.725 6.815 2753.815 ;
        RECT 2912.805 2753.815 2913.325 2754.355 ;
        RECT 2912.805 2752.725 2914.015 2753.815 ;
        RECT 5.520 2752.555 6.900 2752.725 ;
        RECT 2909.960 2752.555 2910.420 2752.725 ;
        RECT 2912.720 2752.555 2914.100 2752.725 ;
        RECT 5.605 2751.465 6.815 2752.555 ;
        RECT 6.295 2750.925 6.815 2751.465 ;
        RECT 2910.045 2751.390 2910.335 2752.555 ;
        RECT 2912.805 2751.465 2914.015 2752.555 ;
        RECT 2912.805 2750.925 2913.325 2751.465 ;
        RECT 6.295 2748.375 6.815 2748.915 ;
        RECT 5.605 2747.285 6.815 2748.375 ;
        RECT 2912.805 2748.375 2913.325 2748.915 ;
        RECT 2912.805 2747.285 2914.015 2748.375 ;
        RECT 5.520 2747.115 6.900 2747.285 ;
        RECT 2909.960 2747.115 2910.420 2747.285 ;
        RECT 2912.720 2747.115 2914.100 2747.285 ;
        RECT 5.605 2746.025 6.815 2747.115 ;
        RECT 6.295 2745.485 6.815 2746.025 ;
        RECT 2910.045 2745.950 2910.335 2747.115 ;
        RECT 2912.805 2746.025 2914.015 2747.115 ;
        RECT 2912.805 2745.485 2913.325 2746.025 ;
        RECT 6.295 2742.935 6.815 2743.475 ;
        RECT 5.605 2741.845 6.815 2742.935 ;
        RECT 2912.805 2742.935 2913.325 2743.475 ;
        RECT 2912.805 2741.845 2914.015 2742.935 ;
        RECT 5.520 2741.675 6.900 2741.845 ;
        RECT 2909.960 2741.675 2910.420 2741.845 ;
        RECT 2912.720 2741.675 2914.100 2741.845 ;
        RECT 5.605 2740.585 6.815 2741.675 ;
        RECT 6.295 2740.045 6.815 2740.585 ;
        RECT 2910.045 2740.510 2910.335 2741.675 ;
        RECT 2912.805 2740.585 2914.015 2741.675 ;
        RECT 2912.805 2740.045 2913.325 2740.585 ;
        RECT 6.295 2737.495 6.815 2738.035 ;
        RECT 5.605 2736.405 6.815 2737.495 ;
        RECT 2912.805 2737.495 2913.325 2738.035 ;
        RECT 2912.805 2736.405 2914.015 2737.495 ;
        RECT 5.520 2736.235 6.900 2736.405 ;
        RECT 2909.960 2736.235 2910.420 2736.405 ;
        RECT 2912.720 2736.235 2914.100 2736.405 ;
        RECT 5.605 2735.145 6.815 2736.235 ;
        RECT 6.295 2734.605 6.815 2735.145 ;
        RECT 2910.045 2735.070 2910.335 2736.235 ;
        RECT 2912.805 2735.145 2914.015 2736.235 ;
        RECT 2912.805 2734.605 2913.325 2735.145 ;
        RECT 6.295 2732.055 6.815 2732.595 ;
        RECT 5.605 2730.965 6.815 2732.055 ;
        RECT 2912.805 2732.055 2913.325 2732.595 ;
        RECT 2912.805 2730.965 2914.015 2732.055 ;
        RECT 5.520 2730.795 6.900 2730.965 ;
        RECT 2909.960 2730.795 2910.420 2730.965 ;
        RECT 2912.720 2730.795 2914.100 2730.965 ;
        RECT 5.605 2729.705 6.815 2730.795 ;
        RECT 6.295 2729.165 6.815 2729.705 ;
        RECT 2910.045 2729.630 2910.335 2730.795 ;
        RECT 2912.805 2729.705 2914.015 2730.795 ;
        RECT 2912.805 2729.165 2913.325 2729.705 ;
        RECT 6.295 2726.615 6.815 2727.155 ;
        RECT 5.605 2725.525 6.815 2726.615 ;
        RECT 2912.805 2726.615 2913.325 2727.155 ;
        RECT 2912.805 2725.525 2914.015 2726.615 ;
        RECT 5.520 2725.355 6.900 2725.525 ;
        RECT 2909.960 2725.355 2910.420 2725.525 ;
        RECT 2912.720 2725.355 2914.100 2725.525 ;
        RECT 5.605 2724.265 6.815 2725.355 ;
        RECT 6.295 2723.725 6.815 2724.265 ;
        RECT 2910.045 2724.190 2910.335 2725.355 ;
        RECT 2912.805 2724.265 2914.015 2725.355 ;
        RECT 2912.805 2723.725 2913.325 2724.265 ;
        RECT 6.295 2721.175 6.815 2721.715 ;
        RECT 5.605 2720.085 6.815 2721.175 ;
        RECT 2912.805 2721.175 2913.325 2721.715 ;
        RECT 2912.805 2720.085 2914.015 2721.175 ;
        RECT 5.520 2719.915 6.900 2720.085 ;
        RECT 2909.960 2719.915 2910.420 2720.085 ;
        RECT 2912.720 2719.915 2914.100 2720.085 ;
        RECT 5.605 2718.825 6.815 2719.915 ;
        RECT 6.295 2718.285 6.815 2718.825 ;
        RECT 2910.045 2718.750 2910.335 2719.915 ;
        RECT 2912.805 2718.825 2914.015 2719.915 ;
        RECT 2912.805 2718.285 2913.325 2718.825 ;
        RECT 6.295 2715.735 6.815 2716.275 ;
        RECT 5.605 2714.645 6.815 2715.735 ;
        RECT 2912.805 2715.735 2913.325 2716.275 ;
        RECT 2912.805 2714.645 2914.015 2715.735 ;
        RECT 5.520 2714.475 6.900 2714.645 ;
        RECT 2909.960 2714.475 2910.420 2714.645 ;
        RECT 2912.720 2714.475 2914.100 2714.645 ;
        RECT 5.605 2713.385 6.815 2714.475 ;
        RECT 6.295 2712.845 6.815 2713.385 ;
        RECT 2910.045 2713.310 2910.335 2714.475 ;
        RECT 2912.805 2713.385 2914.015 2714.475 ;
        RECT 2912.805 2712.845 2913.325 2713.385 ;
        RECT 6.295 2710.295 6.815 2710.835 ;
        RECT 5.605 2709.205 6.815 2710.295 ;
        RECT 2912.805 2710.295 2913.325 2710.835 ;
        RECT 2912.805 2709.205 2914.015 2710.295 ;
        RECT 5.520 2709.035 6.900 2709.205 ;
        RECT 2909.960 2709.035 2910.420 2709.205 ;
        RECT 2912.720 2709.035 2914.100 2709.205 ;
        RECT 5.605 2707.945 6.815 2709.035 ;
        RECT 6.295 2707.405 6.815 2707.945 ;
        RECT 2910.045 2707.870 2910.335 2709.035 ;
        RECT 2912.805 2707.945 2914.015 2709.035 ;
        RECT 2912.805 2707.405 2913.325 2707.945 ;
        RECT 6.295 2704.855 6.815 2705.395 ;
        RECT 5.605 2703.765 6.815 2704.855 ;
        RECT 2912.805 2704.855 2913.325 2705.395 ;
        RECT 2912.805 2703.765 2914.015 2704.855 ;
        RECT 5.520 2703.595 6.900 2703.765 ;
        RECT 2909.960 2703.595 2910.420 2703.765 ;
        RECT 2912.720 2703.595 2914.100 2703.765 ;
        RECT 5.605 2702.505 6.815 2703.595 ;
        RECT 6.295 2701.965 6.815 2702.505 ;
        RECT 2910.045 2702.430 2910.335 2703.595 ;
        RECT 2912.805 2702.505 2914.015 2703.595 ;
        RECT 2912.805 2701.965 2913.325 2702.505 ;
        RECT 6.295 2699.415 6.815 2699.955 ;
        RECT 5.605 2698.325 6.815 2699.415 ;
        RECT 2912.805 2699.415 2913.325 2699.955 ;
        RECT 2912.805 2698.325 2914.015 2699.415 ;
        RECT 5.520 2698.155 6.900 2698.325 ;
        RECT 2909.960 2698.155 2910.420 2698.325 ;
        RECT 2912.720 2698.155 2914.100 2698.325 ;
        RECT 5.605 2697.065 6.815 2698.155 ;
        RECT 6.295 2696.525 6.815 2697.065 ;
        RECT 2910.045 2696.990 2910.335 2698.155 ;
        RECT 2912.805 2697.065 2914.015 2698.155 ;
        RECT 2912.805 2696.525 2913.325 2697.065 ;
        RECT 6.295 2693.975 6.815 2694.515 ;
        RECT 5.605 2692.885 6.815 2693.975 ;
        RECT 2912.805 2693.975 2913.325 2694.515 ;
        RECT 2912.805 2692.885 2914.015 2693.975 ;
        RECT 5.520 2692.715 6.900 2692.885 ;
        RECT 2912.720 2692.715 2914.100 2692.885 ;
        RECT 5.605 2691.625 6.815 2692.715 ;
        RECT 6.295 2691.085 6.815 2691.625 ;
        RECT 2912.805 2691.625 2914.015 2692.715 ;
        RECT 2912.805 2691.085 2913.325 2691.625 ;
        RECT 6.295 2688.535 6.815 2689.075 ;
        RECT 5.605 2687.445 6.815 2688.535 ;
        RECT 2906.365 2687.445 2906.655 2688.610 ;
        RECT 2912.805 2688.535 2913.325 2689.075 ;
        RECT 2912.805 2687.445 2914.015 2688.535 ;
        RECT 5.520 2687.275 6.900 2687.445 ;
        RECT 2906.300 2687.275 2906.740 2687.445 ;
        RECT 2912.720 2687.275 2914.100 2687.445 ;
        RECT 5.605 2686.185 6.815 2687.275 ;
        RECT 6.295 2685.645 6.815 2686.185 ;
        RECT 2912.805 2686.185 2914.015 2687.275 ;
        RECT 2912.805 2685.645 2913.325 2686.185 ;
        RECT 6.295 2683.095 6.815 2683.635 ;
        RECT 5.605 2682.005 6.815 2683.095 ;
        RECT 2906.365 2682.005 2906.655 2683.170 ;
        RECT 2912.805 2683.095 2913.325 2683.635 ;
        RECT 2912.805 2682.005 2914.015 2683.095 ;
        RECT 5.520 2681.835 6.900 2682.005 ;
        RECT 2906.300 2681.835 2906.740 2682.005 ;
        RECT 2912.720 2681.835 2914.100 2682.005 ;
        RECT 5.605 2680.745 6.815 2681.835 ;
        RECT 6.295 2680.205 6.815 2680.745 ;
        RECT 2912.805 2680.745 2914.015 2681.835 ;
        RECT 2912.805 2680.205 2913.325 2680.745 ;
        RECT 6.295 2677.655 6.815 2678.195 ;
        RECT 5.605 2676.565 6.815 2677.655 ;
        RECT 2906.365 2676.565 2906.655 2677.730 ;
        RECT 2912.805 2677.655 2913.325 2678.195 ;
        RECT 2912.805 2676.565 2914.015 2677.655 ;
        RECT 5.520 2676.395 6.900 2676.565 ;
        RECT 2906.300 2676.395 2906.740 2676.565 ;
        RECT 2912.720 2676.395 2914.100 2676.565 ;
        RECT 5.605 2675.305 6.815 2676.395 ;
        RECT 6.295 2674.765 6.815 2675.305 ;
        RECT 2912.805 2675.305 2914.015 2676.395 ;
        RECT 2912.805 2674.765 2913.325 2675.305 ;
        RECT 6.295 2672.215 6.815 2672.755 ;
        RECT 5.605 2671.125 6.815 2672.215 ;
        RECT 2906.365 2671.125 2906.655 2672.290 ;
        RECT 2912.805 2672.215 2913.325 2672.755 ;
        RECT 2912.805 2671.125 2914.015 2672.215 ;
        RECT 5.520 2670.955 6.900 2671.125 ;
        RECT 2906.300 2670.955 2906.740 2671.125 ;
        RECT 2912.720 2670.955 2914.100 2671.125 ;
        RECT 5.605 2669.865 6.815 2670.955 ;
        RECT 6.295 2669.325 6.815 2669.865 ;
        RECT 2912.805 2669.865 2914.015 2670.955 ;
        RECT 2912.805 2669.325 2913.325 2669.865 ;
        RECT 6.295 2666.775 6.815 2667.315 ;
        RECT 5.605 2665.685 6.815 2666.775 ;
        RECT 2906.365 2665.685 2906.655 2666.850 ;
        RECT 2912.805 2666.775 2913.325 2667.315 ;
        RECT 2912.805 2665.685 2914.015 2666.775 ;
        RECT 5.520 2665.515 6.900 2665.685 ;
        RECT 2906.300 2665.515 2906.740 2665.685 ;
        RECT 2912.720 2665.515 2914.100 2665.685 ;
        RECT 5.605 2664.425 6.815 2665.515 ;
        RECT 6.295 2663.885 6.815 2664.425 ;
        RECT 2912.805 2664.425 2914.015 2665.515 ;
        RECT 2912.805 2663.885 2913.325 2664.425 ;
        RECT 6.295 2661.335 6.815 2661.875 ;
        RECT 5.605 2660.245 6.815 2661.335 ;
        RECT 2906.365 2660.245 2906.655 2661.410 ;
        RECT 2912.805 2661.335 2913.325 2661.875 ;
        RECT 2912.805 2660.245 2914.015 2661.335 ;
        RECT 5.520 2660.075 6.900 2660.245 ;
        RECT 2906.300 2660.075 2906.740 2660.245 ;
        RECT 2912.720 2660.075 2914.100 2660.245 ;
        RECT 5.605 2658.985 6.815 2660.075 ;
        RECT 6.295 2658.445 6.815 2658.985 ;
        RECT 2912.805 2658.985 2914.015 2660.075 ;
        RECT 2912.805 2658.445 2913.325 2658.985 ;
        RECT 6.295 2655.895 6.815 2656.435 ;
        RECT 5.605 2654.805 6.815 2655.895 ;
        RECT 2906.365 2654.805 2906.655 2655.970 ;
        RECT 2912.805 2655.895 2913.325 2656.435 ;
        RECT 2912.805 2654.805 2914.015 2655.895 ;
        RECT 5.520 2654.635 6.900 2654.805 ;
        RECT 2906.300 2654.635 2906.740 2654.805 ;
        RECT 2912.720 2654.635 2914.100 2654.805 ;
        RECT 5.605 2653.545 6.815 2654.635 ;
        RECT 6.295 2653.005 6.815 2653.545 ;
        RECT 2912.805 2653.545 2914.015 2654.635 ;
        RECT 2912.805 2653.005 2913.325 2653.545 ;
        RECT 6.295 2650.455 6.815 2650.995 ;
        RECT 5.605 2649.365 6.815 2650.455 ;
        RECT 2906.365 2649.365 2906.655 2650.530 ;
        RECT 2912.805 2650.455 2913.325 2650.995 ;
        RECT 2912.805 2649.365 2914.015 2650.455 ;
        RECT 5.520 2649.195 6.900 2649.365 ;
        RECT 2906.300 2649.195 2906.740 2649.365 ;
        RECT 2912.720 2649.195 2914.100 2649.365 ;
        RECT 5.605 2648.105 6.815 2649.195 ;
        RECT 6.295 2647.565 6.815 2648.105 ;
        RECT 2912.805 2648.105 2914.015 2649.195 ;
        RECT 2912.805 2647.565 2913.325 2648.105 ;
        RECT 6.295 2645.015 6.815 2645.555 ;
        RECT 5.605 2643.925 6.815 2645.015 ;
        RECT 2906.365 2643.925 2906.655 2645.090 ;
        RECT 2912.805 2645.015 2913.325 2645.555 ;
        RECT 2912.805 2643.925 2914.015 2645.015 ;
        RECT 5.520 2643.755 6.900 2643.925 ;
        RECT 2906.300 2643.755 2906.740 2643.925 ;
        RECT 2912.720 2643.755 2914.100 2643.925 ;
        RECT 5.605 2642.665 6.815 2643.755 ;
        RECT 6.295 2642.125 6.815 2642.665 ;
        RECT 2912.805 2642.665 2914.015 2643.755 ;
        RECT 2912.805 2642.125 2913.325 2642.665 ;
        RECT 6.295 2639.575 6.815 2640.115 ;
        RECT 5.605 2638.485 6.815 2639.575 ;
        RECT 2906.365 2638.485 2906.655 2639.650 ;
        RECT 2912.805 2639.575 2913.325 2640.115 ;
        RECT 2912.805 2638.485 2914.015 2639.575 ;
        RECT 5.520 2638.315 6.900 2638.485 ;
        RECT 2906.300 2638.315 2906.740 2638.485 ;
        RECT 2912.720 2638.315 2914.100 2638.485 ;
        RECT 5.605 2637.225 6.815 2638.315 ;
        RECT 6.295 2636.685 6.815 2637.225 ;
        RECT 2912.805 2637.225 2914.015 2638.315 ;
        RECT 2912.805 2636.685 2913.325 2637.225 ;
        RECT 6.295 2634.135 6.815 2634.675 ;
        RECT 5.605 2633.045 6.815 2634.135 ;
        RECT 2906.365 2633.045 2906.655 2634.210 ;
        RECT 2912.805 2634.135 2913.325 2634.675 ;
        RECT 2912.805 2633.045 2914.015 2634.135 ;
        RECT 5.520 2632.875 6.900 2633.045 ;
        RECT 2906.300 2632.875 2906.740 2633.045 ;
        RECT 2912.720 2632.875 2914.100 2633.045 ;
        RECT 5.605 2631.785 6.815 2632.875 ;
        RECT 6.295 2631.245 6.815 2631.785 ;
        RECT 2912.805 2631.785 2914.015 2632.875 ;
        RECT 2912.805 2631.245 2913.325 2631.785 ;
        RECT 6.295 2628.695 6.815 2629.235 ;
        RECT 5.605 2627.605 6.815 2628.695 ;
        RECT 2906.365 2627.605 2906.655 2628.770 ;
        RECT 2912.805 2628.695 2913.325 2629.235 ;
        RECT 2909.315 2627.605 2909.645 2628.330 ;
        RECT 2912.805 2627.605 2914.015 2628.695 ;
        RECT 5.520 2627.435 6.900 2627.605 ;
        RECT 2906.300 2627.435 2906.740 2627.605 ;
        RECT 2909.040 2627.435 2910.420 2627.605 ;
        RECT 2912.720 2627.435 2914.100 2627.605 ;
        RECT 5.605 2626.345 6.815 2627.435 ;
        RECT 6.295 2625.805 6.815 2626.345 ;
        RECT 2912.805 2626.345 2914.015 2627.435 ;
        RECT 2912.805 2625.805 2913.325 2626.345 ;
        RECT 6.295 2623.255 6.815 2623.795 ;
        RECT 5.605 2622.165 6.815 2623.255 ;
        RECT 2906.365 2622.165 2906.655 2623.330 ;
        RECT 2912.805 2623.255 2913.325 2623.795 ;
        RECT 2912.805 2622.165 2914.015 2623.255 ;
        RECT 5.520 2621.995 6.900 2622.165 ;
        RECT 2906.300 2621.995 2906.740 2622.165 ;
        RECT 2912.720 2621.995 2914.100 2622.165 ;
        RECT 5.605 2620.905 6.815 2621.995 ;
        RECT 6.295 2620.365 6.815 2620.905 ;
        RECT 2912.805 2620.905 2914.015 2621.995 ;
        RECT 2912.805 2620.365 2913.325 2620.905 ;
        RECT 6.295 2617.815 6.815 2618.355 ;
        RECT 5.605 2616.725 6.815 2617.815 ;
        RECT 2906.365 2616.725 2906.655 2617.890 ;
        RECT 2912.805 2617.815 2913.325 2618.355 ;
        RECT 2912.805 2616.725 2914.015 2617.815 ;
        RECT 5.520 2616.555 6.900 2616.725 ;
        RECT 2906.300 2616.555 2906.740 2616.725 ;
        RECT 2912.720 2616.555 2914.100 2616.725 ;
        RECT 5.605 2615.465 6.815 2616.555 ;
        RECT 6.295 2614.925 6.815 2615.465 ;
        RECT 2912.805 2615.465 2914.015 2616.555 ;
        RECT 2912.805 2614.925 2913.325 2615.465 ;
        RECT 6.295 2612.375 6.815 2612.915 ;
        RECT 5.605 2611.285 6.815 2612.375 ;
        RECT 2906.365 2611.285 2906.655 2612.450 ;
        RECT 2912.805 2612.375 2913.325 2612.915 ;
        RECT 2912.805 2611.285 2914.015 2612.375 ;
        RECT 5.520 2611.115 6.900 2611.285 ;
        RECT 2906.300 2611.115 2906.740 2611.285 ;
        RECT 2912.720 2611.115 2914.100 2611.285 ;
        RECT 5.605 2610.025 6.815 2611.115 ;
        RECT 6.295 2609.485 6.815 2610.025 ;
        RECT 2912.805 2610.025 2914.015 2611.115 ;
        RECT 2912.805 2609.485 2913.325 2610.025 ;
        RECT 6.295 2606.935 6.815 2607.475 ;
        RECT 5.605 2605.845 6.815 2606.935 ;
        RECT 2906.365 2605.845 2906.655 2607.010 ;
        RECT 2912.805 2606.935 2913.325 2607.475 ;
        RECT 2912.805 2605.845 2914.015 2606.935 ;
        RECT 5.520 2605.675 6.900 2605.845 ;
        RECT 2906.300 2605.675 2906.740 2605.845 ;
        RECT 2912.720 2605.675 2914.100 2605.845 ;
        RECT 5.605 2604.585 6.815 2605.675 ;
        RECT 6.295 2604.045 6.815 2604.585 ;
        RECT 2912.805 2604.585 2914.015 2605.675 ;
        RECT 2912.805 2604.045 2913.325 2604.585 ;
        RECT 6.295 2601.495 6.815 2602.035 ;
        RECT 5.605 2600.405 6.815 2601.495 ;
        RECT 2906.365 2600.405 2906.655 2601.570 ;
        RECT 2912.805 2601.495 2913.325 2602.035 ;
        RECT 2909.315 2600.405 2909.645 2601.130 ;
        RECT 2912.805 2600.405 2914.015 2601.495 ;
        RECT 5.520 2600.235 6.900 2600.405 ;
        RECT 2906.300 2600.235 2906.740 2600.405 ;
        RECT 2909.040 2600.235 2910.420 2600.405 ;
        RECT 2912.720 2600.235 2914.100 2600.405 ;
        RECT 5.605 2599.145 6.815 2600.235 ;
        RECT 6.295 2598.605 6.815 2599.145 ;
        RECT 2912.805 2599.145 2914.015 2600.235 ;
        RECT 2912.805 2598.605 2913.325 2599.145 ;
        RECT 6.295 2596.055 6.815 2596.595 ;
        RECT 5.605 2594.965 6.815 2596.055 ;
        RECT 2906.365 2594.965 2906.655 2596.130 ;
        RECT 2912.805 2596.055 2913.325 2596.595 ;
        RECT 2912.805 2594.965 2914.015 2596.055 ;
        RECT 5.520 2594.795 6.900 2594.965 ;
        RECT 2906.300 2594.795 2906.740 2594.965 ;
        RECT 2912.720 2594.795 2914.100 2594.965 ;
        RECT 5.605 2593.705 6.815 2594.795 ;
        RECT 6.295 2593.165 6.815 2593.705 ;
        RECT 2912.805 2593.705 2914.015 2594.795 ;
        RECT 2912.805 2593.165 2913.325 2593.705 ;
        RECT 6.295 2590.615 6.815 2591.155 ;
        RECT 5.605 2589.525 6.815 2590.615 ;
        RECT 2906.365 2589.525 2906.655 2590.690 ;
        RECT 2912.805 2590.615 2913.325 2591.155 ;
        RECT 2912.805 2589.525 2914.015 2590.615 ;
        RECT 5.520 2589.355 6.900 2589.525 ;
        RECT 2906.300 2589.355 2906.740 2589.525 ;
        RECT 2912.720 2589.355 2914.100 2589.525 ;
        RECT 5.605 2588.265 6.815 2589.355 ;
        RECT 6.295 2587.725 6.815 2588.265 ;
        RECT 2912.805 2588.265 2914.015 2589.355 ;
        RECT 2912.805 2587.725 2913.325 2588.265 ;
        RECT 6.295 2585.175 6.815 2585.715 ;
        RECT 5.605 2584.085 6.815 2585.175 ;
        RECT 2906.365 2584.085 2906.655 2585.250 ;
        RECT 2912.805 2585.175 2913.325 2585.715 ;
        RECT 2912.805 2584.085 2914.015 2585.175 ;
        RECT 5.520 2583.915 6.900 2584.085 ;
        RECT 2906.300 2583.915 2906.740 2584.085 ;
        RECT 2912.720 2583.915 2914.100 2584.085 ;
        RECT 5.605 2582.825 6.815 2583.915 ;
        RECT 6.295 2582.285 6.815 2582.825 ;
        RECT 2912.805 2582.825 2914.015 2583.915 ;
        RECT 2912.805 2582.285 2913.325 2582.825 ;
        RECT 6.295 2579.735 6.815 2580.275 ;
        RECT 5.605 2578.645 6.815 2579.735 ;
        RECT 2906.365 2578.645 2906.655 2579.810 ;
        RECT 2912.805 2579.735 2913.325 2580.275 ;
        RECT 2912.805 2578.645 2914.015 2579.735 ;
        RECT 5.520 2578.475 6.900 2578.645 ;
        RECT 2906.300 2578.475 2906.740 2578.645 ;
        RECT 2912.720 2578.475 2914.100 2578.645 ;
        RECT 5.605 2577.385 6.815 2578.475 ;
        RECT 6.295 2576.845 6.815 2577.385 ;
        RECT 2912.805 2577.385 2914.015 2578.475 ;
        RECT 2912.805 2576.845 2913.325 2577.385 ;
        RECT 6.295 2574.295 6.815 2574.835 ;
        RECT 5.605 2573.205 6.815 2574.295 ;
        RECT 2906.365 2573.205 2906.655 2574.370 ;
        RECT 2912.805 2574.295 2913.325 2574.835 ;
        RECT 2912.805 2573.205 2914.015 2574.295 ;
        RECT 5.520 2573.035 6.900 2573.205 ;
        RECT 2906.300 2573.035 2906.740 2573.205 ;
        RECT 2912.720 2573.035 2914.100 2573.205 ;
        RECT 5.605 2571.945 6.815 2573.035 ;
        RECT 6.295 2571.405 6.815 2571.945 ;
        RECT 2912.805 2571.945 2914.015 2573.035 ;
        RECT 2912.805 2571.405 2913.325 2571.945 ;
        RECT 6.295 2568.855 6.815 2569.395 ;
        RECT 5.605 2567.765 6.815 2568.855 ;
        RECT 2906.365 2567.765 2906.655 2568.930 ;
        RECT 2912.805 2568.855 2913.325 2569.395 ;
        RECT 2912.805 2567.765 2914.015 2568.855 ;
        RECT 5.520 2567.595 6.900 2567.765 ;
        RECT 2906.300 2567.595 2906.740 2567.765 ;
        RECT 2912.720 2567.595 2914.100 2567.765 ;
        RECT 5.605 2566.505 6.815 2567.595 ;
        RECT 6.295 2565.965 6.815 2566.505 ;
        RECT 2912.805 2566.505 2914.015 2567.595 ;
        RECT 2912.805 2565.965 2913.325 2566.505 ;
        RECT 6.295 2563.415 6.815 2563.955 ;
        RECT 5.605 2562.325 6.815 2563.415 ;
        RECT 2906.365 2562.325 2906.655 2563.490 ;
        RECT 2912.805 2563.415 2913.325 2563.955 ;
        RECT 2912.805 2562.325 2914.015 2563.415 ;
        RECT 5.520 2562.155 6.900 2562.325 ;
        RECT 2906.300 2562.155 2906.740 2562.325 ;
        RECT 2912.720 2562.155 2914.100 2562.325 ;
        RECT 5.605 2561.065 6.815 2562.155 ;
        RECT 6.295 2560.525 6.815 2561.065 ;
        RECT 2912.805 2561.065 2914.015 2562.155 ;
        RECT 2912.805 2560.525 2913.325 2561.065 ;
        RECT 6.295 2557.975 6.815 2558.515 ;
        RECT 5.605 2556.885 6.815 2557.975 ;
        RECT 2906.365 2556.885 2906.655 2558.050 ;
        RECT 2912.805 2557.975 2913.325 2558.515 ;
        RECT 2912.805 2556.885 2914.015 2557.975 ;
        RECT 5.520 2556.715 6.900 2556.885 ;
        RECT 2906.300 2556.715 2906.740 2556.885 ;
        RECT 2912.720 2556.715 2914.100 2556.885 ;
        RECT 5.605 2555.625 6.815 2556.715 ;
        RECT 6.295 2555.085 6.815 2555.625 ;
        RECT 2912.805 2555.625 2914.015 2556.715 ;
        RECT 2912.805 2555.085 2913.325 2555.625 ;
        RECT 6.295 2552.535 6.815 2553.075 ;
        RECT 5.605 2551.445 6.815 2552.535 ;
        RECT 2906.365 2551.445 2906.655 2552.610 ;
        RECT 2912.805 2552.535 2913.325 2553.075 ;
        RECT 2912.805 2551.445 2914.015 2552.535 ;
        RECT 5.520 2551.275 6.900 2551.445 ;
        RECT 2906.300 2551.275 2906.740 2551.445 ;
        RECT 2912.720 2551.275 2914.100 2551.445 ;
        RECT 5.605 2550.185 6.815 2551.275 ;
        RECT 6.295 2549.645 6.815 2550.185 ;
        RECT 2912.805 2550.185 2914.015 2551.275 ;
        RECT 2912.805 2549.645 2913.325 2550.185 ;
        RECT 6.295 2547.095 6.815 2547.635 ;
        RECT 5.605 2546.005 6.815 2547.095 ;
        RECT 2906.365 2546.005 2906.655 2547.170 ;
        RECT 2912.805 2547.095 2913.325 2547.635 ;
        RECT 2912.805 2546.005 2914.015 2547.095 ;
        RECT 5.520 2545.835 6.900 2546.005 ;
        RECT 2906.300 2545.835 2906.740 2546.005 ;
        RECT 2912.720 2545.835 2914.100 2546.005 ;
        RECT 5.605 2544.745 6.815 2545.835 ;
        RECT 6.295 2544.205 6.815 2544.745 ;
        RECT 2912.805 2544.745 2914.015 2545.835 ;
        RECT 2912.805 2544.205 2913.325 2544.745 ;
        RECT 6.295 2541.655 6.815 2542.195 ;
        RECT 5.605 2540.565 6.815 2541.655 ;
        RECT 2906.365 2540.565 2906.655 2541.730 ;
        RECT 2912.805 2541.655 2913.325 2542.195 ;
        RECT 2912.805 2540.565 2914.015 2541.655 ;
        RECT 5.520 2540.395 6.900 2540.565 ;
        RECT 2906.300 2540.395 2906.740 2540.565 ;
        RECT 2912.720 2540.395 2914.100 2540.565 ;
        RECT 5.605 2539.305 6.815 2540.395 ;
        RECT 6.295 2538.765 6.815 2539.305 ;
        RECT 2912.805 2539.305 2914.015 2540.395 ;
        RECT 2912.805 2538.765 2913.325 2539.305 ;
        RECT 6.295 2536.215 6.815 2536.755 ;
        RECT 5.605 2535.125 6.815 2536.215 ;
        RECT 2906.365 2535.125 2906.655 2536.290 ;
        RECT 2912.805 2536.215 2913.325 2536.755 ;
        RECT 2912.805 2535.125 2914.015 2536.215 ;
        RECT 5.520 2534.955 6.900 2535.125 ;
        RECT 2906.300 2534.955 2906.740 2535.125 ;
        RECT 2912.720 2534.955 2914.100 2535.125 ;
        RECT 5.605 2533.865 6.815 2534.955 ;
        RECT 6.295 2533.325 6.815 2533.865 ;
        RECT 2912.805 2533.865 2914.015 2534.955 ;
        RECT 2912.805 2533.325 2913.325 2533.865 ;
        RECT 6.295 2530.775 6.815 2531.315 ;
        RECT 5.605 2529.685 6.815 2530.775 ;
        RECT 2906.365 2529.685 2906.655 2530.850 ;
        RECT 2912.805 2530.775 2913.325 2531.315 ;
        RECT 2912.805 2529.685 2914.015 2530.775 ;
        RECT 5.520 2529.515 6.900 2529.685 ;
        RECT 2906.300 2529.515 2906.740 2529.685 ;
        RECT 2912.720 2529.515 2914.100 2529.685 ;
        RECT 5.605 2528.425 6.815 2529.515 ;
        RECT 6.295 2527.885 6.815 2528.425 ;
        RECT 2912.805 2528.425 2914.015 2529.515 ;
        RECT 2912.805 2527.885 2913.325 2528.425 ;
        RECT 6.295 2525.335 6.815 2525.875 ;
        RECT 5.605 2524.245 6.815 2525.335 ;
        RECT 2906.365 2524.245 2906.655 2525.410 ;
        RECT 2912.805 2525.335 2913.325 2525.875 ;
        RECT 2912.805 2524.245 2914.015 2525.335 ;
        RECT 5.520 2524.075 6.900 2524.245 ;
        RECT 2906.300 2524.075 2906.740 2524.245 ;
        RECT 2912.720 2524.075 2914.100 2524.245 ;
        RECT 5.605 2522.985 6.815 2524.075 ;
        RECT 6.295 2522.445 6.815 2522.985 ;
        RECT 2912.805 2522.985 2914.015 2524.075 ;
        RECT 2912.805 2522.445 2913.325 2522.985 ;
        RECT 6.295 2519.895 6.815 2520.435 ;
        RECT 5.605 2518.805 6.815 2519.895 ;
        RECT 2906.365 2518.805 2906.655 2519.970 ;
        RECT 2912.805 2519.895 2913.325 2520.435 ;
        RECT 2912.805 2518.805 2914.015 2519.895 ;
        RECT 5.520 2518.635 6.900 2518.805 ;
        RECT 2906.300 2518.635 2906.740 2518.805 ;
        RECT 2912.720 2518.635 2914.100 2518.805 ;
        RECT 5.605 2517.545 6.815 2518.635 ;
        RECT 6.295 2517.005 6.815 2517.545 ;
        RECT 2912.805 2517.545 2914.015 2518.635 ;
        RECT 2912.805 2517.005 2913.325 2517.545 ;
        RECT 6.295 2514.455 6.815 2514.995 ;
        RECT 5.605 2513.365 6.815 2514.455 ;
        RECT 2906.365 2513.365 2906.655 2514.530 ;
        RECT 2912.805 2514.455 2913.325 2514.995 ;
        RECT 2912.805 2513.365 2914.015 2514.455 ;
        RECT 5.520 2513.195 6.900 2513.365 ;
        RECT 2906.300 2513.195 2906.740 2513.365 ;
        RECT 2912.720 2513.195 2914.100 2513.365 ;
        RECT 5.605 2512.105 6.815 2513.195 ;
        RECT 6.295 2511.565 6.815 2512.105 ;
        RECT 2912.805 2512.105 2914.015 2513.195 ;
        RECT 2912.805 2511.565 2913.325 2512.105 ;
        RECT 6.295 2509.015 6.815 2509.555 ;
        RECT 5.605 2507.925 6.815 2509.015 ;
        RECT 2906.365 2507.925 2906.655 2509.090 ;
        RECT 2912.805 2509.015 2913.325 2509.555 ;
        RECT 2912.805 2507.925 2914.015 2509.015 ;
        RECT 5.520 2507.755 6.900 2507.925 ;
        RECT 2906.300 2507.755 2906.740 2507.925 ;
        RECT 2912.720 2507.755 2914.100 2507.925 ;
        RECT 5.605 2506.665 6.815 2507.755 ;
        RECT 6.295 2506.125 6.815 2506.665 ;
        RECT 2912.805 2506.665 2914.015 2507.755 ;
        RECT 2912.805 2506.125 2913.325 2506.665 ;
        RECT 6.295 2503.575 6.815 2504.115 ;
        RECT 5.605 2502.485 6.815 2503.575 ;
        RECT 2906.365 2502.485 2906.655 2503.650 ;
        RECT 2912.805 2503.575 2913.325 2504.115 ;
        RECT 2912.805 2502.485 2914.015 2503.575 ;
        RECT 5.520 2502.315 6.900 2502.485 ;
        RECT 8.740 2502.315 10.120 2502.485 ;
        RECT 2906.300 2502.315 2906.740 2502.485 ;
        RECT 2912.720 2502.315 2914.100 2502.485 ;
        RECT 5.605 2501.225 6.815 2502.315 ;
        RECT 9.015 2501.590 9.345 2502.315 ;
        RECT 6.295 2500.685 6.815 2501.225 ;
        RECT 2912.805 2501.225 2914.015 2502.315 ;
        RECT 2912.805 2500.685 2913.325 2501.225 ;
        RECT 6.295 2498.135 6.815 2498.675 ;
        RECT 5.605 2497.045 6.815 2498.135 ;
        RECT 2906.365 2497.045 2906.655 2498.210 ;
        RECT 2912.805 2498.135 2913.325 2498.675 ;
        RECT 2912.805 2497.045 2914.015 2498.135 ;
        RECT 5.520 2496.875 6.900 2497.045 ;
        RECT 2906.300 2496.875 2906.740 2497.045 ;
        RECT 2912.720 2496.875 2914.100 2497.045 ;
        RECT 5.605 2495.785 6.815 2496.875 ;
        RECT 6.295 2495.245 6.815 2495.785 ;
        RECT 2912.805 2495.785 2914.015 2496.875 ;
        RECT 2912.805 2495.245 2913.325 2495.785 ;
        RECT 6.295 2492.695 6.815 2493.235 ;
        RECT 5.605 2491.605 6.815 2492.695 ;
        RECT 2906.365 2491.605 2906.655 2492.770 ;
        RECT 2912.805 2492.695 2913.325 2493.235 ;
        RECT 2912.805 2491.605 2914.015 2492.695 ;
        RECT 5.520 2491.435 6.900 2491.605 ;
        RECT 2906.300 2491.435 2906.740 2491.605 ;
        RECT 2912.720 2491.435 2914.100 2491.605 ;
        RECT 5.605 2490.345 6.815 2491.435 ;
        RECT 6.295 2489.805 6.815 2490.345 ;
        RECT 2912.805 2490.345 2914.015 2491.435 ;
        RECT 2912.805 2489.805 2913.325 2490.345 ;
        RECT 6.295 2487.255 6.815 2487.795 ;
        RECT 5.605 2486.165 6.815 2487.255 ;
        RECT 2906.365 2486.165 2906.655 2487.330 ;
        RECT 2912.805 2487.255 2913.325 2487.795 ;
        RECT 2912.805 2486.165 2914.015 2487.255 ;
        RECT 5.520 2485.995 6.900 2486.165 ;
        RECT 2906.300 2485.995 2906.740 2486.165 ;
        RECT 2912.720 2485.995 2914.100 2486.165 ;
        RECT 5.605 2484.905 6.815 2485.995 ;
        RECT 6.295 2484.365 6.815 2484.905 ;
        RECT 2912.805 2484.905 2914.015 2485.995 ;
        RECT 2912.805 2484.365 2913.325 2484.905 ;
        RECT 6.295 2481.815 6.815 2482.355 ;
        RECT 5.605 2480.725 6.815 2481.815 ;
        RECT 2906.365 2480.725 2906.655 2481.890 ;
        RECT 2912.805 2481.815 2913.325 2482.355 ;
        RECT 2912.805 2480.725 2914.015 2481.815 ;
        RECT 5.520 2480.555 6.900 2480.725 ;
        RECT 2906.300 2480.555 2906.740 2480.725 ;
        RECT 2912.720 2480.555 2914.100 2480.725 ;
        RECT 5.605 2479.465 6.815 2480.555 ;
        RECT 6.295 2478.925 6.815 2479.465 ;
        RECT 2912.805 2479.465 2914.015 2480.555 ;
        RECT 2912.805 2478.925 2913.325 2479.465 ;
        RECT 6.295 2476.375 6.815 2476.915 ;
        RECT 5.605 2475.285 6.815 2476.375 ;
        RECT 2906.365 2475.285 2906.655 2476.450 ;
        RECT 2912.805 2476.375 2913.325 2476.915 ;
        RECT 2912.805 2475.285 2914.015 2476.375 ;
        RECT 5.520 2475.115 6.900 2475.285 ;
        RECT 2906.300 2475.115 2906.740 2475.285 ;
        RECT 2912.720 2475.115 2914.100 2475.285 ;
        RECT 5.605 2474.025 6.815 2475.115 ;
        RECT 6.295 2473.485 6.815 2474.025 ;
        RECT 2912.805 2474.025 2914.015 2475.115 ;
        RECT 2912.805 2473.485 2913.325 2474.025 ;
        RECT 6.295 2470.935 6.815 2471.475 ;
        RECT 5.605 2469.845 6.815 2470.935 ;
        RECT 2906.365 2469.845 2906.655 2471.010 ;
        RECT 2912.805 2470.935 2913.325 2471.475 ;
        RECT 2912.805 2469.845 2914.015 2470.935 ;
        RECT 5.520 2469.675 6.900 2469.845 ;
        RECT 2906.300 2469.675 2906.740 2469.845 ;
        RECT 2912.720 2469.675 2914.100 2469.845 ;
        RECT 5.605 2468.585 6.815 2469.675 ;
        RECT 6.295 2468.045 6.815 2468.585 ;
        RECT 2912.805 2468.585 2914.015 2469.675 ;
        RECT 2912.805 2468.045 2913.325 2468.585 ;
        RECT 6.295 2465.495 6.815 2466.035 ;
        RECT 5.605 2464.405 6.815 2465.495 ;
        RECT 2906.365 2464.405 2906.655 2465.570 ;
        RECT 2912.805 2465.495 2913.325 2466.035 ;
        RECT 2912.805 2464.405 2914.015 2465.495 ;
        RECT 5.520 2464.235 6.900 2464.405 ;
        RECT 2906.300 2464.235 2906.740 2464.405 ;
        RECT 2909.040 2464.235 2910.420 2464.405 ;
        RECT 2912.720 2464.235 2914.100 2464.405 ;
        RECT 5.605 2463.145 6.815 2464.235 ;
        RECT 2909.315 2463.510 2909.645 2464.235 ;
        RECT 6.295 2462.605 6.815 2463.145 ;
        RECT 2912.805 2463.145 2914.015 2464.235 ;
        RECT 2912.805 2462.605 2913.325 2463.145 ;
        RECT 6.295 2460.055 6.815 2460.595 ;
        RECT 5.605 2458.965 6.815 2460.055 ;
        RECT 2906.365 2458.965 2906.655 2460.130 ;
        RECT 2912.805 2460.055 2913.325 2460.595 ;
        RECT 2912.805 2458.965 2914.015 2460.055 ;
        RECT 5.520 2458.795 6.900 2458.965 ;
        RECT 2906.300 2458.795 2906.740 2458.965 ;
        RECT 2912.720 2458.795 2914.100 2458.965 ;
        RECT 5.605 2457.705 6.815 2458.795 ;
        RECT 6.295 2457.165 6.815 2457.705 ;
        RECT 2912.805 2457.705 2914.015 2458.795 ;
        RECT 2912.805 2457.165 2913.325 2457.705 ;
        RECT 6.295 2454.615 6.815 2455.155 ;
        RECT 5.605 2453.525 6.815 2454.615 ;
        RECT 2906.365 2453.525 2906.655 2454.690 ;
        RECT 2912.805 2454.615 2913.325 2455.155 ;
        RECT 2912.805 2453.525 2914.015 2454.615 ;
        RECT 5.520 2453.355 6.900 2453.525 ;
        RECT 2906.300 2453.355 2906.740 2453.525 ;
        RECT 2912.720 2453.355 2914.100 2453.525 ;
        RECT 5.605 2452.265 6.815 2453.355 ;
        RECT 6.295 2451.725 6.815 2452.265 ;
        RECT 2912.805 2452.265 2914.015 2453.355 ;
        RECT 2912.805 2451.725 2913.325 2452.265 ;
        RECT 6.295 2449.175 6.815 2449.715 ;
        RECT 5.605 2448.085 6.815 2449.175 ;
        RECT 2906.365 2448.085 2906.655 2449.250 ;
        RECT 2912.805 2449.175 2913.325 2449.715 ;
        RECT 2912.805 2448.085 2914.015 2449.175 ;
        RECT 5.520 2447.915 6.900 2448.085 ;
        RECT 2906.300 2447.915 2906.740 2448.085 ;
        RECT 2912.720 2447.915 2914.100 2448.085 ;
        RECT 5.605 2446.825 6.815 2447.915 ;
        RECT 6.295 2446.285 6.815 2446.825 ;
        RECT 2912.805 2446.825 2914.015 2447.915 ;
        RECT 2912.805 2446.285 2913.325 2446.825 ;
        RECT 6.295 2443.735 6.815 2444.275 ;
        RECT 5.605 2442.645 6.815 2443.735 ;
        RECT 2906.365 2442.645 2906.655 2443.810 ;
        RECT 2912.805 2443.735 2913.325 2444.275 ;
        RECT 2912.805 2442.645 2914.015 2443.735 ;
        RECT 5.520 2442.475 6.900 2442.645 ;
        RECT 2906.300 2442.475 2906.740 2442.645 ;
        RECT 2912.720 2442.475 2914.100 2442.645 ;
        RECT 5.605 2441.385 6.815 2442.475 ;
        RECT 6.295 2440.845 6.815 2441.385 ;
        RECT 2912.805 2441.385 2914.015 2442.475 ;
        RECT 2912.805 2440.845 2913.325 2441.385 ;
        RECT 6.295 2438.295 6.815 2438.835 ;
        RECT 5.605 2437.205 6.815 2438.295 ;
        RECT 2906.365 2437.205 2906.655 2438.370 ;
        RECT 2912.805 2438.295 2913.325 2438.835 ;
        RECT 2912.805 2437.205 2914.015 2438.295 ;
        RECT 5.520 2437.035 6.900 2437.205 ;
        RECT 2906.300 2437.035 2906.740 2437.205 ;
        RECT 2912.720 2437.035 2914.100 2437.205 ;
        RECT 5.605 2435.945 6.815 2437.035 ;
        RECT 6.295 2435.405 6.815 2435.945 ;
        RECT 2912.805 2435.945 2914.015 2437.035 ;
        RECT 2912.805 2435.405 2913.325 2435.945 ;
        RECT 6.295 2432.855 6.815 2433.395 ;
        RECT 5.605 2431.765 6.815 2432.855 ;
        RECT 2906.365 2431.765 2906.655 2432.930 ;
        RECT 2912.805 2432.855 2913.325 2433.395 ;
        RECT 2909.315 2431.765 2909.645 2432.490 ;
        RECT 2912.805 2431.765 2914.015 2432.855 ;
        RECT 5.520 2431.595 6.900 2431.765 ;
        RECT 2906.300 2431.595 2906.740 2431.765 ;
        RECT 2909.040 2431.595 2910.420 2431.765 ;
        RECT 2912.720 2431.595 2914.100 2431.765 ;
        RECT 5.605 2430.505 6.815 2431.595 ;
        RECT 6.295 2429.965 6.815 2430.505 ;
        RECT 2912.805 2430.505 2914.015 2431.595 ;
        RECT 2912.805 2429.965 2913.325 2430.505 ;
        RECT 6.295 2427.415 6.815 2427.955 ;
        RECT 5.605 2426.325 6.815 2427.415 ;
        RECT 2906.365 2426.325 2906.655 2427.490 ;
        RECT 2912.805 2427.415 2913.325 2427.955 ;
        RECT 2912.805 2426.325 2914.015 2427.415 ;
        RECT 5.520 2426.155 6.900 2426.325 ;
        RECT 2906.300 2426.155 2906.740 2426.325 ;
        RECT 2912.720 2426.155 2914.100 2426.325 ;
        RECT 5.605 2425.065 6.815 2426.155 ;
        RECT 6.295 2424.525 6.815 2425.065 ;
        RECT 2912.805 2425.065 2914.015 2426.155 ;
        RECT 2912.805 2424.525 2913.325 2425.065 ;
        RECT 6.295 2421.975 6.815 2422.515 ;
        RECT 5.605 2420.885 6.815 2421.975 ;
        RECT 2906.365 2420.885 2906.655 2422.050 ;
        RECT 2912.805 2421.975 2913.325 2422.515 ;
        RECT 2912.805 2420.885 2914.015 2421.975 ;
        RECT 5.520 2420.715 6.900 2420.885 ;
        RECT 2906.300 2420.715 2906.740 2420.885 ;
        RECT 2912.720 2420.715 2914.100 2420.885 ;
        RECT 5.605 2419.625 6.815 2420.715 ;
        RECT 6.295 2419.085 6.815 2419.625 ;
        RECT 2912.805 2419.625 2914.015 2420.715 ;
        RECT 2912.805 2419.085 2913.325 2419.625 ;
        RECT 6.295 2416.535 6.815 2417.075 ;
        RECT 5.605 2415.445 6.815 2416.535 ;
        RECT 2906.365 2415.445 2906.655 2416.610 ;
        RECT 2912.805 2416.535 2913.325 2417.075 ;
        RECT 2912.805 2415.445 2914.015 2416.535 ;
        RECT 5.520 2415.275 6.900 2415.445 ;
        RECT 2906.300 2415.275 2906.740 2415.445 ;
        RECT 2912.720 2415.275 2914.100 2415.445 ;
        RECT 5.605 2414.185 6.815 2415.275 ;
        RECT 6.295 2413.645 6.815 2414.185 ;
        RECT 2912.805 2414.185 2914.015 2415.275 ;
        RECT 2912.805 2413.645 2913.325 2414.185 ;
        RECT 6.295 2411.095 6.815 2411.635 ;
        RECT 5.605 2410.005 6.815 2411.095 ;
        RECT 2906.365 2410.005 2906.655 2411.170 ;
        RECT 2912.805 2411.095 2913.325 2411.635 ;
        RECT 2912.805 2410.005 2914.015 2411.095 ;
        RECT 5.520 2409.835 6.900 2410.005 ;
        RECT 2906.300 2409.835 2906.740 2410.005 ;
        RECT 2912.720 2409.835 2914.100 2410.005 ;
        RECT 5.605 2408.745 6.815 2409.835 ;
        RECT 6.295 2408.205 6.815 2408.745 ;
        RECT 2912.805 2408.745 2914.015 2409.835 ;
        RECT 2912.805 2408.205 2913.325 2408.745 ;
        RECT 6.295 2405.655 6.815 2406.195 ;
        RECT 5.605 2404.565 6.815 2405.655 ;
        RECT 2906.365 2404.565 2906.655 2405.730 ;
        RECT 2912.805 2405.655 2913.325 2406.195 ;
        RECT 2912.805 2404.565 2914.015 2405.655 ;
        RECT 5.520 2404.395 6.900 2404.565 ;
        RECT 2906.300 2404.395 2906.740 2404.565 ;
        RECT 2912.720 2404.395 2914.100 2404.565 ;
        RECT 5.605 2403.305 6.815 2404.395 ;
        RECT 6.295 2402.765 6.815 2403.305 ;
        RECT 2912.805 2403.305 2914.015 2404.395 ;
        RECT 2912.805 2402.765 2913.325 2403.305 ;
        RECT 6.295 2400.215 6.815 2400.755 ;
        RECT 5.605 2399.125 6.815 2400.215 ;
        RECT 2906.365 2399.125 2906.655 2400.290 ;
        RECT 2912.805 2400.215 2913.325 2400.755 ;
        RECT 2912.805 2399.125 2914.015 2400.215 ;
        RECT 5.520 2398.955 6.900 2399.125 ;
        RECT 2906.300 2398.955 2906.740 2399.125 ;
        RECT 2912.720 2398.955 2914.100 2399.125 ;
        RECT 5.605 2397.865 6.815 2398.955 ;
        RECT 6.295 2397.325 6.815 2397.865 ;
        RECT 2912.805 2397.865 2914.015 2398.955 ;
        RECT 2912.805 2397.325 2913.325 2397.865 ;
        RECT 6.295 2394.775 6.815 2395.315 ;
        RECT 5.605 2393.685 6.815 2394.775 ;
        RECT 2906.365 2393.685 2906.655 2394.850 ;
        RECT 2912.805 2394.775 2913.325 2395.315 ;
        RECT 2912.805 2393.685 2914.015 2394.775 ;
        RECT 5.520 2393.515 6.900 2393.685 ;
        RECT 2906.300 2393.515 2906.740 2393.685 ;
        RECT 2912.720 2393.515 2914.100 2393.685 ;
        RECT 5.605 2392.425 6.815 2393.515 ;
        RECT 6.295 2391.885 6.815 2392.425 ;
        RECT 2912.805 2392.425 2914.015 2393.515 ;
        RECT 2912.805 2391.885 2913.325 2392.425 ;
        RECT 6.295 2389.335 6.815 2389.875 ;
        RECT 5.605 2388.245 6.815 2389.335 ;
        RECT 2906.365 2388.245 2906.655 2389.410 ;
        RECT 2912.805 2389.335 2913.325 2389.875 ;
        RECT 2912.805 2388.245 2914.015 2389.335 ;
        RECT 5.520 2388.075 6.900 2388.245 ;
        RECT 2906.300 2388.075 2906.740 2388.245 ;
        RECT 2909.040 2388.075 2910.420 2388.245 ;
        RECT 2912.720 2388.075 2914.100 2388.245 ;
        RECT 5.605 2386.985 6.815 2388.075 ;
        RECT 2909.315 2387.350 2909.645 2388.075 ;
        RECT 6.295 2386.445 6.815 2386.985 ;
        RECT 2912.805 2386.985 2914.015 2388.075 ;
        RECT 2912.805 2386.445 2913.325 2386.985 ;
        RECT 6.295 2383.895 6.815 2384.435 ;
        RECT 5.605 2382.805 6.815 2383.895 ;
        RECT 2906.365 2382.805 2906.655 2383.970 ;
        RECT 2912.805 2383.895 2913.325 2384.435 ;
        RECT 2912.805 2382.805 2914.015 2383.895 ;
        RECT 5.520 2382.635 6.900 2382.805 ;
        RECT 8.740 2382.635 10.120 2382.805 ;
        RECT 2906.300 2382.635 2906.740 2382.805 ;
        RECT 2912.720 2382.635 2914.100 2382.805 ;
        RECT 5.605 2381.545 6.815 2382.635 ;
        RECT 9.015 2381.910 9.345 2382.635 ;
        RECT 6.295 2381.005 6.815 2381.545 ;
        RECT 2912.805 2381.545 2914.015 2382.635 ;
        RECT 2912.805 2381.005 2913.325 2381.545 ;
        RECT 6.295 2378.455 6.815 2378.995 ;
        RECT 5.605 2377.365 6.815 2378.455 ;
        RECT 2906.365 2377.365 2906.655 2378.530 ;
        RECT 2912.805 2378.455 2913.325 2378.995 ;
        RECT 2912.805 2377.365 2914.015 2378.455 ;
        RECT 5.520 2377.195 6.900 2377.365 ;
        RECT 2906.300 2377.195 2906.740 2377.365 ;
        RECT 2912.720 2377.195 2914.100 2377.365 ;
        RECT 5.605 2376.105 6.815 2377.195 ;
        RECT 6.295 2375.565 6.815 2376.105 ;
        RECT 2912.805 2376.105 2914.015 2377.195 ;
        RECT 2912.805 2375.565 2913.325 2376.105 ;
        RECT 6.295 2373.015 6.815 2373.555 ;
        RECT 5.605 2371.925 6.815 2373.015 ;
        RECT 2906.365 2371.925 2906.655 2373.090 ;
        RECT 2912.805 2373.015 2913.325 2373.555 ;
        RECT 2912.805 2371.925 2914.015 2373.015 ;
        RECT 5.520 2371.755 6.900 2371.925 ;
        RECT 2906.300 2371.755 2906.740 2371.925 ;
        RECT 2912.720 2371.755 2914.100 2371.925 ;
        RECT 5.605 2370.665 6.815 2371.755 ;
        RECT 6.295 2370.125 6.815 2370.665 ;
        RECT 2912.805 2370.665 2914.015 2371.755 ;
        RECT 2912.805 2370.125 2913.325 2370.665 ;
        RECT 6.295 2367.575 6.815 2368.115 ;
        RECT 5.605 2366.485 6.815 2367.575 ;
        RECT 2906.365 2366.485 2906.655 2367.650 ;
        RECT 2912.805 2367.575 2913.325 2368.115 ;
        RECT 2912.805 2366.485 2914.015 2367.575 ;
        RECT 5.520 2366.315 6.900 2366.485 ;
        RECT 2906.300 2366.315 2906.740 2366.485 ;
        RECT 2912.720 2366.315 2914.100 2366.485 ;
        RECT 5.605 2365.225 6.815 2366.315 ;
        RECT 6.295 2364.685 6.815 2365.225 ;
        RECT 2912.805 2365.225 2914.015 2366.315 ;
        RECT 2912.805 2364.685 2913.325 2365.225 ;
        RECT 6.295 2362.135 6.815 2362.675 ;
        RECT 5.605 2361.045 6.815 2362.135 ;
        RECT 2906.365 2361.045 2906.655 2362.210 ;
        RECT 2912.805 2362.135 2913.325 2362.675 ;
        RECT 2912.805 2361.045 2914.015 2362.135 ;
        RECT 5.520 2360.875 6.900 2361.045 ;
        RECT 2906.300 2360.875 2906.740 2361.045 ;
        RECT 2912.720 2360.875 2914.100 2361.045 ;
        RECT 5.605 2359.785 6.815 2360.875 ;
        RECT 6.295 2359.245 6.815 2359.785 ;
        RECT 2912.805 2359.785 2914.015 2360.875 ;
        RECT 2912.805 2359.245 2913.325 2359.785 ;
        RECT 6.295 2356.695 6.815 2357.235 ;
        RECT 5.605 2355.605 6.815 2356.695 ;
        RECT 2906.365 2355.605 2906.655 2356.770 ;
        RECT 2912.805 2356.695 2913.325 2357.235 ;
        RECT 2912.805 2355.605 2914.015 2356.695 ;
        RECT 5.520 2355.435 6.900 2355.605 ;
        RECT 2906.300 2355.435 2906.740 2355.605 ;
        RECT 2912.720 2355.435 2914.100 2355.605 ;
        RECT 5.605 2354.345 6.815 2355.435 ;
        RECT 6.295 2353.805 6.815 2354.345 ;
        RECT 2912.805 2354.345 2914.015 2355.435 ;
        RECT 2912.805 2353.805 2913.325 2354.345 ;
        RECT 6.295 2351.255 6.815 2351.795 ;
        RECT 5.605 2350.165 6.815 2351.255 ;
        RECT 2906.365 2350.165 2906.655 2351.330 ;
        RECT 2912.805 2351.255 2913.325 2351.795 ;
        RECT 2912.805 2350.165 2914.015 2351.255 ;
        RECT 5.520 2349.995 6.900 2350.165 ;
        RECT 2906.300 2349.995 2906.740 2350.165 ;
        RECT 2912.720 2349.995 2914.100 2350.165 ;
        RECT 5.605 2348.905 6.815 2349.995 ;
        RECT 6.295 2348.365 6.815 2348.905 ;
        RECT 2912.805 2348.905 2914.015 2349.995 ;
        RECT 2912.805 2348.365 2913.325 2348.905 ;
        RECT 6.295 2345.815 6.815 2346.355 ;
        RECT 5.605 2344.725 6.815 2345.815 ;
        RECT 2906.365 2344.725 2906.655 2345.890 ;
        RECT 2912.805 2345.815 2913.325 2346.355 ;
        RECT 2912.805 2344.725 2914.015 2345.815 ;
        RECT 5.520 2344.555 6.900 2344.725 ;
        RECT 2906.300 2344.555 2906.740 2344.725 ;
        RECT 2912.720 2344.555 2914.100 2344.725 ;
        RECT 5.605 2343.465 6.815 2344.555 ;
        RECT 6.295 2342.925 6.815 2343.465 ;
        RECT 2912.805 2343.465 2914.015 2344.555 ;
        RECT 2912.805 2342.925 2913.325 2343.465 ;
        RECT 6.295 2340.375 6.815 2340.915 ;
        RECT 5.605 2339.285 6.815 2340.375 ;
        RECT 2906.365 2339.285 2906.655 2340.450 ;
        RECT 2912.805 2340.375 2913.325 2340.915 ;
        RECT 2912.805 2339.285 2914.015 2340.375 ;
        RECT 5.520 2339.115 6.900 2339.285 ;
        RECT 2906.300 2339.115 2906.740 2339.285 ;
        RECT 2912.720 2339.115 2914.100 2339.285 ;
        RECT 5.605 2338.025 6.815 2339.115 ;
        RECT 6.295 2337.485 6.815 2338.025 ;
        RECT 2912.805 2338.025 2914.015 2339.115 ;
        RECT 2912.805 2337.485 2913.325 2338.025 ;
        RECT 6.295 2334.935 6.815 2335.475 ;
        RECT 5.605 2333.845 6.815 2334.935 ;
        RECT 2906.365 2333.845 2906.655 2335.010 ;
        RECT 2912.805 2334.935 2913.325 2335.475 ;
        RECT 2912.805 2333.845 2914.015 2334.935 ;
        RECT 5.520 2333.675 6.900 2333.845 ;
        RECT 2906.300 2333.675 2906.740 2333.845 ;
        RECT 2912.720 2333.675 2914.100 2333.845 ;
        RECT 5.605 2332.585 6.815 2333.675 ;
        RECT 6.295 2332.045 6.815 2332.585 ;
        RECT 2912.805 2332.585 2914.015 2333.675 ;
        RECT 2912.805 2332.045 2913.325 2332.585 ;
        RECT 6.295 2329.495 6.815 2330.035 ;
        RECT 5.605 2328.405 6.815 2329.495 ;
        RECT 2906.365 2328.405 2906.655 2329.570 ;
        RECT 2912.805 2329.495 2913.325 2330.035 ;
        RECT 2912.805 2328.405 2914.015 2329.495 ;
        RECT 5.520 2328.235 6.900 2328.405 ;
        RECT 2906.300 2328.235 2906.740 2328.405 ;
        RECT 2912.720 2328.235 2914.100 2328.405 ;
        RECT 5.605 2327.145 6.815 2328.235 ;
        RECT 6.295 2326.605 6.815 2327.145 ;
        RECT 2912.805 2327.145 2914.015 2328.235 ;
        RECT 2912.805 2326.605 2913.325 2327.145 ;
        RECT 6.295 2324.055 6.815 2324.595 ;
        RECT 5.605 2322.965 6.815 2324.055 ;
        RECT 2906.365 2322.965 2906.655 2324.130 ;
        RECT 2912.805 2324.055 2913.325 2324.595 ;
        RECT 2912.805 2322.965 2914.015 2324.055 ;
        RECT 5.520 2322.795 6.900 2322.965 ;
        RECT 2906.300 2322.795 2906.740 2322.965 ;
        RECT 2912.720 2322.795 2914.100 2322.965 ;
        RECT 5.605 2321.705 6.815 2322.795 ;
        RECT 6.295 2321.165 6.815 2321.705 ;
        RECT 2912.805 2321.705 2914.015 2322.795 ;
        RECT 2912.805 2321.165 2913.325 2321.705 ;
        RECT 6.295 2318.615 6.815 2319.155 ;
        RECT 5.605 2317.525 6.815 2318.615 ;
        RECT 2906.365 2317.525 2906.655 2318.690 ;
        RECT 2912.805 2318.615 2913.325 2319.155 ;
        RECT 2912.805 2317.525 2914.015 2318.615 ;
        RECT 5.520 2317.355 6.900 2317.525 ;
        RECT 2906.300 2317.355 2906.740 2317.525 ;
        RECT 2912.720 2317.355 2914.100 2317.525 ;
        RECT 5.605 2316.265 6.815 2317.355 ;
        RECT 6.295 2315.725 6.815 2316.265 ;
        RECT 2912.805 2316.265 2914.015 2317.355 ;
        RECT 2912.805 2315.725 2913.325 2316.265 ;
        RECT 6.295 2313.175 6.815 2313.715 ;
        RECT 5.605 2312.085 6.815 2313.175 ;
        RECT 2906.365 2312.085 2906.655 2313.250 ;
        RECT 2912.805 2313.175 2913.325 2313.715 ;
        RECT 2912.805 2312.085 2914.015 2313.175 ;
        RECT 5.520 2311.915 6.900 2312.085 ;
        RECT 2906.300 2311.915 2906.740 2312.085 ;
        RECT 2912.720 2311.915 2914.100 2312.085 ;
        RECT 5.605 2310.825 6.815 2311.915 ;
        RECT 6.295 2310.285 6.815 2310.825 ;
        RECT 2912.805 2310.825 2914.015 2311.915 ;
        RECT 2912.805 2310.285 2913.325 2310.825 ;
        RECT 6.295 2307.735 6.815 2308.275 ;
        RECT 5.605 2306.645 6.815 2307.735 ;
        RECT 2906.365 2306.645 2906.655 2307.810 ;
        RECT 2912.805 2307.735 2913.325 2308.275 ;
        RECT 2912.805 2306.645 2914.015 2307.735 ;
        RECT 5.520 2306.475 6.900 2306.645 ;
        RECT 2906.300 2306.475 2906.740 2306.645 ;
        RECT 2912.720 2306.475 2914.100 2306.645 ;
        RECT 5.605 2305.385 6.815 2306.475 ;
        RECT 6.295 2304.845 6.815 2305.385 ;
        RECT 2912.805 2305.385 2914.015 2306.475 ;
        RECT 2912.805 2304.845 2913.325 2305.385 ;
        RECT 6.295 2302.295 6.815 2302.835 ;
        RECT 5.605 2301.205 6.815 2302.295 ;
        RECT 2906.365 2301.205 2906.655 2302.370 ;
        RECT 2912.805 2302.295 2913.325 2302.835 ;
        RECT 2912.805 2301.205 2914.015 2302.295 ;
        RECT 5.520 2301.035 6.900 2301.205 ;
        RECT 2906.300 2301.035 2906.740 2301.205 ;
        RECT 2912.720 2301.035 2914.100 2301.205 ;
        RECT 5.605 2299.945 6.815 2301.035 ;
        RECT 6.295 2299.405 6.815 2299.945 ;
        RECT 2912.805 2299.945 2914.015 2301.035 ;
        RECT 2912.805 2299.405 2913.325 2299.945 ;
        RECT 6.295 2296.855 6.815 2297.395 ;
        RECT 5.605 2295.765 6.815 2296.855 ;
        RECT 2906.365 2295.765 2906.655 2296.930 ;
        RECT 2912.805 2296.855 2913.325 2297.395 ;
        RECT 2912.805 2295.765 2914.015 2296.855 ;
        RECT 5.520 2295.595 6.900 2295.765 ;
        RECT 2906.300 2295.595 2906.740 2295.765 ;
        RECT 2912.720 2295.595 2914.100 2295.765 ;
        RECT 5.605 2294.505 6.815 2295.595 ;
        RECT 6.295 2293.965 6.815 2294.505 ;
        RECT 2912.805 2294.505 2914.015 2295.595 ;
        RECT 2912.805 2293.965 2913.325 2294.505 ;
        RECT 6.295 2291.415 6.815 2291.955 ;
        RECT 5.605 2290.325 6.815 2291.415 ;
        RECT 2906.365 2290.325 2906.655 2291.490 ;
        RECT 2912.805 2291.415 2913.325 2291.955 ;
        RECT 2912.805 2290.325 2914.015 2291.415 ;
        RECT 5.520 2290.155 6.900 2290.325 ;
        RECT 2906.300 2290.155 2906.740 2290.325 ;
        RECT 2912.720 2290.155 2914.100 2290.325 ;
        RECT 5.605 2289.065 6.815 2290.155 ;
        RECT 6.295 2288.525 6.815 2289.065 ;
        RECT 2912.805 2289.065 2914.015 2290.155 ;
        RECT 2912.805 2288.525 2913.325 2289.065 ;
        RECT 6.295 2285.975 6.815 2286.515 ;
        RECT 5.605 2284.885 6.815 2285.975 ;
        RECT 2906.365 2284.885 2906.655 2286.050 ;
        RECT 2912.805 2285.975 2913.325 2286.515 ;
        RECT 2912.805 2284.885 2914.015 2285.975 ;
        RECT 5.520 2284.715 6.900 2284.885 ;
        RECT 2906.300 2284.715 2906.740 2284.885 ;
        RECT 2912.720 2284.715 2914.100 2284.885 ;
        RECT 5.605 2283.625 6.815 2284.715 ;
        RECT 6.295 2283.085 6.815 2283.625 ;
        RECT 2912.805 2283.625 2914.015 2284.715 ;
        RECT 2912.805 2283.085 2913.325 2283.625 ;
        RECT 6.295 2280.535 6.815 2281.075 ;
        RECT 5.605 2279.445 6.815 2280.535 ;
        RECT 2906.365 2279.445 2906.655 2280.610 ;
        RECT 2912.805 2280.535 2913.325 2281.075 ;
        RECT 2912.805 2279.445 2914.015 2280.535 ;
        RECT 5.520 2279.275 6.900 2279.445 ;
        RECT 2906.300 2279.275 2906.740 2279.445 ;
        RECT 2912.720 2279.275 2914.100 2279.445 ;
        RECT 5.605 2278.185 6.815 2279.275 ;
        RECT 6.295 2277.645 6.815 2278.185 ;
        RECT 2912.805 2278.185 2914.015 2279.275 ;
        RECT 2912.805 2277.645 2913.325 2278.185 ;
        RECT 6.295 2275.095 6.815 2275.635 ;
        RECT 5.605 2274.005 6.815 2275.095 ;
        RECT 2906.365 2274.005 2906.655 2275.170 ;
        RECT 2912.805 2275.095 2913.325 2275.635 ;
        RECT 2912.805 2274.005 2914.015 2275.095 ;
        RECT 5.520 2273.835 6.900 2274.005 ;
        RECT 2906.300 2273.835 2906.740 2274.005 ;
        RECT 2912.720 2273.835 2914.100 2274.005 ;
        RECT 5.605 2272.745 6.815 2273.835 ;
        RECT 6.295 2272.205 6.815 2272.745 ;
        RECT 2912.805 2272.745 2914.015 2273.835 ;
        RECT 2912.805 2272.205 2913.325 2272.745 ;
        RECT 6.295 2269.655 6.815 2270.195 ;
        RECT 5.605 2268.565 6.815 2269.655 ;
        RECT 2906.365 2268.565 2906.655 2269.730 ;
        RECT 2912.805 2269.655 2913.325 2270.195 ;
        RECT 2912.805 2268.565 2914.015 2269.655 ;
        RECT 5.520 2268.395 6.900 2268.565 ;
        RECT 2906.300 2268.395 2906.740 2268.565 ;
        RECT 2912.720 2268.395 2914.100 2268.565 ;
        RECT 5.605 2267.305 6.815 2268.395 ;
        RECT 6.295 2266.765 6.815 2267.305 ;
        RECT 2912.805 2267.305 2914.015 2268.395 ;
        RECT 2912.805 2266.765 2913.325 2267.305 ;
        RECT 6.295 2264.215 6.815 2264.755 ;
        RECT 5.605 2263.125 6.815 2264.215 ;
        RECT 2906.365 2263.125 2906.655 2264.290 ;
        RECT 2912.805 2264.215 2913.325 2264.755 ;
        RECT 2909.315 2263.125 2909.645 2263.850 ;
        RECT 2912.805 2263.125 2914.015 2264.215 ;
        RECT 5.520 2262.955 6.900 2263.125 ;
        RECT 2906.300 2262.955 2906.740 2263.125 ;
        RECT 2909.040 2262.955 2910.420 2263.125 ;
        RECT 2912.720 2262.955 2914.100 2263.125 ;
        RECT 5.605 2261.865 6.815 2262.955 ;
        RECT 6.295 2261.325 6.815 2261.865 ;
        RECT 2912.805 2261.865 2914.015 2262.955 ;
        RECT 2912.805 2261.325 2913.325 2261.865 ;
        RECT 6.295 2258.775 6.815 2259.315 ;
        RECT 5.605 2257.685 6.815 2258.775 ;
        RECT 2906.365 2257.685 2906.655 2258.850 ;
        RECT 2912.805 2258.775 2913.325 2259.315 ;
        RECT 2912.805 2257.685 2914.015 2258.775 ;
        RECT 5.520 2257.515 6.900 2257.685 ;
        RECT 2906.300 2257.515 2906.740 2257.685 ;
        RECT 2912.720 2257.515 2914.100 2257.685 ;
        RECT 5.605 2256.425 6.815 2257.515 ;
        RECT 6.295 2255.885 6.815 2256.425 ;
        RECT 2912.805 2256.425 2914.015 2257.515 ;
        RECT 2912.805 2255.885 2913.325 2256.425 ;
        RECT 6.295 2253.335 6.815 2253.875 ;
        RECT 5.605 2252.245 6.815 2253.335 ;
        RECT 2906.365 2252.245 2906.655 2253.410 ;
        RECT 2912.805 2253.335 2913.325 2253.875 ;
        RECT 2912.805 2252.245 2914.015 2253.335 ;
        RECT 5.520 2252.075 6.900 2252.245 ;
        RECT 2906.300 2252.075 2906.740 2252.245 ;
        RECT 2912.720 2252.075 2914.100 2252.245 ;
        RECT 5.605 2250.985 6.815 2252.075 ;
        RECT 6.295 2250.445 6.815 2250.985 ;
        RECT 2912.805 2250.985 2914.015 2252.075 ;
        RECT 2912.805 2250.445 2913.325 2250.985 ;
        RECT 6.295 2247.895 6.815 2248.435 ;
        RECT 5.605 2246.805 6.815 2247.895 ;
        RECT 2906.365 2246.805 2906.655 2247.970 ;
        RECT 2912.805 2247.895 2913.325 2248.435 ;
        RECT 2912.805 2246.805 2914.015 2247.895 ;
        RECT 5.520 2246.635 6.900 2246.805 ;
        RECT 2906.300 2246.635 2906.740 2246.805 ;
        RECT 2912.720 2246.635 2914.100 2246.805 ;
        RECT 5.605 2245.545 6.815 2246.635 ;
        RECT 6.295 2245.005 6.815 2245.545 ;
        RECT 2912.805 2245.545 2914.015 2246.635 ;
        RECT 2912.805 2245.005 2913.325 2245.545 ;
        RECT 6.295 2242.455 6.815 2242.995 ;
        RECT 5.605 2241.365 6.815 2242.455 ;
        RECT 2906.365 2241.365 2906.655 2242.530 ;
        RECT 2912.805 2242.455 2913.325 2242.995 ;
        RECT 2912.805 2241.365 2914.015 2242.455 ;
        RECT 5.520 2241.195 6.900 2241.365 ;
        RECT 2906.300 2241.195 2906.740 2241.365 ;
        RECT 2912.720 2241.195 2914.100 2241.365 ;
        RECT 5.605 2240.105 6.815 2241.195 ;
        RECT 6.295 2239.565 6.815 2240.105 ;
        RECT 2912.805 2240.105 2914.015 2241.195 ;
        RECT 2912.805 2239.565 2913.325 2240.105 ;
        RECT 6.295 2237.015 6.815 2237.555 ;
        RECT 5.605 2235.925 6.815 2237.015 ;
        RECT 2906.365 2235.925 2906.655 2237.090 ;
        RECT 2912.805 2237.015 2913.325 2237.555 ;
        RECT 2912.805 2235.925 2914.015 2237.015 ;
        RECT 5.520 2235.755 6.900 2235.925 ;
        RECT 2906.300 2235.755 2906.740 2235.925 ;
        RECT 2912.720 2235.755 2914.100 2235.925 ;
        RECT 5.605 2234.665 6.815 2235.755 ;
        RECT 6.295 2234.125 6.815 2234.665 ;
        RECT 2912.805 2234.665 2914.015 2235.755 ;
        RECT 2912.805 2234.125 2913.325 2234.665 ;
        RECT 6.295 2231.575 6.815 2232.115 ;
        RECT 5.605 2230.485 6.815 2231.575 ;
        RECT 2906.365 2230.485 2906.655 2231.650 ;
        RECT 2912.805 2231.575 2913.325 2232.115 ;
        RECT 2912.805 2230.485 2914.015 2231.575 ;
        RECT 5.520 2230.315 6.900 2230.485 ;
        RECT 2906.300 2230.315 2906.740 2230.485 ;
        RECT 2912.720 2230.315 2914.100 2230.485 ;
        RECT 5.605 2229.225 6.815 2230.315 ;
        RECT 6.295 2228.685 6.815 2229.225 ;
        RECT 2912.805 2229.225 2914.015 2230.315 ;
        RECT 2912.805 2228.685 2913.325 2229.225 ;
        RECT 6.295 2226.135 6.815 2226.675 ;
        RECT 5.605 2225.045 6.815 2226.135 ;
        RECT 2906.365 2225.045 2906.655 2226.210 ;
        RECT 2912.805 2226.135 2913.325 2226.675 ;
        RECT 2912.805 2225.045 2914.015 2226.135 ;
        RECT 5.520 2224.875 6.900 2225.045 ;
        RECT 2906.300 2224.875 2906.740 2225.045 ;
        RECT 2912.720 2224.875 2914.100 2225.045 ;
        RECT 5.605 2223.785 6.815 2224.875 ;
        RECT 6.295 2223.245 6.815 2223.785 ;
        RECT 2912.805 2223.785 2914.015 2224.875 ;
        RECT 2912.805 2223.245 2913.325 2223.785 ;
        RECT 6.295 2220.695 6.815 2221.235 ;
        RECT 5.605 2219.605 6.815 2220.695 ;
        RECT 2906.365 2219.605 2906.655 2220.770 ;
        RECT 2912.805 2220.695 2913.325 2221.235 ;
        RECT 2912.805 2219.605 2914.015 2220.695 ;
        RECT 5.520 2219.435 6.900 2219.605 ;
        RECT 2906.300 2219.435 2906.740 2219.605 ;
        RECT 2912.720 2219.435 2914.100 2219.605 ;
        RECT 5.605 2218.345 6.815 2219.435 ;
        RECT 6.295 2217.805 6.815 2218.345 ;
        RECT 2912.805 2218.345 2914.015 2219.435 ;
        RECT 2912.805 2217.805 2913.325 2218.345 ;
        RECT 6.295 2215.255 6.815 2215.795 ;
        RECT 5.605 2214.165 6.815 2215.255 ;
        RECT 2906.365 2214.165 2906.655 2215.330 ;
        RECT 2912.805 2215.255 2913.325 2215.795 ;
        RECT 2912.805 2214.165 2914.015 2215.255 ;
        RECT 5.520 2213.995 6.900 2214.165 ;
        RECT 2906.300 2213.995 2906.740 2214.165 ;
        RECT 2912.720 2213.995 2914.100 2214.165 ;
        RECT 5.605 2212.905 6.815 2213.995 ;
        RECT 6.295 2212.365 6.815 2212.905 ;
        RECT 2912.805 2212.905 2914.015 2213.995 ;
        RECT 2912.805 2212.365 2913.325 2212.905 ;
        RECT 6.295 2209.815 6.815 2210.355 ;
        RECT 5.605 2208.725 6.815 2209.815 ;
        RECT 2906.365 2208.725 2906.655 2209.890 ;
        RECT 2912.805 2209.815 2913.325 2210.355 ;
        RECT 2912.805 2208.725 2914.015 2209.815 ;
        RECT 5.520 2208.555 6.900 2208.725 ;
        RECT 2906.300 2208.555 2906.740 2208.725 ;
        RECT 2912.720 2208.555 2914.100 2208.725 ;
        RECT 5.605 2207.465 6.815 2208.555 ;
        RECT 6.295 2206.925 6.815 2207.465 ;
        RECT 2912.805 2207.465 2914.015 2208.555 ;
        RECT 2912.805 2206.925 2913.325 2207.465 ;
        RECT 6.295 2204.375 6.815 2204.915 ;
        RECT 5.605 2203.285 6.815 2204.375 ;
        RECT 2906.365 2203.285 2906.655 2204.450 ;
        RECT 2912.805 2204.375 2913.325 2204.915 ;
        RECT 2912.805 2203.285 2914.015 2204.375 ;
        RECT 5.520 2203.115 6.900 2203.285 ;
        RECT 2906.300 2203.115 2906.740 2203.285 ;
        RECT 2912.720 2203.115 2914.100 2203.285 ;
        RECT 5.605 2202.025 6.815 2203.115 ;
        RECT 6.295 2201.485 6.815 2202.025 ;
        RECT 2912.805 2202.025 2914.015 2203.115 ;
        RECT 2912.805 2201.485 2913.325 2202.025 ;
        RECT 6.295 2198.935 6.815 2199.475 ;
        RECT 5.605 2197.845 6.815 2198.935 ;
        RECT 2906.365 2197.845 2906.655 2199.010 ;
        RECT 2912.805 2198.935 2913.325 2199.475 ;
        RECT 2912.805 2197.845 2914.015 2198.935 ;
        RECT 5.520 2197.675 6.900 2197.845 ;
        RECT 2906.300 2197.675 2906.740 2197.845 ;
        RECT 2912.720 2197.675 2914.100 2197.845 ;
        RECT 5.605 2196.585 6.815 2197.675 ;
        RECT 6.295 2196.045 6.815 2196.585 ;
        RECT 2912.805 2196.585 2914.015 2197.675 ;
        RECT 2912.805 2196.045 2913.325 2196.585 ;
        RECT 6.295 2193.495 6.815 2194.035 ;
        RECT 5.605 2192.405 6.815 2193.495 ;
        RECT 2906.365 2192.405 2906.655 2193.570 ;
        RECT 2912.805 2193.495 2913.325 2194.035 ;
        RECT 2912.805 2192.405 2914.015 2193.495 ;
        RECT 5.520 2192.235 6.900 2192.405 ;
        RECT 2906.300 2192.235 2906.740 2192.405 ;
        RECT 2912.720 2192.235 2914.100 2192.405 ;
        RECT 5.605 2191.145 6.815 2192.235 ;
        RECT 6.295 2190.605 6.815 2191.145 ;
        RECT 2912.805 2191.145 2914.015 2192.235 ;
        RECT 2912.805 2190.605 2913.325 2191.145 ;
        RECT 6.295 2188.055 6.815 2188.595 ;
        RECT 5.605 2186.965 6.815 2188.055 ;
        RECT 2906.365 2186.965 2906.655 2188.130 ;
        RECT 2912.805 2188.055 2913.325 2188.595 ;
        RECT 2912.805 2186.965 2914.015 2188.055 ;
        RECT 5.520 2186.795 6.900 2186.965 ;
        RECT 2906.300 2186.795 2906.740 2186.965 ;
        RECT 2912.720 2186.795 2914.100 2186.965 ;
        RECT 5.605 2185.705 6.815 2186.795 ;
        RECT 6.295 2185.165 6.815 2185.705 ;
        RECT 2912.805 2185.705 2914.015 2186.795 ;
        RECT 2912.805 2185.165 2913.325 2185.705 ;
        RECT 6.295 2182.615 6.815 2183.155 ;
        RECT 5.605 2181.525 6.815 2182.615 ;
        RECT 2906.365 2181.525 2906.655 2182.690 ;
        RECT 2912.805 2182.615 2913.325 2183.155 ;
        RECT 2912.805 2181.525 2914.015 2182.615 ;
        RECT 5.520 2181.355 6.900 2181.525 ;
        RECT 2906.300 2181.355 2906.740 2181.525 ;
        RECT 2912.720 2181.355 2914.100 2181.525 ;
        RECT 5.605 2180.265 6.815 2181.355 ;
        RECT 6.295 2179.725 6.815 2180.265 ;
        RECT 2912.805 2180.265 2914.015 2181.355 ;
        RECT 2912.805 2179.725 2913.325 2180.265 ;
        RECT 6.295 2177.175 6.815 2177.715 ;
        RECT 5.605 2176.085 6.815 2177.175 ;
        RECT 2906.365 2176.085 2906.655 2177.250 ;
        RECT 2912.805 2177.175 2913.325 2177.715 ;
        RECT 2912.805 2176.085 2914.015 2177.175 ;
        RECT 5.520 2175.915 6.900 2176.085 ;
        RECT 2906.300 2175.915 2906.740 2176.085 ;
        RECT 2912.720 2175.915 2914.100 2176.085 ;
        RECT 5.605 2174.825 6.815 2175.915 ;
        RECT 6.295 2174.285 6.815 2174.825 ;
        RECT 2912.805 2174.825 2914.015 2175.915 ;
        RECT 2912.805 2174.285 2913.325 2174.825 ;
        RECT 6.295 2171.735 6.815 2172.275 ;
        RECT 5.605 2170.645 6.815 2171.735 ;
        RECT 2906.365 2170.645 2906.655 2171.810 ;
        RECT 2912.805 2171.735 2913.325 2172.275 ;
        RECT 2912.805 2170.645 2914.015 2171.735 ;
        RECT 5.520 2170.475 6.900 2170.645 ;
        RECT 2906.300 2170.475 2906.740 2170.645 ;
        RECT 2912.720 2170.475 2914.100 2170.645 ;
        RECT 5.605 2169.385 6.815 2170.475 ;
        RECT 6.295 2168.845 6.815 2169.385 ;
        RECT 2912.805 2169.385 2914.015 2170.475 ;
        RECT 2912.805 2168.845 2913.325 2169.385 ;
        RECT 6.295 2166.295 6.815 2166.835 ;
        RECT 5.605 2165.205 6.815 2166.295 ;
        RECT 2906.365 2165.205 2906.655 2166.370 ;
        RECT 2912.805 2166.295 2913.325 2166.835 ;
        RECT 2912.805 2165.205 2914.015 2166.295 ;
        RECT 5.520 2165.035 6.900 2165.205 ;
        RECT 2906.300 2165.035 2906.740 2165.205 ;
        RECT 2912.720 2165.035 2914.100 2165.205 ;
        RECT 5.605 2163.945 6.815 2165.035 ;
        RECT 6.295 2163.405 6.815 2163.945 ;
        RECT 2912.805 2163.945 2914.015 2165.035 ;
        RECT 2912.805 2163.405 2913.325 2163.945 ;
        RECT 6.295 2160.855 6.815 2161.395 ;
        RECT 5.605 2159.765 6.815 2160.855 ;
        RECT 2906.365 2159.765 2906.655 2160.930 ;
        RECT 2912.805 2160.855 2913.325 2161.395 ;
        RECT 2912.805 2159.765 2914.015 2160.855 ;
        RECT 5.520 2159.595 6.900 2159.765 ;
        RECT 2906.300 2159.595 2906.740 2159.765 ;
        RECT 2912.720 2159.595 2914.100 2159.765 ;
        RECT 5.605 2158.505 6.815 2159.595 ;
        RECT 6.295 2157.965 6.815 2158.505 ;
        RECT 2912.805 2158.505 2914.015 2159.595 ;
        RECT 2912.805 2157.965 2913.325 2158.505 ;
        RECT 6.295 2155.415 6.815 2155.955 ;
        RECT 5.605 2154.325 6.815 2155.415 ;
        RECT 2906.365 2154.325 2906.655 2155.490 ;
        RECT 2912.805 2155.415 2913.325 2155.955 ;
        RECT 2912.805 2154.325 2914.015 2155.415 ;
        RECT 5.520 2154.155 6.900 2154.325 ;
        RECT 2906.300 2154.155 2906.740 2154.325 ;
        RECT 2912.720 2154.155 2914.100 2154.325 ;
        RECT 5.605 2153.065 6.815 2154.155 ;
        RECT 6.295 2152.525 6.815 2153.065 ;
        RECT 2912.805 2153.065 2914.015 2154.155 ;
        RECT 2912.805 2152.525 2913.325 2153.065 ;
        RECT 6.295 2149.975 6.815 2150.515 ;
        RECT 5.605 2148.885 6.815 2149.975 ;
        RECT 2906.365 2148.885 2906.655 2150.050 ;
        RECT 2912.805 2149.975 2913.325 2150.515 ;
        RECT 2912.805 2148.885 2914.015 2149.975 ;
        RECT 5.520 2148.715 6.900 2148.885 ;
        RECT 2906.300 2148.715 2906.740 2148.885 ;
        RECT 2912.720 2148.715 2914.100 2148.885 ;
        RECT 5.605 2147.625 6.815 2148.715 ;
        RECT 6.295 2147.085 6.815 2147.625 ;
        RECT 2912.805 2147.625 2914.015 2148.715 ;
        RECT 2912.805 2147.085 2913.325 2147.625 ;
        RECT 6.295 2144.535 6.815 2145.075 ;
        RECT 5.605 2143.445 6.815 2144.535 ;
        RECT 2906.365 2143.445 2906.655 2144.610 ;
        RECT 2912.805 2144.535 2913.325 2145.075 ;
        RECT 2912.805 2143.445 2914.015 2144.535 ;
        RECT 5.520 2143.275 6.900 2143.445 ;
        RECT 2906.300 2143.275 2906.740 2143.445 ;
        RECT 2912.720 2143.275 2914.100 2143.445 ;
        RECT 5.605 2142.185 6.815 2143.275 ;
        RECT 6.295 2141.645 6.815 2142.185 ;
        RECT 2912.805 2142.185 2914.015 2143.275 ;
        RECT 2912.805 2141.645 2913.325 2142.185 ;
        RECT 6.295 2139.095 6.815 2139.635 ;
        RECT 5.605 2138.005 6.815 2139.095 ;
        RECT 2906.365 2138.005 2906.655 2139.170 ;
        RECT 2912.805 2139.095 2913.325 2139.635 ;
        RECT 2912.805 2138.005 2914.015 2139.095 ;
        RECT 5.520 2137.835 6.900 2138.005 ;
        RECT 2906.300 2137.835 2906.740 2138.005 ;
        RECT 2912.720 2137.835 2914.100 2138.005 ;
        RECT 5.605 2136.745 6.815 2137.835 ;
        RECT 6.295 2136.205 6.815 2136.745 ;
        RECT 2912.805 2136.745 2914.015 2137.835 ;
        RECT 2912.805 2136.205 2913.325 2136.745 ;
        RECT 6.295 2133.655 6.815 2134.195 ;
        RECT 5.605 2132.565 6.815 2133.655 ;
        RECT 2906.365 2132.565 2906.655 2133.730 ;
        RECT 2912.805 2133.655 2913.325 2134.195 ;
        RECT 2912.805 2132.565 2914.015 2133.655 ;
        RECT 5.520 2132.395 6.900 2132.565 ;
        RECT 2906.300 2132.395 2906.740 2132.565 ;
        RECT 2912.720 2132.395 2914.100 2132.565 ;
        RECT 5.605 2131.305 6.815 2132.395 ;
        RECT 6.295 2130.765 6.815 2131.305 ;
        RECT 2912.805 2131.305 2914.015 2132.395 ;
        RECT 2912.805 2130.765 2913.325 2131.305 ;
        RECT 6.295 2128.215 6.815 2128.755 ;
        RECT 5.605 2127.125 6.815 2128.215 ;
        RECT 2906.365 2127.125 2906.655 2128.290 ;
        RECT 2912.805 2128.215 2913.325 2128.755 ;
        RECT 2912.805 2127.125 2914.015 2128.215 ;
        RECT 5.520 2126.955 6.900 2127.125 ;
        RECT 2906.300 2126.955 2906.740 2127.125 ;
        RECT 2912.720 2126.955 2914.100 2127.125 ;
        RECT 5.605 2125.865 6.815 2126.955 ;
        RECT 6.295 2125.325 6.815 2125.865 ;
        RECT 2912.805 2125.865 2914.015 2126.955 ;
        RECT 2912.805 2125.325 2913.325 2125.865 ;
        RECT 6.295 2122.775 6.815 2123.315 ;
        RECT 5.605 2121.685 6.815 2122.775 ;
        RECT 2906.365 2121.685 2906.655 2122.850 ;
        RECT 2912.805 2122.775 2913.325 2123.315 ;
        RECT 2912.805 2121.685 2914.015 2122.775 ;
        RECT 5.520 2121.515 6.900 2121.685 ;
        RECT 2906.300 2121.515 2906.740 2121.685 ;
        RECT 2912.720 2121.515 2914.100 2121.685 ;
        RECT 5.605 2120.425 6.815 2121.515 ;
        RECT 6.295 2119.885 6.815 2120.425 ;
        RECT 2912.805 2120.425 2914.015 2121.515 ;
        RECT 2912.805 2119.885 2913.325 2120.425 ;
        RECT 6.295 2117.335 6.815 2117.875 ;
        RECT 5.605 2116.245 6.815 2117.335 ;
        RECT 2906.365 2116.245 2906.655 2117.410 ;
        RECT 2912.805 2117.335 2913.325 2117.875 ;
        RECT 2909.315 2116.245 2909.645 2116.970 ;
        RECT 2912.805 2116.245 2914.015 2117.335 ;
        RECT 5.520 2116.075 6.900 2116.245 ;
        RECT 2906.300 2116.075 2906.740 2116.245 ;
        RECT 2909.040 2116.075 2910.420 2116.245 ;
        RECT 2912.720 2116.075 2914.100 2116.245 ;
        RECT 5.605 2114.985 6.815 2116.075 ;
        RECT 6.295 2114.445 6.815 2114.985 ;
        RECT 2912.805 2114.985 2914.015 2116.075 ;
        RECT 2912.805 2114.445 2913.325 2114.985 ;
        RECT 6.295 2111.895 6.815 2112.435 ;
        RECT 5.605 2110.805 6.815 2111.895 ;
        RECT 2906.365 2110.805 2906.655 2111.970 ;
        RECT 2912.805 2111.895 2913.325 2112.435 ;
        RECT 2912.805 2110.805 2914.015 2111.895 ;
        RECT 5.520 2110.635 6.900 2110.805 ;
        RECT 2906.300 2110.635 2906.740 2110.805 ;
        RECT 2912.720 2110.635 2914.100 2110.805 ;
        RECT 5.605 2109.545 6.815 2110.635 ;
        RECT 6.295 2109.005 6.815 2109.545 ;
        RECT 2912.805 2109.545 2914.015 2110.635 ;
        RECT 2912.805 2109.005 2913.325 2109.545 ;
        RECT 6.295 2106.455 6.815 2106.995 ;
        RECT 5.605 2105.365 6.815 2106.455 ;
        RECT 2906.365 2105.365 2906.655 2106.530 ;
        RECT 2912.805 2106.455 2913.325 2106.995 ;
        RECT 2912.805 2105.365 2914.015 2106.455 ;
        RECT 5.520 2105.195 6.900 2105.365 ;
        RECT 2906.300 2105.195 2906.740 2105.365 ;
        RECT 2912.720 2105.195 2914.100 2105.365 ;
        RECT 5.605 2104.105 6.815 2105.195 ;
        RECT 6.295 2103.565 6.815 2104.105 ;
        RECT 2912.805 2104.105 2914.015 2105.195 ;
        RECT 2912.805 2103.565 2913.325 2104.105 ;
        RECT 6.295 2101.015 6.815 2101.555 ;
        RECT 5.605 2099.925 6.815 2101.015 ;
        RECT 2906.365 2099.925 2906.655 2101.090 ;
        RECT 2912.805 2101.015 2913.325 2101.555 ;
        RECT 2912.805 2099.925 2914.015 2101.015 ;
        RECT 5.520 2099.755 6.900 2099.925 ;
        RECT 2906.300 2099.755 2906.740 2099.925 ;
        RECT 2912.720 2099.755 2914.100 2099.925 ;
        RECT 5.605 2098.665 6.815 2099.755 ;
        RECT 6.295 2098.125 6.815 2098.665 ;
        RECT 2912.805 2098.665 2914.015 2099.755 ;
        RECT 2912.805 2098.125 2913.325 2098.665 ;
        RECT 6.295 2095.575 6.815 2096.115 ;
        RECT 5.605 2094.485 6.815 2095.575 ;
        RECT 2906.365 2094.485 2906.655 2095.650 ;
        RECT 2912.805 2095.575 2913.325 2096.115 ;
        RECT 2912.805 2094.485 2914.015 2095.575 ;
        RECT 5.520 2094.315 6.900 2094.485 ;
        RECT 2906.300 2094.315 2906.740 2094.485 ;
        RECT 2912.720 2094.315 2914.100 2094.485 ;
        RECT 5.605 2093.225 6.815 2094.315 ;
        RECT 6.295 2092.685 6.815 2093.225 ;
        RECT 2912.805 2093.225 2914.015 2094.315 ;
        RECT 2912.805 2092.685 2913.325 2093.225 ;
        RECT 6.295 2090.135 6.815 2090.675 ;
        RECT 5.605 2089.045 6.815 2090.135 ;
        RECT 2906.365 2089.045 2906.655 2090.210 ;
        RECT 2912.805 2090.135 2913.325 2090.675 ;
        RECT 2912.805 2089.045 2914.015 2090.135 ;
        RECT 5.520 2088.875 6.900 2089.045 ;
        RECT 2906.300 2088.875 2906.740 2089.045 ;
        RECT 2912.720 2088.875 2914.100 2089.045 ;
        RECT 5.605 2087.785 6.815 2088.875 ;
        RECT 6.295 2087.245 6.815 2087.785 ;
        RECT 2912.805 2087.785 2914.015 2088.875 ;
        RECT 2912.805 2087.245 2913.325 2087.785 ;
        RECT 6.295 2084.695 6.815 2085.235 ;
        RECT 5.605 2083.605 6.815 2084.695 ;
        RECT 2906.365 2083.605 2906.655 2084.770 ;
        RECT 2912.805 2084.695 2913.325 2085.235 ;
        RECT 2912.805 2083.605 2914.015 2084.695 ;
        RECT 5.520 2083.435 6.900 2083.605 ;
        RECT 2906.300 2083.435 2906.740 2083.605 ;
        RECT 2912.720 2083.435 2914.100 2083.605 ;
        RECT 5.605 2082.345 6.815 2083.435 ;
        RECT 6.295 2081.805 6.815 2082.345 ;
        RECT 2912.805 2082.345 2914.015 2083.435 ;
        RECT 2912.805 2081.805 2913.325 2082.345 ;
        RECT 6.295 2079.255 6.815 2079.795 ;
        RECT 5.605 2078.165 6.815 2079.255 ;
        RECT 2906.365 2078.165 2906.655 2079.330 ;
        RECT 2912.805 2079.255 2913.325 2079.795 ;
        RECT 2912.805 2078.165 2914.015 2079.255 ;
        RECT 5.520 2077.995 6.900 2078.165 ;
        RECT 2906.300 2077.995 2906.740 2078.165 ;
        RECT 2912.720 2077.995 2914.100 2078.165 ;
        RECT 5.605 2076.905 6.815 2077.995 ;
        RECT 6.295 2076.365 6.815 2076.905 ;
        RECT 2912.805 2076.905 2914.015 2077.995 ;
        RECT 2912.805 2076.365 2913.325 2076.905 ;
        RECT 6.295 2073.815 6.815 2074.355 ;
        RECT 5.605 2072.725 6.815 2073.815 ;
        RECT 2906.365 2072.725 2906.655 2073.890 ;
        RECT 2912.805 2073.815 2913.325 2074.355 ;
        RECT 2912.805 2072.725 2914.015 2073.815 ;
        RECT 5.520 2072.555 6.900 2072.725 ;
        RECT 2906.300 2072.555 2906.740 2072.725 ;
        RECT 2912.720 2072.555 2914.100 2072.725 ;
        RECT 5.605 2071.465 6.815 2072.555 ;
        RECT 6.295 2070.925 6.815 2071.465 ;
        RECT 2912.805 2071.465 2914.015 2072.555 ;
        RECT 2912.805 2070.925 2913.325 2071.465 ;
        RECT 6.295 2068.375 6.815 2068.915 ;
        RECT 5.605 2067.285 6.815 2068.375 ;
        RECT 2906.365 2067.285 2906.655 2068.450 ;
        RECT 2912.805 2068.375 2913.325 2068.915 ;
        RECT 2912.805 2067.285 2914.015 2068.375 ;
        RECT 5.520 2067.115 6.900 2067.285 ;
        RECT 2906.300 2067.115 2906.740 2067.285 ;
        RECT 2912.720 2067.115 2914.100 2067.285 ;
        RECT 5.605 2066.025 6.815 2067.115 ;
        RECT 6.295 2065.485 6.815 2066.025 ;
        RECT 2912.805 2066.025 2914.015 2067.115 ;
        RECT 2912.805 2065.485 2913.325 2066.025 ;
        RECT 6.295 2062.935 6.815 2063.475 ;
        RECT 5.605 2061.845 6.815 2062.935 ;
        RECT 2906.365 2061.845 2906.655 2063.010 ;
        RECT 2912.805 2062.935 2913.325 2063.475 ;
        RECT 2912.805 2061.845 2914.015 2062.935 ;
        RECT 5.520 2061.675 6.900 2061.845 ;
        RECT 2906.300 2061.675 2906.740 2061.845 ;
        RECT 2912.720 2061.675 2914.100 2061.845 ;
        RECT 5.605 2060.585 6.815 2061.675 ;
        RECT 6.295 2060.045 6.815 2060.585 ;
        RECT 2912.805 2060.585 2914.015 2061.675 ;
        RECT 2912.805 2060.045 2913.325 2060.585 ;
        RECT 6.295 2057.495 6.815 2058.035 ;
        RECT 5.605 2056.405 6.815 2057.495 ;
        RECT 2906.365 2056.405 2906.655 2057.570 ;
        RECT 2912.805 2057.495 2913.325 2058.035 ;
        RECT 2912.805 2056.405 2914.015 2057.495 ;
        RECT 5.520 2056.235 6.900 2056.405 ;
        RECT 2906.300 2056.235 2906.740 2056.405 ;
        RECT 2912.720 2056.235 2914.100 2056.405 ;
        RECT 5.605 2055.145 6.815 2056.235 ;
        RECT 6.295 2054.605 6.815 2055.145 ;
        RECT 2912.805 2055.145 2914.015 2056.235 ;
        RECT 2912.805 2054.605 2913.325 2055.145 ;
        RECT 6.295 2052.055 6.815 2052.595 ;
        RECT 5.605 2050.965 6.815 2052.055 ;
        RECT 2906.365 2050.965 2906.655 2052.130 ;
        RECT 2912.805 2052.055 2913.325 2052.595 ;
        RECT 2912.805 2050.965 2914.015 2052.055 ;
        RECT 5.520 2050.795 6.900 2050.965 ;
        RECT 2906.300 2050.795 2906.740 2050.965 ;
        RECT 2912.720 2050.795 2914.100 2050.965 ;
        RECT 5.605 2049.705 6.815 2050.795 ;
        RECT 6.295 2049.165 6.815 2049.705 ;
        RECT 2912.805 2049.705 2914.015 2050.795 ;
        RECT 2912.805 2049.165 2913.325 2049.705 ;
        RECT 6.295 2046.615 6.815 2047.155 ;
        RECT 5.605 2045.525 6.815 2046.615 ;
        RECT 2906.365 2045.525 2906.655 2046.690 ;
        RECT 2912.805 2046.615 2913.325 2047.155 ;
        RECT 2912.805 2045.525 2914.015 2046.615 ;
        RECT 5.520 2045.355 6.900 2045.525 ;
        RECT 2906.300 2045.355 2906.740 2045.525 ;
        RECT 2912.720 2045.355 2914.100 2045.525 ;
        RECT 5.605 2044.265 6.815 2045.355 ;
        RECT 6.295 2043.725 6.815 2044.265 ;
        RECT 2912.805 2044.265 2914.015 2045.355 ;
        RECT 2912.805 2043.725 2913.325 2044.265 ;
        RECT 6.295 2041.175 6.815 2041.715 ;
        RECT 5.605 2040.085 6.815 2041.175 ;
        RECT 2906.365 2040.085 2906.655 2041.250 ;
        RECT 2912.805 2041.175 2913.325 2041.715 ;
        RECT 2912.805 2040.085 2914.015 2041.175 ;
        RECT 5.520 2039.915 6.900 2040.085 ;
        RECT 2906.300 2039.915 2906.740 2040.085 ;
        RECT 2912.720 2039.915 2914.100 2040.085 ;
        RECT 5.605 2038.825 6.815 2039.915 ;
        RECT 6.295 2038.285 6.815 2038.825 ;
        RECT 2912.805 2038.825 2914.015 2039.915 ;
        RECT 2912.805 2038.285 2913.325 2038.825 ;
        RECT 6.295 2035.735 6.815 2036.275 ;
        RECT 5.605 2034.645 6.815 2035.735 ;
        RECT 2906.365 2034.645 2906.655 2035.810 ;
        RECT 2912.805 2035.735 2913.325 2036.275 ;
        RECT 2912.805 2034.645 2914.015 2035.735 ;
        RECT 5.520 2034.475 6.900 2034.645 ;
        RECT 2906.300 2034.475 2906.740 2034.645 ;
        RECT 2912.720 2034.475 2914.100 2034.645 ;
        RECT 5.605 2033.385 6.815 2034.475 ;
        RECT 6.295 2032.845 6.815 2033.385 ;
        RECT 2912.805 2033.385 2914.015 2034.475 ;
        RECT 2912.805 2032.845 2913.325 2033.385 ;
        RECT 6.295 2030.295 6.815 2030.835 ;
        RECT 5.605 2029.205 6.815 2030.295 ;
        RECT 2906.365 2029.205 2906.655 2030.370 ;
        RECT 2912.805 2030.295 2913.325 2030.835 ;
        RECT 2912.805 2029.205 2914.015 2030.295 ;
        RECT 5.520 2029.035 6.900 2029.205 ;
        RECT 2906.300 2029.035 2906.740 2029.205 ;
        RECT 2912.720 2029.035 2914.100 2029.205 ;
        RECT 5.605 2027.945 6.815 2029.035 ;
        RECT 6.295 2027.405 6.815 2027.945 ;
        RECT 2912.805 2027.945 2914.015 2029.035 ;
        RECT 2912.805 2027.405 2913.325 2027.945 ;
        RECT 6.295 2024.855 6.815 2025.395 ;
        RECT 5.605 2023.765 6.815 2024.855 ;
        RECT 2906.365 2023.765 2906.655 2024.930 ;
        RECT 2912.805 2024.855 2913.325 2025.395 ;
        RECT 2912.805 2023.765 2914.015 2024.855 ;
        RECT 5.520 2023.595 6.900 2023.765 ;
        RECT 2906.300 2023.595 2906.740 2023.765 ;
        RECT 2912.720 2023.595 2914.100 2023.765 ;
        RECT 5.605 2022.505 6.815 2023.595 ;
        RECT 6.295 2021.965 6.815 2022.505 ;
        RECT 2912.805 2022.505 2914.015 2023.595 ;
        RECT 2912.805 2021.965 2913.325 2022.505 ;
        RECT 6.295 2019.415 6.815 2019.955 ;
        RECT 5.605 2018.325 6.815 2019.415 ;
        RECT 2906.365 2018.325 2906.655 2019.490 ;
        RECT 2912.805 2019.415 2913.325 2019.955 ;
        RECT 2912.805 2018.325 2914.015 2019.415 ;
        RECT 5.520 2018.155 6.900 2018.325 ;
        RECT 2906.300 2018.155 2906.740 2018.325 ;
        RECT 2912.720 2018.155 2914.100 2018.325 ;
        RECT 5.605 2017.065 6.815 2018.155 ;
        RECT 6.295 2016.525 6.815 2017.065 ;
        RECT 2912.805 2017.065 2914.015 2018.155 ;
        RECT 2912.805 2016.525 2913.325 2017.065 ;
        RECT 6.295 2013.975 6.815 2014.515 ;
        RECT 5.605 2012.885 6.815 2013.975 ;
        RECT 2906.365 2012.885 2906.655 2014.050 ;
        RECT 2912.805 2013.975 2913.325 2014.515 ;
        RECT 2912.805 2012.885 2914.015 2013.975 ;
        RECT 5.520 2012.715 6.900 2012.885 ;
        RECT 2906.300 2012.715 2906.740 2012.885 ;
        RECT 2912.720 2012.715 2914.100 2012.885 ;
        RECT 5.605 2011.625 6.815 2012.715 ;
        RECT 6.295 2011.085 6.815 2011.625 ;
        RECT 2912.805 2011.625 2914.015 2012.715 ;
        RECT 2912.805 2011.085 2913.325 2011.625 ;
        RECT 6.295 2008.535 6.815 2009.075 ;
        RECT 5.605 2007.445 6.815 2008.535 ;
        RECT 2906.365 2007.445 2906.655 2008.610 ;
        RECT 2912.805 2008.535 2913.325 2009.075 ;
        RECT 2912.805 2007.445 2914.015 2008.535 ;
        RECT 5.520 2007.275 6.900 2007.445 ;
        RECT 2906.300 2007.275 2906.740 2007.445 ;
        RECT 2912.720 2007.275 2914.100 2007.445 ;
        RECT 5.605 2006.185 6.815 2007.275 ;
        RECT 6.295 2005.645 6.815 2006.185 ;
        RECT 2912.805 2006.185 2914.015 2007.275 ;
        RECT 2912.805 2005.645 2913.325 2006.185 ;
        RECT 6.295 2003.095 6.815 2003.635 ;
        RECT 5.605 2002.005 6.815 2003.095 ;
        RECT 2906.365 2002.005 2906.655 2003.170 ;
        RECT 2912.805 2003.095 2913.325 2003.635 ;
        RECT 2912.805 2002.005 2914.015 2003.095 ;
        RECT 5.520 2001.835 6.900 2002.005 ;
        RECT 2906.300 2001.835 2906.740 2002.005 ;
        RECT 2912.720 2001.835 2914.100 2002.005 ;
        RECT 5.605 2000.745 6.815 2001.835 ;
        RECT 6.295 2000.205 6.815 2000.745 ;
        RECT 2912.805 2000.745 2914.015 2001.835 ;
        RECT 2912.805 2000.205 2913.325 2000.745 ;
        RECT 6.295 1997.655 6.815 1998.195 ;
        RECT 5.605 1996.565 6.815 1997.655 ;
        RECT 2906.365 1996.565 2906.655 1997.730 ;
        RECT 2912.805 1997.655 2913.325 1998.195 ;
        RECT 2912.805 1996.565 2914.015 1997.655 ;
        RECT 5.520 1996.395 6.900 1996.565 ;
        RECT 2906.300 1996.395 2906.740 1996.565 ;
        RECT 2912.720 1996.395 2914.100 1996.565 ;
        RECT 5.605 1995.305 6.815 1996.395 ;
        RECT 6.295 1994.765 6.815 1995.305 ;
        RECT 2912.805 1995.305 2914.015 1996.395 ;
        RECT 2912.805 1994.765 2913.325 1995.305 ;
        RECT 6.295 1992.215 6.815 1992.755 ;
        RECT 5.605 1991.125 6.815 1992.215 ;
        RECT 2906.365 1991.125 2906.655 1992.290 ;
        RECT 2912.805 1992.215 2913.325 1992.755 ;
        RECT 2912.805 1991.125 2914.015 1992.215 ;
        RECT 5.520 1990.955 6.900 1991.125 ;
        RECT 2906.300 1990.955 2906.740 1991.125 ;
        RECT 2912.720 1990.955 2914.100 1991.125 ;
        RECT 5.605 1989.865 6.815 1990.955 ;
        RECT 6.295 1989.325 6.815 1989.865 ;
        RECT 2912.805 1989.865 2914.015 1990.955 ;
        RECT 2912.805 1989.325 2913.325 1989.865 ;
        RECT 6.295 1986.775 6.815 1987.315 ;
        RECT 5.605 1985.685 6.815 1986.775 ;
        RECT 2906.365 1985.685 2906.655 1986.850 ;
        RECT 2912.805 1986.775 2913.325 1987.315 ;
        RECT 2912.805 1985.685 2914.015 1986.775 ;
        RECT 5.520 1985.515 6.900 1985.685 ;
        RECT 8.740 1985.515 10.120 1985.685 ;
        RECT 2906.300 1985.515 2906.740 1985.685 ;
        RECT 2912.720 1985.515 2914.100 1985.685 ;
        RECT 5.605 1984.425 6.815 1985.515 ;
        RECT 9.015 1984.790 9.345 1985.515 ;
        RECT 6.295 1983.885 6.815 1984.425 ;
        RECT 2912.805 1984.425 2914.015 1985.515 ;
        RECT 2912.805 1983.885 2913.325 1984.425 ;
        RECT 6.295 1981.335 6.815 1981.875 ;
        RECT 5.605 1980.245 6.815 1981.335 ;
        RECT 2906.365 1980.245 2906.655 1981.410 ;
        RECT 2912.805 1981.335 2913.325 1981.875 ;
        RECT 2912.805 1980.245 2914.015 1981.335 ;
        RECT 5.520 1980.075 6.900 1980.245 ;
        RECT 2906.300 1980.075 2906.740 1980.245 ;
        RECT 2912.720 1980.075 2914.100 1980.245 ;
        RECT 5.605 1978.985 6.815 1980.075 ;
        RECT 6.295 1978.445 6.815 1978.985 ;
        RECT 2912.805 1978.985 2914.015 1980.075 ;
        RECT 2912.805 1978.445 2913.325 1978.985 ;
        RECT 6.295 1975.895 6.815 1976.435 ;
        RECT 5.605 1974.805 6.815 1975.895 ;
        RECT 2906.365 1974.805 2906.655 1975.970 ;
        RECT 2912.805 1975.895 2913.325 1976.435 ;
        RECT 2912.805 1974.805 2914.015 1975.895 ;
        RECT 5.520 1974.635 6.900 1974.805 ;
        RECT 2906.300 1974.635 2906.740 1974.805 ;
        RECT 2912.720 1974.635 2914.100 1974.805 ;
        RECT 5.605 1973.545 6.815 1974.635 ;
        RECT 6.295 1973.005 6.815 1973.545 ;
        RECT 2912.805 1973.545 2914.015 1974.635 ;
        RECT 2912.805 1973.005 2913.325 1973.545 ;
        RECT 6.295 1970.455 6.815 1970.995 ;
        RECT 5.605 1969.365 6.815 1970.455 ;
        RECT 2906.365 1969.365 2906.655 1970.530 ;
        RECT 2912.805 1970.455 2913.325 1970.995 ;
        RECT 2912.805 1969.365 2914.015 1970.455 ;
        RECT 5.520 1969.195 6.900 1969.365 ;
        RECT 2906.300 1969.195 2906.740 1969.365 ;
        RECT 2912.720 1969.195 2914.100 1969.365 ;
        RECT 5.605 1968.105 6.815 1969.195 ;
        RECT 6.295 1967.565 6.815 1968.105 ;
        RECT 2912.805 1968.105 2914.015 1969.195 ;
        RECT 2912.805 1967.565 2913.325 1968.105 ;
        RECT 6.295 1965.015 6.815 1965.555 ;
        RECT 5.605 1963.925 6.815 1965.015 ;
        RECT 2906.365 1963.925 2906.655 1965.090 ;
        RECT 2912.805 1965.015 2913.325 1965.555 ;
        RECT 2912.805 1963.925 2914.015 1965.015 ;
        RECT 5.520 1963.755 6.900 1963.925 ;
        RECT 2906.300 1963.755 2906.740 1963.925 ;
        RECT 2912.720 1963.755 2914.100 1963.925 ;
        RECT 5.605 1962.665 6.815 1963.755 ;
        RECT 6.295 1962.125 6.815 1962.665 ;
        RECT 2912.805 1962.665 2914.015 1963.755 ;
        RECT 2912.805 1962.125 2913.325 1962.665 ;
        RECT 6.295 1959.575 6.815 1960.115 ;
        RECT 5.605 1958.485 6.815 1959.575 ;
        RECT 2906.365 1958.485 2906.655 1959.650 ;
        RECT 2912.805 1959.575 2913.325 1960.115 ;
        RECT 2912.805 1958.485 2914.015 1959.575 ;
        RECT 5.520 1958.315 6.900 1958.485 ;
        RECT 2906.300 1958.315 2906.740 1958.485 ;
        RECT 2912.720 1958.315 2914.100 1958.485 ;
        RECT 5.605 1957.225 6.815 1958.315 ;
        RECT 6.295 1956.685 6.815 1957.225 ;
        RECT 2912.805 1957.225 2914.015 1958.315 ;
        RECT 2912.805 1956.685 2913.325 1957.225 ;
        RECT 6.295 1954.135 6.815 1954.675 ;
        RECT 5.605 1953.045 6.815 1954.135 ;
        RECT 9.015 1953.045 9.345 1953.770 ;
        RECT 2906.365 1953.045 2906.655 1954.210 ;
        RECT 2912.805 1954.135 2913.325 1954.675 ;
        RECT 2912.805 1953.045 2914.015 1954.135 ;
        RECT 5.520 1952.875 6.900 1953.045 ;
        RECT 8.740 1952.875 10.120 1953.045 ;
        RECT 2906.300 1952.875 2906.740 1953.045 ;
        RECT 2912.720 1952.875 2914.100 1953.045 ;
        RECT 5.605 1951.785 6.815 1952.875 ;
        RECT 6.295 1951.245 6.815 1951.785 ;
        RECT 2912.805 1951.785 2914.015 1952.875 ;
        RECT 2912.805 1951.245 2913.325 1951.785 ;
        RECT 6.295 1948.695 6.815 1949.235 ;
        RECT 5.605 1947.605 6.815 1948.695 ;
        RECT 2906.365 1947.605 2906.655 1948.770 ;
        RECT 2912.805 1948.695 2913.325 1949.235 ;
        RECT 2912.805 1947.605 2914.015 1948.695 ;
        RECT 5.520 1947.435 6.900 1947.605 ;
        RECT 2906.300 1947.435 2906.740 1947.605 ;
        RECT 2912.720 1947.435 2914.100 1947.605 ;
        RECT 5.605 1946.345 6.815 1947.435 ;
        RECT 6.295 1945.805 6.815 1946.345 ;
        RECT 2912.805 1946.345 2914.015 1947.435 ;
        RECT 2912.805 1945.805 2913.325 1946.345 ;
        RECT 6.295 1943.255 6.815 1943.795 ;
        RECT 5.605 1942.165 6.815 1943.255 ;
        RECT 2906.365 1942.165 2906.655 1943.330 ;
        RECT 2912.805 1943.255 2913.325 1943.795 ;
        RECT 2912.805 1942.165 2914.015 1943.255 ;
        RECT 5.520 1941.995 6.900 1942.165 ;
        RECT 2906.300 1941.995 2906.740 1942.165 ;
        RECT 2912.720 1941.995 2914.100 1942.165 ;
        RECT 5.605 1940.905 6.815 1941.995 ;
        RECT 6.295 1940.365 6.815 1940.905 ;
        RECT 2912.805 1940.905 2914.015 1941.995 ;
        RECT 2912.805 1940.365 2913.325 1940.905 ;
        RECT 6.295 1937.815 6.815 1938.355 ;
        RECT 5.605 1936.725 6.815 1937.815 ;
        RECT 2906.365 1936.725 2906.655 1937.890 ;
        RECT 2912.805 1937.815 2913.325 1938.355 ;
        RECT 2912.805 1936.725 2914.015 1937.815 ;
        RECT 5.520 1936.555 6.900 1936.725 ;
        RECT 2906.300 1936.555 2906.740 1936.725 ;
        RECT 2909.040 1936.555 2910.420 1936.725 ;
        RECT 2912.720 1936.555 2914.100 1936.725 ;
        RECT 5.605 1935.465 6.815 1936.555 ;
        RECT 2909.315 1935.830 2909.645 1936.555 ;
        RECT 6.295 1934.925 6.815 1935.465 ;
        RECT 2912.805 1935.465 2914.015 1936.555 ;
        RECT 2912.805 1934.925 2913.325 1935.465 ;
        RECT 6.295 1932.375 6.815 1932.915 ;
        RECT 5.605 1931.285 6.815 1932.375 ;
        RECT 2906.365 1931.285 2906.655 1932.450 ;
        RECT 2912.805 1932.375 2913.325 1932.915 ;
        RECT 2912.805 1931.285 2914.015 1932.375 ;
        RECT 5.520 1931.115 6.900 1931.285 ;
        RECT 2906.300 1931.115 2906.740 1931.285 ;
        RECT 2912.720 1931.115 2914.100 1931.285 ;
        RECT 5.605 1930.025 6.815 1931.115 ;
        RECT 6.295 1929.485 6.815 1930.025 ;
        RECT 2912.805 1930.025 2914.015 1931.115 ;
        RECT 2912.805 1929.485 2913.325 1930.025 ;
        RECT 6.295 1926.935 6.815 1927.475 ;
        RECT 5.605 1925.845 6.815 1926.935 ;
        RECT 2906.365 1925.845 2906.655 1927.010 ;
        RECT 2912.805 1926.935 2913.325 1927.475 ;
        RECT 2912.805 1925.845 2914.015 1926.935 ;
        RECT 5.520 1925.675 6.900 1925.845 ;
        RECT 2906.300 1925.675 2906.740 1925.845 ;
        RECT 2912.720 1925.675 2914.100 1925.845 ;
        RECT 5.605 1924.585 6.815 1925.675 ;
        RECT 6.295 1924.045 6.815 1924.585 ;
        RECT 2912.805 1924.585 2914.015 1925.675 ;
        RECT 2912.805 1924.045 2913.325 1924.585 ;
        RECT 6.295 1921.495 6.815 1922.035 ;
        RECT 5.605 1920.405 6.815 1921.495 ;
        RECT 2906.365 1920.405 2906.655 1921.570 ;
        RECT 2912.805 1921.495 2913.325 1922.035 ;
        RECT 2912.805 1920.405 2914.015 1921.495 ;
        RECT 5.520 1920.235 6.900 1920.405 ;
        RECT 2906.300 1920.235 2906.740 1920.405 ;
        RECT 2912.720 1920.235 2914.100 1920.405 ;
        RECT 5.605 1919.145 6.815 1920.235 ;
        RECT 6.295 1918.605 6.815 1919.145 ;
        RECT 2912.805 1919.145 2914.015 1920.235 ;
        RECT 2912.805 1918.605 2913.325 1919.145 ;
        RECT 6.295 1916.055 6.815 1916.595 ;
        RECT 5.605 1914.965 6.815 1916.055 ;
        RECT 2906.365 1914.965 2906.655 1916.130 ;
        RECT 2912.805 1916.055 2913.325 1916.595 ;
        RECT 2912.805 1914.965 2914.015 1916.055 ;
        RECT 5.520 1914.795 6.900 1914.965 ;
        RECT 2906.300 1914.795 2906.740 1914.965 ;
        RECT 2912.720 1914.795 2914.100 1914.965 ;
        RECT 5.605 1913.705 6.815 1914.795 ;
        RECT 6.295 1913.165 6.815 1913.705 ;
        RECT 2912.805 1913.705 2914.015 1914.795 ;
        RECT 2912.805 1913.165 2913.325 1913.705 ;
        RECT 6.295 1910.615 6.815 1911.155 ;
        RECT 5.605 1909.525 6.815 1910.615 ;
        RECT 2906.365 1909.525 2906.655 1910.690 ;
        RECT 2912.805 1910.615 2913.325 1911.155 ;
        RECT 2912.805 1909.525 2914.015 1910.615 ;
        RECT 5.520 1909.355 6.900 1909.525 ;
        RECT 2906.300 1909.355 2906.740 1909.525 ;
        RECT 2912.720 1909.355 2914.100 1909.525 ;
        RECT 5.605 1908.265 6.815 1909.355 ;
        RECT 6.295 1907.725 6.815 1908.265 ;
        RECT 2912.805 1908.265 2914.015 1909.355 ;
        RECT 2912.805 1907.725 2913.325 1908.265 ;
        RECT 6.295 1905.175 6.815 1905.715 ;
        RECT 5.605 1904.085 6.815 1905.175 ;
        RECT 2906.365 1904.085 2906.655 1905.250 ;
        RECT 2912.805 1905.175 2913.325 1905.715 ;
        RECT 2912.805 1904.085 2914.015 1905.175 ;
        RECT 5.520 1903.915 6.900 1904.085 ;
        RECT 2906.300 1903.915 2906.740 1904.085 ;
        RECT 2912.720 1903.915 2914.100 1904.085 ;
        RECT 5.605 1902.825 6.815 1903.915 ;
        RECT 6.295 1902.285 6.815 1902.825 ;
        RECT 2912.805 1902.825 2914.015 1903.915 ;
        RECT 2912.805 1902.285 2913.325 1902.825 ;
        RECT 6.295 1899.735 6.815 1900.275 ;
        RECT 5.605 1898.645 6.815 1899.735 ;
        RECT 2906.365 1898.645 2906.655 1899.810 ;
        RECT 2912.805 1899.735 2913.325 1900.275 ;
        RECT 2912.805 1898.645 2914.015 1899.735 ;
        RECT 5.520 1898.475 6.900 1898.645 ;
        RECT 2906.300 1898.475 2906.740 1898.645 ;
        RECT 2912.720 1898.475 2914.100 1898.645 ;
        RECT 5.605 1897.385 6.815 1898.475 ;
        RECT 6.295 1896.845 6.815 1897.385 ;
        RECT 2912.805 1897.385 2914.015 1898.475 ;
        RECT 2912.805 1896.845 2913.325 1897.385 ;
        RECT 6.295 1894.295 6.815 1894.835 ;
        RECT 5.605 1893.205 6.815 1894.295 ;
        RECT 2906.365 1893.205 2906.655 1894.370 ;
        RECT 2912.805 1894.295 2913.325 1894.835 ;
        RECT 2912.805 1893.205 2914.015 1894.295 ;
        RECT 5.520 1893.035 6.900 1893.205 ;
        RECT 2906.300 1893.035 2906.740 1893.205 ;
        RECT 2912.720 1893.035 2914.100 1893.205 ;
        RECT 5.605 1891.945 6.815 1893.035 ;
        RECT 6.295 1891.405 6.815 1891.945 ;
        RECT 2912.805 1891.945 2914.015 1893.035 ;
        RECT 2912.805 1891.405 2913.325 1891.945 ;
        RECT 6.295 1888.855 6.815 1889.395 ;
        RECT 5.605 1887.765 6.815 1888.855 ;
        RECT 2906.365 1887.765 2906.655 1888.930 ;
        RECT 2912.805 1888.855 2913.325 1889.395 ;
        RECT 2912.805 1887.765 2914.015 1888.855 ;
        RECT 5.520 1887.595 6.900 1887.765 ;
        RECT 2906.300 1887.595 2906.740 1887.765 ;
        RECT 2912.720 1887.595 2914.100 1887.765 ;
        RECT 5.605 1886.505 6.815 1887.595 ;
        RECT 6.295 1885.965 6.815 1886.505 ;
        RECT 2912.805 1886.505 2914.015 1887.595 ;
        RECT 2912.805 1885.965 2913.325 1886.505 ;
        RECT 6.295 1883.415 6.815 1883.955 ;
        RECT 5.605 1882.325 6.815 1883.415 ;
        RECT 2906.365 1882.325 2906.655 1883.490 ;
        RECT 2912.805 1883.415 2913.325 1883.955 ;
        RECT 2912.805 1882.325 2914.015 1883.415 ;
        RECT 5.520 1882.155 6.900 1882.325 ;
        RECT 2906.300 1882.155 2906.740 1882.325 ;
        RECT 2912.720 1882.155 2914.100 1882.325 ;
        RECT 5.605 1881.065 6.815 1882.155 ;
        RECT 6.295 1880.525 6.815 1881.065 ;
        RECT 2912.805 1881.065 2914.015 1882.155 ;
        RECT 2912.805 1880.525 2913.325 1881.065 ;
        RECT 6.295 1877.975 6.815 1878.515 ;
        RECT 5.605 1876.885 6.815 1877.975 ;
        RECT 2906.365 1876.885 2906.655 1878.050 ;
        RECT 2912.805 1877.975 2913.325 1878.515 ;
        RECT 2912.805 1876.885 2914.015 1877.975 ;
        RECT 5.520 1876.715 6.900 1876.885 ;
        RECT 2906.300 1876.715 2906.740 1876.885 ;
        RECT 2912.720 1876.715 2914.100 1876.885 ;
        RECT 5.605 1875.625 6.815 1876.715 ;
        RECT 6.295 1875.085 6.815 1875.625 ;
        RECT 2912.805 1875.625 2914.015 1876.715 ;
        RECT 2912.805 1875.085 2913.325 1875.625 ;
        RECT 6.295 1872.535 6.815 1873.075 ;
        RECT 5.605 1871.445 6.815 1872.535 ;
        RECT 2906.365 1871.445 2906.655 1872.610 ;
        RECT 2912.805 1872.535 2913.325 1873.075 ;
        RECT 2912.805 1871.445 2914.015 1872.535 ;
        RECT 5.520 1871.275 6.900 1871.445 ;
        RECT 2906.300 1871.275 2906.740 1871.445 ;
        RECT 2912.720 1871.275 2914.100 1871.445 ;
        RECT 5.605 1870.185 6.815 1871.275 ;
        RECT 6.295 1869.645 6.815 1870.185 ;
        RECT 2912.805 1870.185 2914.015 1871.275 ;
        RECT 2912.805 1869.645 2913.325 1870.185 ;
        RECT 6.295 1867.095 6.815 1867.635 ;
        RECT 5.605 1866.005 6.815 1867.095 ;
        RECT 2906.365 1866.005 2906.655 1867.170 ;
        RECT 2912.805 1867.095 2913.325 1867.635 ;
        RECT 2912.805 1866.005 2914.015 1867.095 ;
        RECT 5.520 1865.835 6.900 1866.005 ;
        RECT 2906.300 1865.835 2906.740 1866.005 ;
        RECT 2912.720 1865.835 2914.100 1866.005 ;
        RECT 5.605 1864.745 6.815 1865.835 ;
        RECT 6.295 1864.205 6.815 1864.745 ;
        RECT 2912.805 1864.745 2914.015 1865.835 ;
        RECT 2912.805 1864.205 2913.325 1864.745 ;
        RECT 6.295 1861.655 6.815 1862.195 ;
        RECT 5.605 1860.565 6.815 1861.655 ;
        RECT 2906.365 1860.565 2906.655 1861.730 ;
        RECT 2912.805 1861.655 2913.325 1862.195 ;
        RECT 2912.805 1860.565 2914.015 1861.655 ;
        RECT 5.520 1860.395 6.900 1860.565 ;
        RECT 2906.300 1860.395 2906.740 1860.565 ;
        RECT 2912.720 1860.395 2914.100 1860.565 ;
        RECT 5.605 1859.305 6.815 1860.395 ;
        RECT 6.295 1858.765 6.815 1859.305 ;
        RECT 2912.805 1859.305 2914.015 1860.395 ;
        RECT 2912.805 1858.765 2913.325 1859.305 ;
        RECT 6.295 1856.215 6.815 1856.755 ;
        RECT 5.605 1855.125 6.815 1856.215 ;
        RECT 2906.365 1855.125 2906.655 1856.290 ;
        RECT 2912.805 1856.215 2913.325 1856.755 ;
        RECT 2912.805 1855.125 2914.015 1856.215 ;
        RECT 5.520 1854.955 6.900 1855.125 ;
        RECT 2906.300 1854.955 2906.740 1855.125 ;
        RECT 2912.720 1854.955 2914.100 1855.125 ;
        RECT 5.605 1853.865 6.815 1854.955 ;
        RECT 6.295 1853.325 6.815 1853.865 ;
        RECT 2912.805 1853.865 2914.015 1854.955 ;
        RECT 2912.805 1853.325 2913.325 1853.865 ;
        RECT 6.295 1850.775 6.815 1851.315 ;
        RECT 5.605 1849.685 6.815 1850.775 ;
        RECT 2906.365 1849.685 2906.655 1850.850 ;
        RECT 2912.805 1850.775 2913.325 1851.315 ;
        RECT 2912.805 1849.685 2914.015 1850.775 ;
        RECT 5.520 1849.515 6.900 1849.685 ;
        RECT 2906.300 1849.515 2906.740 1849.685 ;
        RECT 2912.720 1849.515 2914.100 1849.685 ;
        RECT 5.605 1848.425 6.815 1849.515 ;
        RECT 6.295 1847.885 6.815 1848.425 ;
        RECT 2912.805 1848.425 2914.015 1849.515 ;
        RECT 2912.805 1847.885 2913.325 1848.425 ;
        RECT 6.295 1845.335 6.815 1845.875 ;
        RECT 5.605 1844.245 6.815 1845.335 ;
        RECT 2906.365 1844.245 2906.655 1845.410 ;
        RECT 2912.805 1845.335 2913.325 1845.875 ;
        RECT 2912.805 1844.245 2914.015 1845.335 ;
        RECT 5.520 1844.075 6.900 1844.245 ;
        RECT 2906.300 1844.075 2906.740 1844.245 ;
        RECT 2912.720 1844.075 2914.100 1844.245 ;
        RECT 5.605 1842.985 6.815 1844.075 ;
        RECT 6.295 1842.445 6.815 1842.985 ;
        RECT 2912.805 1842.985 2914.015 1844.075 ;
        RECT 2912.805 1842.445 2913.325 1842.985 ;
        RECT 6.295 1839.895 6.815 1840.435 ;
        RECT 5.605 1838.805 6.815 1839.895 ;
        RECT 2906.365 1838.805 2906.655 1839.970 ;
        RECT 2912.805 1839.895 2913.325 1840.435 ;
        RECT 2912.805 1838.805 2914.015 1839.895 ;
        RECT 5.520 1838.635 6.900 1838.805 ;
        RECT 2906.300 1838.635 2906.740 1838.805 ;
        RECT 2912.720 1838.635 2914.100 1838.805 ;
        RECT 5.605 1837.545 6.815 1838.635 ;
        RECT 6.295 1837.005 6.815 1837.545 ;
        RECT 2912.805 1837.545 2914.015 1838.635 ;
        RECT 2912.805 1837.005 2913.325 1837.545 ;
        RECT 6.295 1834.455 6.815 1834.995 ;
        RECT 5.605 1833.365 6.815 1834.455 ;
        RECT 2906.365 1833.365 2906.655 1834.530 ;
        RECT 2912.805 1834.455 2913.325 1834.995 ;
        RECT 2912.805 1833.365 2914.015 1834.455 ;
        RECT 5.520 1833.195 6.900 1833.365 ;
        RECT 2906.300 1833.195 2906.740 1833.365 ;
        RECT 2912.720 1833.195 2914.100 1833.365 ;
        RECT 5.605 1832.105 6.815 1833.195 ;
        RECT 6.295 1831.565 6.815 1832.105 ;
        RECT 2912.805 1832.105 2914.015 1833.195 ;
        RECT 2912.805 1831.565 2913.325 1832.105 ;
        RECT 6.295 1829.015 6.815 1829.555 ;
        RECT 5.605 1827.925 6.815 1829.015 ;
        RECT 2906.365 1827.925 2906.655 1829.090 ;
        RECT 2912.805 1829.015 2913.325 1829.555 ;
        RECT 2912.805 1827.925 2914.015 1829.015 ;
        RECT 5.520 1827.755 6.900 1827.925 ;
        RECT 2906.300 1827.755 2906.740 1827.925 ;
        RECT 2912.720 1827.755 2914.100 1827.925 ;
        RECT 5.605 1826.665 6.815 1827.755 ;
        RECT 6.295 1826.125 6.815 1826.665 ;
        RECT 2912.805 1826.665 2914.015 1827.755 ;
        RECT 2912.805 1826.125 2913.325 1826.665 ;
        RECT 6.295 1823.575 6.815 1824.115 ;
        RECT 5.605 1822.485 6.815 1823.575 ;
        RECT 2906.365 1822.485 2906.655 1823.650 ;
        RECT 2912.805 1823.575 2913.325 1824.115 ;
        RECT 2912.805 1822.485 2914.015 1823.575 ;
        RECT 5.520 1822.315 6.900 1822.485 ;
        RECT 2906.300 1822.315 2906.740 1822.485 ;
        RECT 2912.720 1822.315 2914.100 1822.485 ;
        RECT 5.605 1821.225 6.815 1822.315 ;
        RECT 6.295 1820.685 6.815 1821.225 ;
        RECT 2912.805 1821.225 2914.015 1822.315 ;
        RECT 2912.805 1820.685 2913.325 1821.225 ;
        RECT 6.295 1818.135 6.815 1818.675 ;
        RECT 5.605 1817.045 6.815 1818.135 ;
        RECT 2906.365 1817.045 2906.655 1818.210 ;
        RECT 2912.805 1818.135 2913.325 1818.675 ;
        RECT 2912.805 1817.045 2914.015 1818.135 ;
        RECT 5.520 1816.875 6.900 1817.045 ;
        RECT 2906.300 1816.875 2906.740 1817.045 ;
        RECT 2912.720 1816.875 2914.100 1817.045 ;
        RECT 5.605 1815.785 6.815 1816.875 ;
        RECT 6.295 1815.245 6.815 1815.785 ;
        RECT 2912.805 1815.785 2914.015 1816.875 ;
        RECT 2912.805 1815.245 2913.325 1815.785 ;
        RECT 6.295 1812.695 6.815 1813.235 ;
        RECT 5.605 1811.605 6.815 1812.695 ;
        RECT 2906.365 1811.605 2906.655 1812.770 ;
        RECT 2912.805 1812.695 2913.325 1813.235 ;
        RECT 2912.805 1811.605 2914.015 1812.695 ;
        RECT 5.520 1811.435 6.900 1811.605 ;
        RECT 2906.300 1811.435 2906.740 1811.605 ;
        RECT 2912.720 1811.435 2914.100 1811.605 ;
        RECT 5.605 1810.345 6.815 1811.435 ;
        RECT 6.295 1809.805 6.815 1810.345 ;
        RECT 2912.805 1810.345 2914.015 1811.435 ;
        RECT 2912.805 1809.805 2913.325 1810.345 ;
        RECT 6.295 1807.255 6.815 1807.795 ;
        RECT 5.605 1806.165 6.815 1807.255 ;
        RECT 2906.365 1806.165 2906.655 1807.330 ;
        RECT 2912.805 1807.255 2913.325 1807.795 ;
        RECT 2912.805 1806.165 2914.015 1807.255 ;
        RECT 5.520 1805.995 6.900 1806.165 ;
        RECT 2906.300 1805.995 2906.740 1806.165 ;
        RECT 2912.720 1805.995 2914.100 1806.165 ;
        RECT 5.605 1804.905 6.815 1805.995 ;
        RECT 6.295 1804.365 6.815 1804.905 ;
        RECT 2912.805 1804.905 2914.015 1805.995 ;
        RECT 2912.805 1804.365 2913.325 1804.905 ;
        RECT 6.295 1801.815 6.815 1802.355 ;
        RECT 5.605 1800.725 6.815 1801.815 ;
        RECT 2906.365 1800.725 2906.655 1801.890 ;
        RECT 2912.805 1801.815 2913.325 1802.355 ;
        RECT 2912.805 1800.725 2914.015 1801.815 ;
        RECT 5.520 1800.555 6.900 1800.725 ;
        RECT 2906.300 1800.555 2906.740 1800.725 ;
        RECT 2912.720 1800.555 2914.100 1800.725 ;
        RECT 5.605 1799.465 6.815 1800.555 ;
        RECT 6.295 1798.925 6.815 1799.465 ;
        RECT 2912.805 1799.465 2914.015 1800.555 ;
        RECT 2912.805 1798.925 2913.325 1799.465 ;
        RECT 6.295 1796.375 6.815 1796.915 ;
        RECT 5.605 1795.285 6.815 1796.375 ;
        RECT 2906.365 1795.285 2906.655 1796.450 ;
        RECT 2912.805 1796.375 2913.325 1796.915 ;
        RECT 2912.805 1795.285 2914.015 1796.375 ;
        RECT 5.520 1795.115 6.900 1795.285 ;
        RECT 2906.300 1795.115 2906.740 1795.285 ;
        RECT 2912.720 1795.115 2914.100 1795.285 ;
        RECT 5.605 1794.025 6.815 1795.115 ;
        RECT 6.295 1793.485 6.815 1794.025 ;
        RECT 2912.805 1794.025 2914.015 1795.115 ;
        RECT 2912.805 1793.485 2913.325 1794.025 ;
        RECT 6.295 1790.935 6.815 1791.475 ;
        RECT 5.605 1789.845 6.815 1790.935 ;
        RECT 2906.365 1789.845 2906.655 1791.010 ;
        RECT 2912.805 1790.935 2913.325 1791.475 ;
        RECT 2912.805 1789.845 2914.015 1790.935 ;
        RECT 5.520 1789.675 6.900 1789.845 ;
        RECT 2906.300 1789.675 2906.740 1789.845 ;
        RECT 2912.720 1789.675 2914.100 1789.845 ;
        RECT 5.605 1788.585 6.815 1789.675 ;
        RECT 6.295 1788.045 6.815 1788.585 ;
        RECT 2912.805 1788.585 2914.015 1789.675 ;
        RECT 2912.805 1788.045 2913.325 1788.585 ;
        RECT 6.295 1785.495 6.815 1786.035 ;
        RECT 5.605 1784.405 6.815 1785.495 ;
        RECT 2906.365 1784.405 2906.655 1785.570 ;
        RECT 2912.805 1785.495 2913.325 1786.035 ;
        RECT 2912.805 1784.405 2914.015 1785.495 ;
        RECT 5.520 1784.235 6.900 1784.405 ;
        RECT 2906.300 1784.235 2906.740 1784.405 ;
        RECT 2912.720 1784.235 2914.100 1784.405 ;
        RECT 5.605 1783.145 6.815 1784.235 ;
        RECT 6.295 1782.605 6.815 1783.145 ;
        RECT 2912.805 1783.145 2914.015 1784.235 ;
        RECT 2912.805 1782.605 2913.325 1783.145 ;
        RECT 6.295 1780.055 6.815 1780.595 ;
        RECT 5.605 1778.965 6.815 1780.055 ;
        RECT 2906.365 1778.965 2906.655 1780.130 ;
        RECT 2912.805 1780.055 2913.325 1780.595 ;
        RECT 2912.805 1778.965 2914.015 1780.055 ;
        RECT 5.520 1778.795 6.900 1778.965 ;
        RECT 8.740 1778.795 10.120 1778.965 ;
        RECT 2906.300 1778.795 2906.740 1778.965 ;
        RECT 2912.720 1778.795 2914.100 1778.965 ;
        RECT 5.605 1777.705 6.815 1778.795 ;
        RECT 9.015 1778.070 9.345 1778.795 ;
        RECT 6.295 1777.165 6.815 1777.705 ;
        RECT 2912.805 1777.705 2914.015 1778.795 ;
        RECT 2912.805 1777.165 2913.325 1777.705 ;
        RECT 6.295 1774.615 6.815 1775.155 ;
        RECT 5.605 1773.525 6.815 1774.615 ;
        RECT 2906.365 1773.525 2906.655 1774.690 ;
        RECT 2912.805 1774.615 2913.325 1775.155 ;
        RECT 2912.805 1773.525 2914.015 1774.615 ;
        RECT 5.520 1773.355 6.900 1773.525 ;
        RECT 2906.300 1773.355 2906.740 1773.525 ;
        RECT 2912.720 1773.355 2914.100 1773.525 ;
        RECT 5.605 1772.265 6.815 1773.355 ;
        RECT 6.295 1771.725 6.815 1772.265 ;
        RECT 2912.805 1772.265 2914.015 1773.355 ;
        RECT 2912.805 1771.725 2913.325 1772.265 ;
        RECT 6.295 1769.175 6.815 1769.715 ;
        RECT 5.605 1768.085 6.815 1769.175 ;
        RECT 2906.365 1768.085 2906.655 1769.250 ;
        RECT 2912.805 1769.175 2913.325 1769.715 ;
        RECT 2912.805 1768.085 2914.015 1769.175 ;
        RECT 5.520 1767.915 6.900 1768.085 ;
        RECT 2906.300 1767.915 2906.740 1768.085 ;
        RECT 2912.720 1767.915 2914.100 1768.085 ;
        RECT 5.605 1766.825 6.815 1767.915 ;
        RECT 6.295 1766.285 6.815 1766.825 ;
        RECT 2912.805 1766.825 2914.015 1767.915 ;
        RECT 2912.805 1766.285 2913.325 1766.825 ;
        RECT 6.295 1763.735 6.815 1764.275 ;
        RECT 5.605 1762.645 6.815 1763.735 ;
        RECT 2906.365 1762.645 2906.655 1763.810 ;
        RECT 2912.805 1763.735 2913.325 1764.275 ;
        RECT 2912.805 1762.645 2914.015 1763.735 ;
        RECT 5.520 1762.475 6.900 1762.645 ;
        RECT 2906.300 1762.475 2906.740 1762.645 ;
        RECT 2912.720 1762.475 2914.100 1762.645 ;
        RECT 5.605 1761.385 6.815 1762.475 ;
        RECT 6.295 1760.845 6.815 1761.385 ;
        RECT 2912.805 1761.385 2914.015 1762.475 ;
        RECT 2912.805 1760.845 2913.325 1761.385 ;
        RECT 6.295 1758.295 6.815 1758.835 ;
        RECT 5.605 1757.205 6.815 1758.295 ;
        RECT 2906.365 1757.205 2906.655 1758.370 ;
        RECT 2912.805 1758.295 2913.325 1758.835 ;
        RECT 2912.805 1757.205 2914.015 1758.295 ;
        RECT 5.520 1757.035 6.900 1757.205 ;
        RECT 2906.300 1757.035 2906.740 1757.205 ;
        RECT 2912.720 1757.035 2914.100 1757.205 ;
        RECT 5.605 1755.945 6.815 1757.035 ;
        RECT 6.295 1755.405 6.815 1755.945 ;
        RECT 2912.805 1755.945 2914.015 1757.035 ;
        RECT 2912.805 1755.405 2913.325 1755.945 ;
        RECT 6.295 1752.855 6.815 1753.395 ;
        RECT 5.605 1751.765 6.815 1752.855 ;
        RECT 2906.365 1751.765 2906.655 1752.930 ;
        RECT 2912.805 1752.855 2913.325 1753.395 ;
        RECT 2912.805 1751.765 2914.015 1752.855 ;
        RECT 5.520 1751.595 6.900 1751.765 ;
        RECT 2906.300 1751.595 2906.740 1751.765 ;
        RECT 2912.720 1751.595 2914.100 1751.765 ;
        RECT 5.605 1750.505 6.815 1751.595 ;
        RECT 6.295 1749.965 6.815 1750.505 ;
        RECT 2912.805 1750.505 2914.015 1751.595 ;
        RECT 2912.805 1749.965 2913.325 1750.505 ;
        RECT 6.295 1747.415 6.815 1747.955 ;
        RECT 5.605 1746.325 6.815 1747.415 ;
        RECT 2906.365 1746.325 2906.655 1747.490 ;
        RECT 2912.805 1747.415 2913.325 1747.955 ;
        RECT 2912.805 1746.325 2914.015 1747.415 ;
        RECT 5.520 1746.155 6.900 1746.325 ;
        RECT 2906.300 1746.155 2906.740 1746.325 ;
        RECT 2912.720 1746.155 2914.100 1746.325 ;
        RECT 5.605 1745.065 6.815 1746.155 ;
        RECT 6.295 1744.525 6.815 1745.065 ;
        RECT 2912.805 1745.065 2914.015 1746.155 ;
        RECT 2912.805 1744.525 2913.325 1745.065 ;
        RECT 6.295 1741.975 6.815 1742.515 ;
        RECT 5.605 1740.885 6.815 1741.975 ;
        RECT 2906.365 1740.885 2906.655 1742.050 ;
        RECT 2912.805 1741.975 2913.325 1742.515 ;
        RECT 2912.805 1740.885 2914.015 1741.975 ;
        RECT 5.520 1740.715 6.900 1740.885 ;
        RECT 2906.300 1740.715 2906.740 1740.885 ;
        RECT 2912.720 1740.715 2914.100 1740.885 ;
        RECT 5.605 1739.625 6.815 1740.715 ;
        RECT 6.295 1739.085 6.815 1739.625 ;
        RECT 2912.805 1739.625 2914.015 1740.715 ;
        RECT 2912.805 1739.085 2913.325 1739.625 ;
        RECT 6.295 1736.535 6.815 1737.075 ;
        RECT 5.605 1735.445 6.815 1736.535 ;
        RECT 2906.365 1735.445 2906.655 1736.610 ;
        RECT 2912.805 1736.535 2913.325 1737.075 ;
        RECT 2912.805 1735.445 2914.015 1736.535 ;
        RECT 5.520 1735.275 6.900 1735.445 ;
        RECT 2906.300 1735.275 2906.740 1735.445 ;
        RECT 2912.720 1735.275 2914.100 1735.445 ;
        RECT 5.605 1734.185 6.815 1735.275 ;
        RECT 6.295 1733.645 6.815 1734.185 ;
        RECT 2912.805 1734.185 2914.015 1735.275 ;
        RECT 2912.805 1733.645 2913.325 1734.185 ;
        RECT 6.295 1731.095 6.815 1731.635 ;
        RECT 5.605 1730.005 6.815 1731.095 ;
        RECT 2906.365 1730.005 2906.655 1731.170 ;
        RECT 2912.805 1731.095 2913.325 1731.635 ;
        RECT 2912.805 1730.005 2914.015 1731.095 ;
        RECT 5.520 1729.835 6.900 1730.005 ;
        RECT 2906.300 1729.835 2906.740 1730.005 ;
        RECT 2912.720 1729.835 2914.100 1730.005 ;
        RECT 5.605 1728.745 6.815 1729.835 ;
        RECT 6.295 1728.205 6.815 1728.745 ;
        RECT 2912.805 1728.745 2914.015 1729.835 ;
        RECT 2912.805 1728.205 2913.325 1728.745 ;
        RECT 6.295 1725.655 6.815 1726.195 ;
        RECT 5.605 1724.565 6.815 1725.655 ;
        RECT 2906.365 1724.565 2906.655 1725.730 ;
        RECT 2912.805 1725.655 2913.325 1726.195 ;
        RECT 2912.805 1724.565 2914.015 1725.655 ;
        RECT 5.520 1724.395 6.900 1724.565 ;
        RECT 2906.300 1724.395 2906.740 1724.565 ;
        RECT 2912.720 1724.395 2914.100 1724.565 ;
        RECT 5.605 1723.305 6.815 1724.395 ;
        RECT 6.295 1722.765 6.815 1723.305 ;
        RECT 2912.805 1723.305 2914.015 1724.395 ;
        RECT 2912.805 1722.765 2913.325 1723.305 ;
        RECT 6.295 1720.215 6.815 1720.755 ;
        RECT 5.605 1719.125 6.815 1720.215 ;
        RECT 2906.365 1719.125 2906.655 1720.290 ;
        RECT 2912.805 1720.215 2913.325 1720.755 ;
        RECT 2912.805 1719.125 2914.015 1720.215 ;
        RECT 5.520 1718.955 6.900 1719.125 ;
        RECT 2906.300 1718.955 2906.740 1719.125 ;
        RECT 2912.720 1718.955 2914.100 1719.125 ;
        RECT 5.605 1717.865 6.815 1718.955 ;
        RECT 6.295 1717.325 6.815 1717.865 ;
        RECT 2912.805 1717.865 2914.015 1718.955 ;
        RECT 2912.805 1717.325 2913.325 1717.865 ;
        RECT 6.295 1714.775 6.815 1715.315 ;
        RECT 5.605 1713.685 6.815 1714.775 ;
        RECT 2906.365 1713.685 2906.655 1714.850 ;
        RECT 2912.805 1714.775 2913.325 1715.315 ;
        RECT 2912.805 1713.685 2914.015 1714.775 ;
        RECT 5.520 1713.515 6.900 1713.685 ;
        RECT 2906.300 1713.515 2906.740 1713.685 ;
        RECT 2912.720 1713.515 2914.100 1713.685 ;
        RECT 5.605 1712.425 6.815 1713.515 ;
        RECT 6.295 1711.885 6.815 1712.425 ;
        RECT 2912.805 1712.425 2914.015 1713.515 ;
        RECT 2912.805 1711.885 2913.325 1712.425 ;
        RECT 6.295 1709.335 6.815 1709.875 ;
        RECT 5.605 1708.245 6.815 1709.335 ;
        RECT 2906.365 1708.245 2906.655 1709.410 ;
        RECT 2912.805 1709.335 2913.325 1709.875 ;
        RECT 2912.805 1708.245 2914.015 1709.335 ;
        RECT 5.520 1708.075 6.900 1708.245 ;
        RECT 8.740 1708.075 10.120 1708.245 ;
        RECT 2906.300 1708.075 2906.740 1708.245 ;
        RECT 2912.720 1708.075 2914.100 1708.245 ;
        RECT 5.605 1706.985 6.815 1708.075 ;
        RECT 9.015 1707.350 9.345 1708.075 ;
        RECT 6.295 1706.445 6.815 1706.985 ;
        RECT 2912.805 1706.985 2914.015 1708.075 ;
        RECT 2912.805 1706.445 2913.325 1706.985 ;
        RECT 6.295 1703.895 6.815 1704.435 ;
        RECT 5.605 1702.805 6.815 1703.895 ;
        RECT 2906.365 1702.805 2906.655 1703.970 ;
        RECT 2912.805 1703.895 2913.325 1704.435 ;
        RECT 2912.805 1702.805 2914.015 1703.895 ;
        RECT 5.520 1702.635 6.900 1702.805 ;
        RECT 2906.300 1702.635 2906.740 1702.805 ;
        RECT 2912.720 1702.635 2914.100 1702.805 ;
        RECT 5.605 1701.545 6.815 1702.635 ;
        RECT 6.295 1701.005 6.815 1701.545 ;
        RECT 2912.805 1701.545 2914.015 1702.635 ;
        RECT 2912.805 1701.005 2913.325 1701.545 ;
        RECT 6.295 1698.455 6.815 1698.995 ;
        RECT 5.605 1697.365 6.815 1698.455 ;
        RECT 2906.365 1697.365 2906.655 1698.530 ;
        RECT 2912.805 1698.455 2913.325 1698.995 ;
        RECT 2912.805 1697.365 2914.015 1698.455 ;
        RECT 5.520 1697.195 6.900 1697.365 ;
        RECT 2906.300 1697.195 2906.740 1697.365 ;
        RECT 2912.720 1697.195 2914.100 1697.365 ;
        RECT 5.605 1696.105 6.815 1697.195 ;
        RECT 6.295 1695.565 6.815 1696.105 ;
        RECT 2912.805 1696.105 2914.015 1697.195 ;
        RECT 2912.805 1695.565 2913.325 1696.105 ;
        RECT 6.295 1693.015 6.815 1693.555 ;
        RECT 5.605 1691.925 6.815 1693.015 ;
        RECT 2906.365 1691.925 2906.655 1693.090 ;
        RECT 2912.805 1693.015 2913.325 1693.555 ;
        RECT 2912.805 1691.925 2914.015 1693.015 ;
        RECT 5.520 1691.755 6.900 1691.925 ;
        RECT 2906.300 1691.755 2906.740 1691.925 ;
        RECT 2912.720 1691.755 2914.100 1691.925 ;
        RECT 5.605 1690.665 6.815 1691.755 ;
        RECT 6.295 1690.125 6.815 1690.665 ;
        RECT 2912.805 1690.665 2914.015 1691.755 ;
        RECT 2912.805 1690.125 2913.325 1690.665 ;
        RECT 6.295 1687.575 6.815 1688.115 ;
        RECT 5.605 1686.485 6.815 1687.575 ;
        RECT 2906.365 1686.485 2906.655 1687.650 ;
        RECT 2912.805 1687.575 2913.325 1688.115 ;
        RECT 2912.805 1686.485 2914.015 1687.575 ;
        RECT 5.520 1686.315 6.900 1686.485 ;
        RECT 2906.300 1686.315 2906.740 1686.485 ;
        RECT 2912.720 1686.315 2914.100 1686.485 ;
        RECT 5.605 1685.225 6.815 1686.315 ;
        RECT 6.295 1684.685 6.815 1685.225 ;
        RECT 2912.805 1685.225 2914.015 1686.315 ;
        RECT 2912.805 1684.685 2913.325 1685.225 ;
        RECT 6.295 1682.135 6.815 1682.675 ;
        RECT 5.605 1681.045 6.815 1682.135 ;
        RECT 2906.365 1681.045 2906.655 1682.210 ;
        RECT 2912.805 1682.135 2913.325 1682.675 ;
        RECT 2912.805 1681.045 2914.015 1682.135 ;
        RECT 5.520 1680.875 6.900 1681.045 ;
        RECT 2906.300 1680.875 2906.740 1681.045 ;
        RECT 2912.720 1680.875 2914.100 1681.045 ;
        RECT 5.605 1679.785 6.815 1680.875 ;
        RECT 6.295 1679.245 6.815 1679.785 ;
        RECT 2912.805 1679.785 2914.015 1680.875 ;
        RECT 2912.805 1679.245 2913.325 1679.785 ;
        RECT 6.295 1676.695 6.815 1677.235 ;
        RECT 5.605 1675.605 6.815 1676.695 ;
        RECT 2906.365 1675.605 2906.655 1676.770 ;
        RECT 2912.805 1676.695 2913.325 1677.235 ;
        RECT 2912.805 1675.605 2914.015 1676.695 ;
        RECT 5.520 1675.435 6.900 1675.605 ;
        RECT 2906.300 1675.435 2906.740 1675.605 ;
        RECT 2912.720 1675.435 2914.100 1675.605 ;
        RECT 5.605 1674.345 6.815 1675.435 ;
        RECT 6.295 1673.805 6.815 1674.345 ;
        RECT 2912.805 1674.345 2914.015 1675.435 ;
        RECT 2912.805 1673.805 2913.325 1674.345 ;
        RECT 6.295 1671.255 6.815 1671.795 ;
        RECT 5.605 1670.165 6.815 1671.255 ;
        RECT 2906.365 1670.165 2906.655 1671.330 ;
        RECT 2912.805 1671.255 2913.325 1671.795 ;
        RECT 2909.315 1670.165 2909.645 1670.890 ;
        RECT 2912.805 1670.165 2914.015 1671.255 ;
        RECT 5.520 1669.995 6.900 1670.165 ;
        RECT 2906.300 1669.995 2906.740 1670.165 ;
        RECT 2909.040 1669.995 2910.420 1670.165 ;
        RECT 2912.720 1669.995 2914.100 1670.165 ;
        RECT 5.605 1668.905 6.815 1669.995 ;
        RECT 6.295 1668.365 6.815 1668.905 ;
        RECT 2912.805 1668.905 2914.015 1669.995 ;
        RECT 2912.805 1668.365 2913.325 1668.905 ;
        RECT 6.295 1665.815 6.815 1666.355 ;
        RECT 5.605 1664.725 6.815 1665.815 ;
        RECT 2906.365 1664.725 2906.655 1665.890 ;
        RECT 2912.805 1665.815 2913.325 1666.355 ;
        RECT 2912.805 1664.725 2914.015 1665.815 ;
        RECT 5.520 1664.555 6.900 1664.725 ;
        RECT 2906.300 1664.555 2906.740 1664.725 ;
        RECT 2912.720 1664.555 2914.100 1664.725 ;
        RECT 5.605 1663.465 6.815 1664.555 ;
        RECT 6.295 1662.925 6.815 1663.465 ;
        RECT 2912.805 1663.465 2914.015 1664.555 ;
        RECT 2912.805 1662.925 2913.325 1663.465 ;
        RECT 6.295 1660.375 6.815 1660.915 ;
        RECT 5.605 1659.285 6.815 1660.375 ;
        RECT 2906.365 1659.285 2906.655 1660.450 ;
        RECT 2912.805 1660.375 2913.325 1660.915 ;
        RECT 2912.805 1659.285 2914.015 1660.375 ;
        RECT 5.520 1659.115 6.900 1659.285 ;
        RECT 2906.300 1659.115 2906.740 1659.285 ;
        RECT 2912.720 1659.115 2914.100 1659.285 ;
        RECT 5.605 1658.025 6.815 1659.115 ;
        RECT 6.295 1657.485 6.815 1658.025 ;
        RECT 2912.805 1658.025 2914.015 1659.115 ;
        RECT 2912.805 1657.485 2913.325 1658.025 ;
        RECT 6.295 1654.935 6.815 1655.475 ;
        RECT 5.605 1653.845 6.815 1654.935 ;
        RECT 2906.365 1653.845 2906.655 1655.010 ;
        RECT 2912.805 1654.935 2913.325 1655.475 ;
        RECT 2912.805 1653.845 2914.015 1654.935 ;
        RECT 5.520 1653.675 6.900 1653.845 ;
        RECT 2906.300 1653.675 2906.740 1653.845 ;
        RECT 2912.720 1653.675 2914.100 1653.845 ;
        RECT 5.605 1652.585 6.815 1653.675 ;
        RECT 6.295 1652.045 6.815 1652.585 ;
        RECT 2912.805 1652.585 2914.015 1653.675 ;
        RECT 2912.805 1652.045 2913.325 1652.585 ;
        RECT 6.295 1649.495 6.815 1650.035 ;
        RECT 5.605 1648.405 6.815 1649.495 ;
        RECT 2906.365 1648.405 2906.655 1649.570 ;
        RECT 2912.805 1649.495 2913.325 1650.035 ;
        RECT 2912.805 1648.405 2914.015 1649.495 ;
        RECT 5.520 1648.235 6.900 1648.405 ;
        RECT 2906.300 1648.235 2906.740 1648.405 ;
        RECT 2912.720 1648.235 2914.100 1648.405 ;
        RECT 5.605 1647.145 6.815 1648.235 ;
        RECT 6.295 1646.605 6.815 1647.145 ;
        RECT 2912.805 1647.145 2914.015 1648.235 ;
        RECT 2912.805 1646.605 2913.325 1647.145 ;
        RECT 6.295 1644.055 6.815 1644.595 ;
        RECT 5.605 1642.965 6.815 1644.055 ;
        RECT 2906.365 1642.965 2906.655 1644.130 ;
        RECT 2912.805 1644.055 2913.325 1644.595 ;
        RECT 2912.805 1642.965 2914.015 1644.055 ;
        RECT 5.520 1642.795 6.900 1642.965 ;
        RECT 2906.300 1642.795 2906.740 1642.965 ;
        RECT 2912.720 1642.795 2914.100 1642.965 ;
        RECT 5.605 1641.705 6.815 1642.795 ;
        RECT 6.295 1641.165 6.815 1641.705 ;
        RECT 2912.805 1641.705 2914.015 1642.795 ;
        RECT 2912.805 1641.165 2913.325 1641.705 ;
        RECT 6.295 1638.615 6.815 1639.155 ;
        RECT 5.605 1637.525 6.815 1638.615 ;
        RECT 2906.365 1637.525 2906.655 1638.690 ;
        RECT 2912.805 1638.615 2913.325 1639.155 ;
        RECT 2912.805 1637.525 2914.015 1638.615 ;
        RECT 5.520 1637.355 6.900 1637.525 ;
        RECT 2906.300 1637.355 2906.740 1637.525 ;
        RECT 2912.720 1637.355 2914.100 1637.525 ;
        RECT 5.605 1636.265 6.815 1637.355 ;
        RECT 6.295 1635.725 6.815 1636.265 ;
        RECT 2912.805 1636.265 2914.015 1637.355 ;
        RECT 2912.805 1635.725 2913.325 1636.265 ;
        RECT 6.295 1633.175 6.815 1633.715 ;
        RECT 5.605 1632.085 6.815 1633.175 ;
        RECT 2906.365 1632.085 2906.655 1633.250 ;
        RECT 2912.805 1633.175 2913.325 1633.715 ;
        RECT 2912.805 1632.085 2914.015 1633.175 ;
        RECT 5.520 1631.915 6.900 1632.085 ;
        RECT 2906.300 1631.915 2906.740 1632.085 ;
        RECT 2912.720 1631.915 2914.100 1632.085 ;
        RECT 5.605 1630.825 6.815 1631.915 ;
        RECT 6.295 1630.285 6.815 1630.825 ;
        RECT 2912.805 1630.825 2914.015 1631.915 ;
        RECT 2912.805 1630.285 2913.325 1630.825 ;
        RECT 6.295 1627.735 6.815 1628.275 ;
        RECT 5.605 1626.645 6.815 1627.735 ;
        RECT 2906.365 1626.645 2906.655 1627.810 ;
        RECT 2912.805 1627.735 2913.325 1628.275 ;
        RECT 2912.805 1626.645 2914.015 1627.735 ;
        RECT 5.520 1626.475 6.900 1626.645 ;
        RECT 2906.300 1626.475 2906.740 1626.645 ;
        RECT 2912.720 1626.475 2914.100 1626.645 ;
        RECT 5.605 1625.385 6.815 1626.475 ;
        RECT 6.295 1624.845 6.815 1625.385 ;
        RECT 2912.805 1625.385 2914.015 1626.475 ;
        RECT 2912.805 1624.845 2913.325 1625.385 ;
        RECT 6.295 1622.295 6.815 1622.835 ;
        RECT 5.605 1621.205 6.815 1622.295 ;
        RECT 2906.365 1621.205 2906.655 1622.370 ;
        RECT 2912.805 1622.295 2913.325 1622.835 ;
        RECT 2912.805 1621.205 2914.015 1622.295 ;
        RECT 5.520 1621.035 6.900 1621.205 ;
        RECT 2906.300 1621.035 2906.740 1621.205 ;
        RECT 2912.720 1621.035 2914.100 1621.205 ;
        RECT 5.605 1619.945 6.815 1621.035 ;
        RECT 6.295 1619.405 6.815 1619.945 ;
        RECT 2912.805 1619.945 2914.015 1621.035 ;
        RECT 2912.805 1619.405 2913.325 1619.945 ;
        RECT 6.295 1616.855 6.815 1617.395 ;
        RECT 5.605 1615.765 6.815 1616.855 ;
        RECT 2906.365 1615.765 2906.655 1616.930 ;
        RECT 2912.805 1616.855 2913.325 1617.395 ;
        RECT 2912.805 1615.765 2914.015 1616.855 ;
        RECT 5.520 1615.595 6.900 1615.765 ;
        RECT 2906.300 1615.595 2906.740 1615.765 ;
        RECT 2912.720 1615.595 2914.100 1615.765 ;
        RECT 5.605 1614.505 6.815 1615.595 ;
        RECT 6.295 1613.965 6.815 1614.505 ;
        RECT 2912.805 1614.505 2914.015 1615.595 ;
        RECT 2912.805 1613.965 2913.325 1614.505 ;
        RECT 6.295 1611.415 6.815 1611.955 ;
        RECT 5.605 1610.325 6.815 1611.415 ;
        RECT 2906.365 1610.325 2906.655 1611.490 ;
        RECT 2912.805 1611.415 2913.325 1611.955 ;
        RECT 2912.805 1610.325 2914.015 1611.415 ;
        RECT 5.520 1610.155 6.900 1610.325 ;
        RECT 2906.300 1610.155 2906.740 1610.325 ;
        RECT 2912.720 1610.155 2914.100 1610.325 ;
        RECT 5.605 1609.065 6.815 1610.155 ;
        RECT 6.295 1608.525 6.815 1609.065 ;
        RECT 2912.805 1609.065 2914.015 1610.155 ;
        RECT 2912.805 1608.525 2913.325 1609.065 ;
        RECT 6.295 1605.975 6.815 1606.515 ;
        RECT 5.605 1604.885 6.815 1605.975 ;
        RECT 2906.365 1604.885 2906.655 1606.050 ;
        RECT 2912.805 1605.975 2913.325 1606.515 ;
        RECT 2912.805 1604.885 2914.015 1605.975 ;
        RECT 5.520 1604.715 6.900 1604.885 ;
        RECT 2906.300 1604.715 2906.740 1604.885 ;
        RECT 2912.720 1604.715 2914.100 1604.885 ;
        RECT 5.605 1603.625 6.815 1604.715 ;
        RECT 6.295 1603.085 6.815 1603.625 ;
        RECT 2912.805 1603.625 2914.015 1604.715 ;
        RECT 2912.805 1603.085 2913.325 1603.625 ;
        RECT 6.295 1600.535 6.815 1601.075 ;
        RECT 5.605 1599.445 6.815 1600.535 ;
        RECT 2906.365 1599.445 2906.655 1600.610 ;
        RECT 2912.805 1600.535 2913.325 1601.075 ;
        RECT 2912.805 1599.445 2914.015 1600.535 ;
        RECT 5.520 1599.275 6.900 1599.445 ;
        RECT 2906.300 1599.275 2906.740 1599.445 ;
        RECT 2912.720 1599.275 2914.100 1599.445 ;
        RECT 5.605 1598.185 6.815 1599.275 ;
        RECT 6.295 1597.645 6.815 1598.185 ;
        RECT 2912.805 1598.185 2914.015 1599.275 ;
        RECT 2912.805 1597.645 2913.325 1598.185 ;
        RECT 6.295 1595.095 6.815 1595.635 ;
        RECT 5.605 1594.005 6.815 1595.095 ;
        RECT 2906.365 1594.005 2906.655 1595.170 ;
        RECT 2912.805 1595.095 2913.325 1595.635 ;
        RECT 2912.805 1594.005 2914.015 1595.095 ;
        RECT 5.520 1593.835 6.900 1594.005 ;
        RECT 2906.300 1593.835 2906.740 1594.005 ;
        RECT 2912.720 1593.835 2914.100 1594.005 ;
        RECT 5.605 1592.745 6.815 1593.835 ;
        RECT 6.295 1592.205 6.815 1592.745 ;
        RECT 2912.805 1592.745 2914.015 1593.835 ;
        RECT 2912.805 1592.205 2913.325 1592.745 ;
        RECT 6.295 1589.655 6.815 1590.195 ;
        RECT 5.605 1588.565 6.815 1589.655 ;
        RECT 2906.365 1588.565 2906.655 1589.730 ;
        RECT 2912.805 1589.655 2913.325 1590.195 ;
        RECT 2912.805 1588.565 2914.015 1589.655 ;
        RECT 5.520 1588.395 6.900 1588.565 ;
        RECT 2906.300 1588.395 2906.740 1588.565 ;
        RECT 2912.720 1588.395 2914.100 1588.565 ;
        RECT 5.605 1587.305 6.815 1588.395 ;
        RECT 6.295 1586.765 6.815 1587.305 ;
        RECT 2912.805 1587.305 2914.015 1588.395 ;
        RECT 2912.805 1586.765 2913.325 1587.305 ;
        RECT 6.295 1584.215 6.815 1584.755 ;
        RECT 5.605 1583.125 6.815 1584.215 ;
        RECT 2906.365 1583.125 2906.655 1584.290 ;
        RECT 2912.805 1584.215 2913.325 1584.755 ;
        RECT 2912.805 1583.125 2914.015 1584.215 ;
        RECT 5.520 1582.955 6.900 1583.125 ;
        RECT 8.740 1582.955 10.120 1583.125 ;
        RECT 2906.300 1582.955 2906.740 1583.125 ;
        RECT 2912.720 1582.955 2914.100 1583.125 ;
        RECT 5.605 1581.865 6.815 1582.955 ;
        RECT 9.015 1582.230 9.345 1582.955 ;
        RECT 6.295 1581.325 6.815 1581.865 ;
        RECT 2912.805 1581.865 2914.015 1582.955 ;
        RECT 2912.805 1581.325 2913.325 1581.865 ;
        RECT 6.295 1578.775 6.815 1579.315 ;
        RECT 5.605 1577.685 6.815 1578.775 ;
        RECT 2906.365 1577.685 2906.655 1578.850 ;
        RECT 2912.805 1578.775 2913.325 1579.315 ;
        RECT 2912.805 1577.685 2914.015 1578.775 ;
        RECT 5.520 1577.515 6.900 1577.685 ;
        RECT 2906.300 1577.515 2906.740 1577.685 ;
        RECT 2912.720 1577.515 2914.100 1577.685 ;
        RECT 5.605 1576.425 6.815 1577.515 ;
        RECT 6.295 1575.885 6.815 1576.425 ;
        RECT 2912.805 1576.425 2914.015 1577.515 ;
        RECT 2912.805 1575.885 2913.325 1576.425 ;
        RECT 6.295 1573.335 6.815 1573.875 ;
        RECT 5.605 1572.245 6.815 1573.335 ;
        RECT 2906.365 1572.245 2906.655 1573.410 ;
        RECT 2912.805 1573.335 2913.325 1573.875 ;
        RECT 2912.805 1572.245 2914.015 1573.335 ;
        RECT 5.520 1572.075 6.900 1572.245 ;
        RECT 2906.300 1572.075 2906.740 1572.245 ;
        RECT 2912.720 1572.075 2914.100 1572.245 ;
        RECT 5.605 1570.985 6.815 1572.075 ;
        RECT 6.295 1570.445 6.815 1570.985 ;
        RECT 2912.805 1570.985 2914.015 1572.075 ;
        RECT 2912.805 1570.445 2913.325 1570.985 ;
        RECT 6.295 1567.895 6.815 1568.435 ;
        RECT 5.605 1566.805 6.815 1567.895 ;
        RECT 2906.365 1566.805 2906.655 1567.970 ;
        RECT 2912.805 1567.895 2913.325 1568.435 ;
        RECT 2912.805 1566.805 2914.015 1567.895 ;
        RECT 5.520 1566.635 6.900 1566.805 ;
        RECT 2906.300 1566.635 2906.740 1566.805 ;
        RECT 2912.720 1566.635 2914.100 1566.805 ;
        RECT 5.605 1565.545 6.815 1566.635 ;
        RECT 6.295 1565.005 6.815 1565.545 ;
        RECT 2912.805 1565.545 2914.015 1566.635 ;
        RECT 2912.805 1565.005 2913.325 1565.545 ;
        RECT 6.295 1562.455 6.815 1562.995 ;
        RECT 5.605 1561.365 6.815 1562.455 ;
        RECT 2906.365 1561.365 2906.655 1562.530 ;
        RECT 2912.805 1562.455 2913.325 1562.995 ;
        RECT 2912.805 1561.365 2914.015 1562.455 ;
        RECT 5.520 1561.195 6.900 1561.365 ;
        RECT 2906.300 1561.195 2906.740 1561.365 ;
        RECT 2912.720 1561.195 2914.100 1561.365 ;
        RECT 5.605 1560.105 6.815 1561.195 ;
        RECT 6.295 1559.565 6.815 1560.105 ;
        RECT 2912.805 1560.105 2914.015 1561.195 ;
        RECT 2912.805 1559.565 2913.325 1560.105 ;
        RECT 6.295 1557.015 6.815 1557.555 ;
        RECT 5.605 1555.925 6.815 1557.015 ;
        RECT 2906.365 1555.925 2906.655 1557.090 ;
        RECT 2912.805 1557.015 2913.325 1557.555 ;
        RECT 2912.805 1555.925 2914.015 1557.015 ;
        RECT 5.520 1555.755 6.900 1555.925 ;
        RECT 2906.300 1555.755 2906.740 1555.925 ;
        RECT 2912.720 1555.755 2914.100 1555.925 ;
        RECT 5.605 1554.665 6.815 1555.755 ;
        RECT 6.295 1554.125 6.815 1554.665 ;
        RECT 2912.805 1554.665 2914.015 1555.755 ;
        RECT 2912.805 1554.125 2913.325 1554.665 ;
        RECT 6.295 1551.575 6.815 1552.115 ;
        RECT 5.605 1550.485 6.815 1551.575 ;
        RECT 2906.365 1550.485 2906.655 1551.650 ;
        RECT 2912.805 1551.575 2913.325 1552.115 ;
        RECT 2912.805 1550.485 2914.015 1551.575 ;
        RECT 5.520 1550.315 6.900 1550.485 ;
        RECT 2906.300 1550.315 2906.740 1550.485 ;
        RECT 2912.720 1550.315 2914.100 1550.485 ;
        RECT 5.605 1549.225 6.815 1550.315 ;
        RECT 6.295 1548.685 6.815 1549.225 ;
        RECT 2912.805 1549.225 2914.015 1550.315 ;
        RECT 2912.805 1548.685 2913.325 1549.225 ;
        RECT 6.295 1546.135 6.815 1546.675 ;
        RECT 5.605 1545.045 6.815 1546.135 ;
        RECT 2906.365 1545.045 2906.655 1546.210 ;
        RECT 2912.805 1546.135 2913.325 1546.675 ;
        RECT 2912.805 1545.045 2914.015 1546.135 ;
        RECT 5.520 1544.875 6.900 1545.045 ;
        RECT 2906.300 1544.875 2906.740 1545.045 ;
        RECT 2912.720 1544.875 2914.100 1545.045 ;
        RECT 5.605 1543.785 6.815 1544.875 ;
        RECT 6.295 1543.245 6.815 1543.785 ;
        RECT 2912.805 1543.785 2914.015 1544.875 ;
        RECT 2912.805 1543.245 2913.325 1543.785 ;
        RECT 6.295 1540.695 6.815 1541.235 ;
        RECT 5.605 1539.605 6.815 1540.695 ;
        RECT 2906.365 1539.605 2906.655 1540.770 ;
        RECT 2912.805 1540.695 2913.325 1541.235 ;
        RECT 2912.805 1539.605 2914.015 1540.695 ;
        RECT 5.520 1539.435 6.900 1539.605 ;
        RECT 2906.300 1539.435 2906.740 1539.605 ;
        RECT 2912.720 1539.435 2914.100 1539.605 ;
        RECT 5.605 1538.345 6.815 1539.435 ;
        RECT 6.295 1537.805 6.815 1538.345 ;
        RECT 2912.805 1538.345 2914.015 1539.435 ;
        RECT 2912.805 1537.805 2913.325 1538.345 ;
        RECT 6.295 1535.255 6.815 1535.795 ;
        RECT 5.605 1534.165 6.815 1535.255 ;
        RECT 2906.365 1534.165 2906.655 1535.330 ;
        RECT 2912.805 1535.255 2913.325 1535.795 ;
        RECT 2912.805 1534.165 2914.015 1535.255 ;
        RECT 5.520 1533.995 6.900 1534.165 ;
        RECT 2906.300 1533.995 2906.740 1534.165 ;
        RECT 2912.720 1533.995 2914.100 1534.165 ;
        RECT 5.605 1532.905 6.815 1533.995 ;
        RECT 6.295 1532.365 6.815 1532.905 ;
        RECT 2912.805 1532.905 2914.015 1533.995 ;
        RECT 2912.805 1532.365 2913.325 1532.905 ;
        RECT 6.295 1529.815 6.815 1530.355 ;
        RECT 5.605 1528.725 6.815 1529.815 ;
        RECT 2906.365 1528.725 2906.655 1529.890 ;
        RECT 2912.805 1529.815 2913.325 1530.355 ;
        RECT 2912.805 1528.725 2914.015 1529.815 ;
        RECT 5.520 1528.555 6.900 1528.725 ;
        RECT 2906.300 1528.555 2906.740 1528.725 ;
        RECT 2909.040 1528.555 2910.420 1528.725 ;
        RECT 2912.720 1528.555 2914.100 1528.725 ;
        RECT 5.605 1527.465 6.815 1528.555 ;
        RECT 2909.315 1527.830 2909.645 1528.555 ;
        RECT 6.295 1526.925 6.815 1527.465 ;
        RECT 2912.805 1527.465 2914.015 1528.555 ;
        RECT 2912.805 1526.925 2913.325 1527.465 ;
        RECT 6.295 1524.375 6.815 1524.915 ;
        RECT 5.605 1523.285 6.815 1524.375 ;
        RECT 2906.365 1523.285 2906.655 1524.450 ;
        RECT 2912.805 1524.375 2913.325 1524.915 ;
        RECT 2912.805 1523.285 2914.015 1524.375 ;
        RECT 5.520 1523.115 6.900 1523.285 ;
        RECT 2906.300 1523.115 2906.740 1523.285 ;
        RECT 2912.720 1523.115 2914.100 1523.285 ;
        RECT 5.605 1522.025 6.815 1523.115 ;
        RECT 6.295 1521.485 6.815 1522.025 ;
        RECT 2912.805 1522.025 2914.015 1523.115 ;
        RECT 2912.805 1521.485 2913.325 1522.025 ;
        RECT 6.295 1518.935 6.815 1519.475 ;
        RECT 5.605 1517.845 6.815 1518.935 ;
        RECT 2906.365 1517.845 2906.655 1519.010 ;
        RECT 2912.805 1518.935 2913.325 1519.475 ;
        RECT 2912.805 1517.845 2914.015 1518.935 ;
        RECT 5.520 1517.675 6.900 1517.845 ;
        RECT 2906.300 1517.675 2906.740 1517.845 ;
        RECT 2909.040 1517.675 2910.420 1517.845 ;
        RECT 2912.720 1517.675 2914.100 1517.845 ;
        RECT 5.605 1516.585 6.815 1517.675 ;
        RECT 2909.315 1516.950 2909.645 1517.675 ;
        RECT 6.295 1516.045 6.815 1516.585 ;
        RECT 2912.805 1516.585 2914.015 1517.675 ;
        RECT 2912.805 1516.045 2913.325 1516.585 ;
        RECT 6.295 1513.495 6.815 1514.035 ;
        RECT 5.605 1512.405 6.815 1513.495 ;
        RECT 2906.365 1512.405 2906.655 1513.570 ;
        RECT 2912.805 1513.495 2913.325 1514.035 ;
        RECT 2912.805 1512.405 2914.015 1513.495 ;
        RECT 5.520 1512.235 6.900 1512.405 ;
        RECT 2906.300 1512.235 2906.740 1512.405 ;
        RECT 2912.720 1512.235 2914.100 1512.405 ;
        RECT 5.605 1511.145 6.815 1512.235 ;
        RECT 6.295 1510.605 6.815 1511.145 ;
        RECT 2912.805 1511.145 2914.015 1512.235 ;
        RECT 2912.805 1510.605 2913.325 1511.145 ;
        RECT 6.295 1508.055 6.815 1508.595 ;
        RECT 5.605 1506.965 6.815 1508.055 ;
        RECT 2906.365 1506.965 2906.655 1508.130 ;
        RECT 2912.805 1508.055 2913.325 1508.595 ;
        RECT 2912.805 1506.965 2914.015 1508.055 ;
        RECT 5.520 1506.795 6.900 1506.965 ;
        RECT 2906.300 1506.795 2906.740 1506.965 ;
        RECT 2912.720 1506.795 2914.100 1506.965 ;
        RECT 5.605 1505.705 6.815 1506.795 ;
        RECT 6.295 1505.165 6.815 1505.705 ;
        RECT 2912.805 1505.705 2914.015 1506.795 ;
        RECT 2912.805 1505.165 2913.325 1505.705 ;
        RECT 6.295 1502.615 6.815 1503.155 ;
        RECT 5.605 1501.525 6.815 1502.615 ;
        RECT 2906.365 1501.525 2906.655 1502.690 ;
        RECT 2912.805 1502.615 2913.325 1503.155 ;
        RECT 2912.805 1501.525 2914.015 1502.615 ;
        RECT 5.520 1501.355 6.900 1501.525 ;
        RECT 2906.300 1501.355 2906.740 1501.525 ;
        RECT 2912.720 1501.355 2914.100 1501.525 ;
        RECT 5.605 1500.265 6.815 1501.355 ;
        RECT 6.295 1499.725 6.815 1500.265 ;
        RECT 2912.805 1500.265 2914.015 1501.355 ;
        RECT 2912.805 1499.725 2913.325 1500.265 ;
        RECT 6.295 1497.175 6.815 1497.715 ;
        RECT 5.605 1496.085 6.815 1497.175 ;
        RECT 2906.365 1496.085 2906.655 1497.250 ;
        RECT 2912.805 1497.175 2913.325 1497.715 ;
        RECT 2912.805 1496.085 2914.015 1497.175 ;
        RECT 5.520 1495.915 6.900 1496.085 ;
        RECT 2906.300 1495.915 2906.740 1496.085 ;
        RECT 2912.720 1495.915 2914.100 1496.085 ;
        RECT 5.605 1494.825 6.815 1495.915 ;
        RECT 6.295 1494.285 6.815 1494.825 ;
        RECT 2912.805 1494.825 2914.015 1495.915 ;
        RECT 2912.805 1494.285 2913.325 1494.825 ;
        RECT 6.295 1491.735 6.815 1492.275 ;
        RECT 5.605 1490.645 6.815 1491.735 ;
        RECT 2906.365 1490.645 2906.655 1491.810 ;
        RECT 2912.805 1491.735 2913.325 1492.275 ;
        RECT 2912.805 1490.645 2914.015 1491.735 ;
        RECT 5.520 1490.475 6.900 1490.645 ;
        RECT 2906.300 1490.475 2906.740 1490.645 ;
        RECT 2912.720 1490.475 2914.100 1490.645 ;
        RECT 5.605 1489.385 6.815 1490.475 ;
        RECT 6.295 1488.845 6.815 1489.385 ;
        RECT 2912.805 1489.385 2914.015 1490.475 ;
        RECT 2912.805 1488.845 2913.325 1489.385 ;
        RECT 6.295 1486.295 6.815 1486.835 ;
        RECT 5.605 1485.205 6.815 1486.295 ;
        RECT 2906.365 1485.205 2906.655 1486.370 ;
        RECT 2912.805 1486.295 2913.325 1486.835 ;
        RECT 2912.805 1485.205 2914.015 1486.295 ;
        RECT 5.520 1485.035 6.900 1485.205 ;
        RECT 2906.300 1485.035 2906.740 1485.205 ;
        RECT 2912.720 1485.035 2914.100 1485.205 ;
        RECT 5.605 1483.945 6.815 1485.035 ;
        RECT 6.295 1483.405 6.815 1483.945 ;
        RECT 2912.805 1483.945 2914.015 1485.035 ;
        RECT 2912.805 1483.405 2913.325 1483.945 ;
        RECT 6.295 1480.855 6.815 1481.395 ;
        RECT 5.605 1479.765 6.815 1480.855 ;
        RECT 2906.365 1479.765 2906.655 1480.930 ;
        RECT 2912.805 1480.855 2913.325 1481.395 ;
        RECT 2912.805 1479.765 2914.015 1480.855 ;
        RECT 5.520 1479.595 6.900 1479.765 ;
        RECT 2906.300 1479.595 2906.740 1479.765 ;
        RECT 2912.720 1479.595 2914.100 1479.765 ;
        RECT 5.605 1478.505 6.815 1479.595 ;
        RECT 6.295 1477.965 6.815 1478.505 ;
        RECT 2912.805 1478.505 2914.015 1479.595 ;
        RECT 2912.805 1477.965 2913.325 1478.505 ;
        RECT 6.295 1475.415 6.815 1475.955 ;
        RECT 5.605 1474.325 6.815 1475.415 ;
        RECT 2906.365 1474.325 2906.655 1475.490 ;
        RECT 2912.805 1475.415 2913.325 1475.955 ;
        RECT 2912.805 1474.325 2914.015 1475.415 ;
        RECT 5.520 1474.155 6.900 1474.325 ;
        RECT 2906.300 1474.155 2906.740 1474.325 ;
        RECT 2909.040 1474.155 2910.420 1474.325 ;
        RECT 2912.720 1474.155 2914.100 1474.325 ;
        RECT 5.605 1473.065 6.815 1474.155 ;
        RECT 2909.315 1473.430 2909.645 1474.155 ;
        RECT 6.295 1472.525 6.815 1473.065 ;
        RECT 2912.805 1473.065 2914.015 1474.155 ;
        RECT 2912.805 1472.525 2913.325 1473.065 ;
        RECT 6.295 1469.975 6.815 1470.515 ;
        RECT 5.605 1468.885 6.815 1469.975 ;
        RECT 2906.365 1468.885 2906.655 1470.050 ;
        RECT 2912.805 1469.975 2913.325 1470.515 ;
        RECT 2912.805 1468.885 2914.015 1469.975 ;
        RECT 5.520 1468.715 6.900 1468.885 ;
        RECT 2906.300 1468.715 2906.740 1468.885 ;
        RECT 2912.720 1468.715 2914.100 1468.885 ;
        RECT 5.605 1467.625 6.815 1468.715 ;
        RECT 6.295 1467.085 6.815 1467.625 ;
        RECT 2912.805 1467.625 2914.015 1468.715 ;
        RECT 2912.805 1467.085 2913.325 1467.625 ;
        RECT 6.295 1464.535 6.815 1465.075 ;
        RECT 5.605 1463.445 6.815 1464.535 ;
        RECT 2906.365 1463.445 2906.655 1464.610 ;
        RECT 2912.805 1464.535 2913.325 1465.075 ;
        RECT 2912.805 1463.445 2914.015 1464.535 ;
        RECT 5.520 1463.275 6.900 1463.445 ;
        RECT 2906.300 1463.275 2906.740 1463.445 ;
        RECT 2912.720 1463.275 2914.100 1463.445 ;
        RECT 5.605 1462.185 6.815 1463.275 ;
        RECT 6.295 1461.645 6.815 1462.185 ;
        RECT 2912.805 1462.185 2914.015 1463.275 ;
        RECT 2912.805 1461.645 2913.325 1462.185 ;
        RECT 6.295 1459.095 6.815 1459.635 ;
        RECT 5.605 1458.005 6.815 1459.095 ;
        RECT 2906.365 1458.005 2906.655 1459.170 ;
        RECT 2912.805 1459.095 2913.325 1459.635 ;
        RECT 2912.805 1458.005 2914.015 1459.095 ;
        RECT 5.520 1457.835 6.900 1458.005 ;
        RECT 2906.300 1457.835 2906.740 1458.005 ;
        RECT 2912.720 1457.835 2914.100 1458.005 ;
        RECT 5.605 1456.745 6.815 1457.835 ;
        RECT 6.295 1456.205 6.815 1456.745 ;
        RECT 2912.805 1456.745 2914.015 1457.835 ;
        RECT 2912.805 1456.205 2913.325 1456.745 ;
        RECT 6.295 1453.655 6.815 1454.195 ;
        RECT 5.605 1452.565 6.815 1453.655 ;
        RECT 2906.365 1452.565 2906.655 1453.730 ;
        RECT 2912.805 1453.655 2913.325 1454.195 ;
        RECT 2912.805 1452.565 2914.015 1453.655 ;
        RECT 5.520 1452.395 6.900 1452.565 ;
        RECT 2906.300 1452.395 2906.740 1452.565 ;
        RECT 2912.720 1452.395 2914.100 1452.565 ;
        RECT 5.605 1451.305 6.815 1452.395 ;
        RECT 6.295 1450.765 6.815 1451.305 ;
        RECT 2912.805 1451.305 2914.015 1452.395 ;
        RECT 2912.805 1450.765 2913.325 1451.305 ;
        RECT 6.295 1448.215 6.815 1448.755 ;
        RECT 5.605 1447.125 6.815 1448.215 ;
        RECT 2906.365 1447.125 2906.655 1448.290 ;
        RECT 2912.805 1448.215 2913.325 1448.755 ;
        RECT 2912.805 1447.125 2914.015 1448.215 ;
        RECT 5.520 1446.955 6.900 1447.125 ;
        RECT 2906.300 1446.955 2906.740 1447.125 ;
        RECT 2912.720 1446.955 2914.100 1447.125 ;
        RECT 5.605 1445.865 6.815 1446.955 ;
        RECT 6.295 1445.325 6.815 1445.865 ;
        RECT 2912.805 1445.865 2914.015 1446.955 ;
        RECT 2912.805 1445.325 2913.325 1445.865 ;
        RECT 6.295 1442.775 6.815 1443.315 ;
        RECT 5.605 1441.685 6.815 1442.775 ;
        RECT 2906.365 1441.685 2906.655 1442.850 ;
        RECT 2912.805 1442.775 2913.325 1443.315 ;
        RECT 2912.805 1441.685 2914.015 1442.775 ;
        RECT 5.520 1441.515 6.900 1441.685 ;
        RECT 2906.300 1441.515 2906.740 1441.685 ;
        RECT 2912.720 1441.515 2914.100 1441.685 ;
        RECT 5.605 1440.425 6.815 1441.515 ;
        RECT 6.295 1439.885 6.815 1440.425 ;
        RECT 2912.805 1440.425 2914.015 1441.515 ;
        RECT 2912.805 1439.885 2913.325 1440.425 ;
        RECT 6.295 1437.335 6.815 1437.875 ;
        RECT 5.605 1436.245 6.815 1437.335 ;
        RECT 2906.365 1436.245 2906.655 1437.410 ;
        RECT 2912.805 1437.335 2913.325 1437.875 ;
        RECT 2912.805 1436.245 2914.015 1437.335 ;
        RECT 5.520 1436.075 6.900 1436.245 ;
        RECT 2906.300 1436.075 2906.740 1436.245 ;
        RECT 2912.720 1436.075 2914.100 1436.245 ;
        RECT 5.605 1434.985 6.815 1436.075 ;
        RECT 6.295 1434.445 6.815 1434.985 ;
        RECT 2912.805 1434.985 2914.015 1436.075 ;
        RECT 2912.805 1434.445 2913.325 1434.985 ;
        RECT 6.295 1431.895 6.815 1432.435 ;
        RECT 5.605 1430.805 6.815 1431.895 ;
        RECT 2906.365 1430.805 2906.655 1431.970 ;
        RECT 2912.805 1431.895 2913.325 1432.435 ;
        RECT 2912.805 1430.805 2914.015 1431.895 ;
        RECT 5.520 1430.635 6.900 1430.805 ;
        RECT 2906.300 1430.635 2906.740 1430.805 ;
        RECT 2912.720 1430.635 2914.100 1430.805 ;
        RECT 5.605 1429.545 6.815 1430.635 ;
        RECT 6.295 1429.005 6.815 1429.545 ;
        RECT 2912.805 1429.545 2914.015 1430.635 ;
        RECT 2912.805 1429.005 2913.325 1429.545 ;
        RECT 6.295 1426.455 6.815 1426.995 ;
        RECT 5.605 1425.365 6.815 1426.455 ;
        RECT 2906.365 1425.365 2906.655 1426.530 ;
        RECT 2912.805 1426.455 2913.325 1426.995 ;
        RECT 2912.805 1425.365 2914.015 1426.455 ;
        RECT 5.520 1425.195 6.900 1425.365 ;
        RECT 2906.300 1425.195 2906.740 1425.365 ;
        RECT 2912.720 1425.195 2914.100 1425.365 ;
        RECT 5.605 1424.105 6.815 1425.195 ;
        RECT 6.295 1423.565 6.815 1424.105 ;
        RECT 2912.805 1424.105 2914.015 1425.195 ;
        RECT 2912.805 1423.565 2913.325 1424.105 ;
        RECT 6.295 1421.015 6.815 1421.555 ;
        RECT 5.605 1419.925 6.815 1421.015 ;
        RECT 2906.365 1419.925 2906.655 1421.090 ;
        RECT 2912.805 1421.015 2913.325 1421.555 ;
        RECT 2912.805 1419.925 2914.015 1421.015 ;
        RECT 5.520 1419.755 6.900 1419.925 ;
        RECT 2906.300 1419.755 2906.740 1419.925 ;
        RECT 2912.720 1419.755 2914.100 1419.925 ;
        RECT 5.605 1418.665 6.815 1419.755 ;
        RECT 6.295 1418.125 6.815 1418.665 ;
        RECT 2912.805 1418.665 2914.015 1419.755 ;
        RECT 2912.805 1418.125 2913.325 1418.665 ;
        RECT 6.295 1415.575 6.815 1416.115 ;
        RECT 5.605 1414.485 6.815 1415.575 ;
        RECT 2906.365 1414.485 2906.655 1415.650 ;
        RECT 2912.805 1415.575 2913.325 1416.115 ;
        RECT 2912.805 1414.485 2914.015 1415.575 ;
        RECT 5.520 1414.315 6.900 1414.485 ;
        RECT 2906.300 1414.315 2906.740 1414.485 ;
        RECT 2912.720 1414.315 2914.100 1414.485 ;
        RECT 5.605 1413.225 6.815 1414.315 ;
        RECT 6.295 1412.685 6.815 1413.225 ;
        RECT 2912.805 1413.225 2914.015 1414.315 ;
        RECT 2912.805 1412.685 2913.325 1413.225 ;
        RECT 6.295 1410.135 6.815 1410.675 ;
        RECT 5.605 1409.045 6.815 1410.135 ;
        RECT 2906.365 1409.045 2906.655 1410.210 ;
        RECT 2912.805 1410.135 2913.325 1410.675 ;
        RECT 2912.805 1409.045 2914.015 1410.135 ;
        RECT 5.520 1408.875 6.900 1409.045 ;
        RECT 2906.300 1408.875 2906.740 1409.045 ;
        RECT 2912.720 1408.875 2914.100 1409.045 ;
        RECT 5.605 1407.785 6.815 1408.875 ;
        RECT 6.295 1407.245 6.815 1407.785 ;
        RECT 2912.805 1407.785 2914.015 1408.875 ;
        RECT 2912.805 1407.245 2913.325 1407.785 ;
        RECT 6.295 1404.695 6.815 1405.235 ;
        RECT 5.605 1403.605 6.815 1404.695 ;
        RECT 2906.365 1403.605 2906.655 1404.770 ;
        RECT 2912.805 1404.695 2913.325 1405.235 ;
        RECT 2912.805 1403.605 2914.015 1404.695 ;
        RECT 5.520 1403.435 6.900 1403.605 ;
        RECT 2906.300 1403.435 2906.740 1403.605 ;
        RECT 2912.720 1403.435 2914.100 1403.605 ;
        RECT 5.605 1402.345 6.815 1403.435 ;
        RECT 6.295 1401.805 6.815 1402.345 ;
        RECT 2912.805 1402.345 2914.015 1403.435 ;
        RECT 2912.805 1401.805 2913.325 1402.345 ;
        RECT 6.295 1399.255 6.815 1399.795 ;
        RECT 5.605 1398.165 6.815 1399.255 ;
        RECT 2906.365 1398.165 2906.655 1399.330 ;
        RECT 2912.805 1399.255 2913.325 1399.795 ;
        RECT 2912.805 1398.165 2914.015 1399.255 ;
        RECT 5.520 1397.995 6.900 1398.165 ;
        RECT 2906.300 1397.995 2906.740 1398.165 ;
        RECT 2912.720 1397.995 2914.100 1398.165 ;
        RECT 5.605 1396.905 6.815 1397.995 ;
        RECT 6.295 1396.365 6.815 1396.905 ;
        RECT 2912.805 1396.905 2914.015 1397.995 ;
        RECT 2912.805 1396.365 2913.325 1396.905 ;
        RECT 6.295 1393.815 6.815 1394.355 ;
        RECT 5.605 1392.725 6.815 1393.815 ;
        RECT 2906.365 1392.725 2906.655 1393.890 ;
        RECT 2912.805 1393.815 2913.325 1394.355 ;
        RECT 2912.805 1392.725 2914.015 1393.815 ;
        RECT 5.520 1392.555 6.900 1392.725 ;
        RECT 2906.300 1392.555 2906.740 1392.725 ;
        RECT 2912.720 1392.555 2914.100 1392.725 ;
        RECT 5.605 1391.465 6.815 1392.555 ;
        RECT 6.295 1390.925 6.815 1391.465 ;
        RECT 2912.805 1391.465 2914.015 1392.555 ;
        RECT 2912.805 1390.925 2913.325 1391.465 ;
        RECT 6.295 1388.375 6.815 1388.915 ;
        RECT 5.605 1387.285 6.815 1388.375 ;
        RECT 2906.365 1387.285 2906.655 1388.450 ;
        RECT 2912.805 1388.375 2913.325 1388.915 ;
        RECT 2912.805 1387.285 2914.015 1388.375 ;
        RECT 5.520 1387.115 6.900 1387.285 ;
        RECT 2906.300 1387.115 2906.740 1387.285 ;
        RECT 2912.720 1387.115 2914.100 1387.285 ;
        RECT 5.605 1386.025 6.815 1387.115 ;
        RECT 6.295 1385.485 6.815 1386.025 ;
        RECT 2912.805 1386.025 2914.015 1387.115 ;
        RECT 2912.805 1385.485 2913.325 1386.025 ;
        RECT 6.295 1382.935 6.815 1383.475 ;
        RECT 5.605 1381.845 6.815 1382.935 ;
        RECT 2906.365 1381.845 2906.655 1383.010 ;
        RECT 2912.805 1382.935 2913.325 1383.475 ;
        RECT 2912.805 1381.845 2914.015 1382.935 ;
        RECT 5.520 1381.675 6.900 1381.845 ;
        RECT 2906.300 1381.675 2906.740 1381.845 ;
        RECT 2912.720 1381.675 2914.100 1381.845 ;
        RECT 5.605 1380.585 6.815 1381.675 ;
        RECT 6.295 1380.045 6.815 1380.585 ;
        RECT 2912.805 1380.585 2914.015 1381.675 ;
        RECT 2912.805 1380.045 2913.325 1380.585 ;
        RECT 6.295 1377.495 6.815 1378.035 ;
        RECT 5.605 1376.405 6.815 1377.495 ;
        RECT 2906.365 1376.405 2906.655 1377.570 ;
        RECT 2912.805 1377.495 2913.325 1378.035 ;
        RECT 2912.805 1376.405 2914.015 1377.495 ;
        RECT 5.520 1376.235 6.900 1376.405 ;
        RECT 2906.300 1376.235 2906.740 1376.405 ;
        RECT 2912.720 1376.235 2914.100 1376.405 ;
        RECT 5.605 1375.145 6.815 1376.235 ;
        RECT 6.295 1374.605 6.815 1375.145 ;
        RECT 2912.805 1375.145 2914.015 1376.235 ;
        RECT 2912.805 1374.605 2913.325 1375.145 ;
        RECT 6.295 1372.055 6.815 1372.595 ;
        RECT 5.605 1370.965 6.815 1372.055 ;
        RECT 2906.365 1370.965 2906.655 1372.130 ;
        RECT 2912.805 1372.055 2913.325 1372.595 ;
        RECT 2912.805 1370.965 2914.015 1372.055 ;
        RECT 5.520 1370.795 6.900 1370.965 ;
        RECT 2906.300 1370.795 2906.740 1370.965 ;
        RECT 2912.720 1370.795 2914.100 1370.965 ;
        RECT 5.605 1369.705 6.815 1370.795 ;
        RECT 6.295 1369.165 6.815 1369.705 ;
        RECT 2912.805 1369.705 2914.015 1370.795 ;
        RECT 2912.805 1369.165 2913.325 1369.705 ;
        RECT 6.295 1366.615 6.815 1367.155 ;
        RECT 5.605 1365.525 6.815 1366.615 ;
        RECT 2906.365 1365.525 2906.655 1366.690 ;
        RECT 2912.805 1366.615 2913.325 1367.155 ;
        RECT 2912.805 1365.525 2914.015 1366.615 ;
        RECT 5.520 1365.355 6.900 1365.525 ;
        RECT 2906.300 1365.355 2906.740 1365.525 ;
        RECT 2912.720 1365.355 2914.100 1365.525 ;
        RECT 5.605 1364.265 6.815 1365.355 ;
        RECT 6.295 1363.725 6.815 1364.265 ;
        RECT 2912.805 1364.265 2914.015 1365.355 ;
        RECT 2912.805 1363.725 2913.325 1364.265 ;
        RECT 6.295 1361.175 6.815 1361.715 ;
        RECT 5.605 1360.085 6.815 1361.175 ;
        RECT 2906.365 1360.085 2906.655 1361.250 ;
        RECT 2912.805 1361.175 2913.325 1361.715 ;
        RECT 2912.805 1360.085 2914.015 1361.175 ;
        RECT 5.520 1359.915 6.900 1360.085 ;
        RECT 2906.300 1359.915 2906.740 1360.085 ;
        RECT 2912.720 1359.915 2914.100 1360.085 ;
        RECT 5.605 1358.825 6.815 1359.915 ;
        RECT 6.295 1358.285 6.815 1358.825 ;
        RECT 2912.805 1358.825 2914.015 1359.915 ;
        RECT 2912.805 1358.285 2913.325 1358.825 ;
        RECT 6.295 1355.735 6.815 1356.275 ;
        RECT 5.605 1354.645 6.815 1355.735 ;
        RECT 2906.365 1354.645 2906.655 1355.810 ;
        RECT 2912.805 1355.735 2913.325 1356.275 ;
        RECT 2912.805 1354.645 2914.015 1355.735 ;
        RECT 5.520 1354.475 6.900 1354.645 ;
        RECT 2906.300 1354.475 2906.740 1354.645 ;
        RECT 2912.720 1354.475 2914.100 1354.645 ;
        RECT 5.605 1353.385 6.815 1354.475 ;
        RECT 6.295 1352.845 6.815 1353.385 ;
        RECT 2912.805 1353.385 2914.015 1354.475 ;
        RECT 2912.805 1352.845 2913.325 1353.385 ;
        RECT 6.295 1350.295 6.815 1350.835 ;
        RECT 5.605 1349.205 6.815 1350.295 ;
        RECT 2906.365 1349.205 2906.655 1350.370 ;
        RECT 2912.805 1350.295 2913.325 1350.835 ;
        RECT 2912.805 1349.205 2914.015 1350.295 ;
        RECT 5.520 1349.035 6.900 1349.205 ;
        RECT 2906.300 1349.035 2906.740 1349.205 ;
        RECT 2912.720 1349.035 2914.100 1349.205 ;
        RECT 5.605 1347.945 6.815 1349.035 ;
        RECT 6.295 1347.405 6.815 1347.945 ;
        RECT 2912.805 1347.945 2914.015 1349.035 ;
        RECT 2912.805 1347.405 2913.325 1347.945 ;
        RECT 6.295 1344.855 6.815 1345.395 ;
        RECT 5.605 1343.765 6.815 1344.855 ;
        RECT 2906.365 1343.765 2906.655 1344.930 ;
        RECT 2912.805 1344.855 2913.325 1345.395 ;
        RECT 2912.805 1343.765 2914.015 1344.855 ;
        RECT 5.520 1343.595 6.900 1343.765 ;
        RECT 2906.300 1343.595 2906.740 1343.765 ;
        RECT 2912.720 1343.595 2914.100 1343.765 ;
        RECT 5.605 1342.505 6.815 1343.595 ;
        RECT 6.295 1341.965 6.815 1342.505 ;
        RECT 2912.805 1342.505 2914.015 1343.595 ;
        RECT 2912.805 1341.965 2913.325 1342.505 ;
        RECT 6.295 1339.415 6.815 1339.955 ;
        RECT 5.605 1338.325 6.815 1339.415 ;
        RECT 2906.365 1338.325 2906.655 1339.490 ;
        RECT 2912.805 1339.415 2913.325 1339.955 ;
        RECT 2912.805 1338.325 2914.015 1339.415 ;
        RECT 5.520 1338.155 6.900 1338.325 ;
        RECT 2906.300 1338.155 2906.740 1338.325 ;
        RECT 2912.720 1338.155 2914.100 1338.325 ;
        RECT 5.605 1337.065 6.815 1338.155 ;
        RECT 6.295 1336.525 6.815 1337.065 ;
        RECT 2912.805 1337.065 2914.015 1338.155 ;
        RECT 2912.805 1336.525 2913.325 1337.065 ;
        RECT 6.295 1333.975 6.815 1334.515 ;
        RECT 5.605 1332.885 6.815 1333.975 ;
        RECT 2906.365 1332.885 2906.655 1334.050 ;
        RECT 2912.805 1333.975 2913.325 1334.515 ;
        RECT 2912.805 1332.885 2914.015 1333.975 ;
        RECT 5.520 1332.715 6.900 1332.885 ;
        RECT 2906.300 1332.715 2906.740 1332.885 ;
        RECT 2912.720 1332.715 2914.100 1332.885 ;
        RECT 5.605 1331.625 6.815 1332.715 ;
        RECT 6.295 1331.085 6.815 1331.625 ;
        RECT 2912.805 1331.625 2914.015 1332.715 ;
        RECT 2912.805 1331.085 2913.325 1331.625 ;
        RECT 6.295 1328.535 6.815 1329.075 ;
        RECT 5.605 1327.445 6.815 1328.535 ;
        RECT 9.015 1327.445 9.345 1328.170 ;
        RECT 2906.365 1327.445 2906.655 1328.610 ;
        RECT 2912.805 1328.535 2913.325 1329.075 ;
        RECT 2912.805 1327.445 2914.015 1328.535 ;
        RECT 5.520 1327.275 6.900 1327.445 ;
        RECT 8.740 1327.275 10.120 1327.445 ;
        RECT 2906.300 1327.275 2906.740 1327.445 ;
        RECT 2912.720 1327.275 2914.100 1327.445 ;
        RECT 5.605 1326.185 6.815 1327.275 ;
        RECT 6.295 1325.645 6.815 1326.185 ;
        RECT 2912.805 1326.185 2914.015 1327.275 ;
        RECT 2912.805 1325.645 2913.325 1326.185 ;
        RECT 6.295 1323.095 6.815 1323.635 ;
        RECT 5.605 1322.005 6.815 1323.095 ;
        RECT 2906.365 1322.005 2906.655 1323.170 ;
        RECT 2912.805 1323.095 2913.325 1323.635 ;
        RECT 2912.805 1322.005 2914.015 1323.095 ;
        RECT 5.520 1321.835 6.900 1322.005 ;
        RECT 2906.300 1321.835 2906.740 1322.005 ;
        RECT 2912.720 1321.835 2914.100 1322.005 ;
        RECT 5.605 1320.745 6.815 1321.835 ;
        RECT 6.295 1320.205 6.815 1320.745 ;
        RECT 2912.805 1320.745 2914.015 1321.835 ;
        RECT 2912.805 1320.205 2913.325 1320.745 ;
        RECT 6.295 1317.655 6.815 1318.195 ;
        RECT 5.605 1316.565 6.815 1317.655 ;
        RECT 2906.365 1316.565 2906.655 1317.730 ;
        RECT 2912.805 1317.655 2913.325 1318.195 ;
        RECT 2912.805 1316.565 2914.015 1317.655 ;
        RECT 5.520 1316.395 6.900 1316.565 ;
        RECT 2906.300 1316.395 2906.740 1316.565 ;
        RECT 2912.720 1316.395 2914.100 1316.565 ;
        RECT 5.605 1315.305 6.815 1316.395 ;
        RECT 6.295 1314.765 6.815 1315.305 ;
        RECT 2912.805 1315.305 2914.015 1316.395 ;
        RECT 2912.805 1314.765 2913.325 1315.305 ;
        RECT 6.295 1312.215 6.815 1312.755 ;
        RECT 5.605 1311.125 6.815 1312.215 ;
        RECT 2906.365 1311.125 2906.655 1312.290 ;
        RECT 2912.805 1312.215 2913.325 1312.755 ;
        RECT 2912.805 1311.125 2914.015 1312.215 ;
        RECT 5.520 1310.955 6.900 1311.125 ;
        RECT 2906.300 1310.955 2906.740 1311.125 ;
        RECT 2912.720 1310.955 2914.100 1311.125 ;
        RECT 5.605 1309.865 6.815 1310.955 ;
        RECT 6.295 1309.325 6.815 1309.865 ;
        RECT 2912.805 1309.865 2914.015 1310.955 ;
        RECT 2912.805 1309.325 2913.325 1309.865 ;
        RECT 6.295 1306.775 6.815 1307.315 ;
        RECT 5.605 1305.685 6.815 1306.775 ;
        RECT 2906.365 1305.685 2906.655 1306.850 ;
        RECT 2912.805 1306.775 2913.325 1307.315 ;
        RECT 2912.805 1305.685 2914.015 1306.775 ;
        RECT 5.520 1305.515 6.900 1305.685 ;
        RECT 2906.300 1305.515 2906.740 1305.685 ;
        RECT 2912.720 1305.515 2914.100 1305.685 ;
        RECT 5.605 1304.425 6.815 1305.515 ;
        RECT 6.295 1303.885 6.815 1304.425 ;
        RECT 2912.805 1304.425 2914.015 1305.515 ;
        RECT 2912.805 1303.885 2913.325 1304.425 ;
        RECT 6.295 1301.335 6.815 1301.875 ;
        RECT 5.605 1300.245 6.815 1301.335 ;
        RECT 2906.365 1300.245 2906.655 1301.410 ;
        RECT 2912.805 1301.335 2913.325 1301.875 ;
        RECT 2909.315 1300.245 2909.645 1300.970 ;
        RECT 2912.805 1300.245 2914.015 1301.335 ;
        RECT 5.520 1300.075 6.900 1300.245 ;
        RECT 2906.300 1300.075 2906.740 1300.245 ;
        RECT 2909.040 1300.075 2910.420 1300.245 ;
        RECT 2912.720 1300.075 2914.100 1300.245 ;
        RECT 5.605 1298.985 6.815 1300.075 ;
        RECT 6.295 1298.445 6.815 1298.985 ;
        RECT 2912.805 1298.985 2914.015 1300.075 ;
        RECT 2912.805 1298.445 2913.325 1298.985 ;
        RECT 6.295 1295.895 6.815 1296.435 ;
        RECT 5.605 1294.805 6.815 1295.895 ;
        RECT 2906.365 1294.805 2906.655 1295.970 ;
        RECT 2912.805 1295.895 2913.325 1296.435 ;
        RECT 2912.805 1294.805 2914.015 1295.895 ;
        RECT 5.520 1294.635 6.900 1294.805 ;
        RECT 2906.300 1294.635 2906.740 1294.805 ;
        RECT 2912.720 1294.635 2914.100 1294.805 ;
        RECT 5.605 1293.545 6.815 1294.635 ;
        RECT 6.295 1293.005 6.815 1293.545 ;
        RECT 2912.805 1293.545 2914.015 1294.635 ;
        RECT 2912.805 1293.005 2913.325 1293.545 ;
        RECT 6.295 1290.455 6.815 1290.995 ;
        RECT 5.605 1289.365 6.815 1290.455 ;
        RECT 2906.365 1289.365 2906.655 1290.530 ;
        RECT 2912.805 1290.455 2913.325 1290.995 ;
        RECT 2912.805 1289.365 2914.015 1290.455 ;
        RECT 5.520 1289.195 6.900 1289.365 ;
        RECT 2906.300 1289.195 2906.740 1289.365 ;
        RECT 2912.720 1289.195 2914.100 1289.365 ;
        RECT 5.605 1288.105 6.815 1289.195 ;
        RECT 6.295 1287.565 6.815 1288.105 ;
        RECT 2912.805 1288.105 2914.015 1289.195 ;
        RECT 2912.805 1287.565 2913.325 1288.105 ;
        RECT 6.295 1285.015 6.815 1285.555 ;
        RECT 5.605 1283.925 6.815 1285.015 ;
        RECT 9.015 1283.925 9.345 1284.650 ;
        RECT 2906.365 1283.925 2906.655 1285.090 ;
        RECT 2912.805 1285.015 2913.325 1285.555 ;
        RECT 2912.805 1283.925 2914.015 1285.015 ;
        RECT 5.520 1283.755 6.900 1283.925 ;
        RECT 8.740 1283.755 10.120 1283.925 ;
        RECT 2906.300 1283.755 2906.740 1283.925 ;
        RECT 2912.720 1283.755 2914.100 1283.925 ;
        RECT 5.605 1282.665 6.815 1283.755 ;
        RECT 6.295 1282.125 6.815 1282.665 ;
        RECT 2912.805 1282.665 2914.015 1283.755 ;
        RECT 2912.805 1282.125 2913.325 1282.665 ;
        RECT 6.295 1279.575 6.815 1280.115 ;
        RECT 5.605 1278.485 6.815 1279.575 ;
        RECT 2906.365 1278.485 2906.655 1279.650 ;
        RECT 2912.805 1279.575 2913.325 1280.115 ;
        RECT 2912.805 1278.485 2914.015 1279.575 ;
        RECT 5.520 1278.315 6.900 1278.485 ;
        RECT 2906.300 1278.315 2906.740 1278.485 ;
        RECT 2912.720 1278.315 2914.100 1278.485 ;
        RECT 5.605 1277.225 6.815 1278.315 ;
        RECT 6.295 1276.685 6.815 1277.225 ;
        RECT 2912.805 1277.225 2914.015 1278.315 ;
        RECT 2912.805 1276.685 2913.325 1277.225 ;
        RECT 6.295 1274.135 6.815 1274.675 ;
        RECT 5.605 1273.045 6.815 1274.135 ;
        RECT 9.015 1273.045 9.345 1273.770 ;
        RECT 2906.365 1273.045 2906.655 1274.210 ;
        RECT 2912.805 1274.135 2913.325 1274.675 ;
        RECT 2912.805 1273.045 2914.015 1274.135 ;
        RECT 5.520 1272.875 6.900 1273.045 ;
        RECT 8.740 1272.875 10.120 1273.045 ;
        RECT 2906.300 1272.875 2906.740 1273.045 ;
        RECT 2912.720 1272.875 2914.100 1273.045 ;
        RECT 5.605 1271.785 6.815 1272.875 ;
        RECT 6.295 1271.245 6.815 1271.785 ;
        RECT 2912.805 1271.785 2914.015 1272.875 ;
        RECT 2912.805 1271.245 2913.325 1271.785 ;
        RECT 6.295 1268.695 6.815 1269.235 ;
        RECT 5.605 1267.605 6.815 1268.695 ;
        RECT 2906.365 1267.605 2906.655 1268.770 ;
        RECT 2912.805 1268.695 2913.325 1269.235 ;
        RECT 2912.805 1267.605 2914.015 1268.695 ;
        RECT 5.520 1267.435 6.900 1267.605 ;
        RECT 2906.300 1267.435 2906.740 1267.605 ;
        RECT 2909.040 1267.435 2910.420 1267.605 ;
        RECT 2912.720 1267.435 2914.100 1267.605 ;
        RECT 5.605 1266.345 6.815 1267.435 ;
        RECT 2909.315 1266.710 2909.645 1267.435 ;
        RECT 6.295 1265.805 6.815 1266.345 ;
        RECT 2912.805 1266.345 2914.015 1267.435 ;
        RECT 2912.805 1265.805 2913.325 1266.345 ;
        RECT 6.295 1263.255 6.815 1263.795 ;
        RECT 5.605 1262.165 6.815 1263.255 ;
        RECT 2906.365 1262.165 2906.655 1263.330 ;
        RECT 2912.805 1263.255 2913.325 1263.795 ;
        RECT 2912.805 1262.165 2914.015 1263.255 ;
        RECT 5.520 1261.995 6.900 1262.165 ;
        RECT 2906.300 1261.995 2906.740 1262.165 ;
        RECT 2912.720 1261.995 2914.100 1262.165 ;
        RECT 5.605 1260.905 6.815 1261.995 ;
        RECT 6.295 1260.365 6.815 1260.905 ;
        RECT 2912.805 1260.905 2914.015 1261.995 ;
        RECT 2912.805 1260.365 2913.325 1260.905 ;
        RECT 6.295 1257.815 6.815 1258.355 ;
        RECT 5.605 1256.725 6.815 1257.815 ;
        RECT 2906.365 1256.725 2906.655 1257.890 ;
        RECT 2912.805 1257.815 2913.325 1258.355 ;
        RECT 2912.805 1256.725 2914.015 1257.815 ;
        RECT 5.520 1256.555 6.900 1256.725 ;
        RECT 2906.300 1256.555 2906.740 1256.725 ;
        RECT 2912.720 1256.555 2914.100 1256.725 ;
        RECT 5.605 1255.465 6.815 1256.555 ;
        RECT 6.295 1254.925 6.815 1255.465 ;
        RECT 2912.805 1255.465 2914.015 1256.555 ;
        RECT 2912.805 1254.925 2913.325 1255.465 ;
        RECT 6.295 1252.375 6.815 1252.915 ;
        RECT 5.605 1251.285 6.815 1252.375 ;
        RECT 2906.365 1251.285 2906.655 1252.450 ;
        RECT 2912.805 1252.375 2913.325 1252.915 ;
        RECT 2912.805 1251.285 2914.015 1252.375 ;
        RECT 5.520 1251.115 6.900 1251.285 ;
        RECT 2906.300 1251.115 2906.740 1251.285 ;
        RECT 2912.720 1251.115 2914.100 1251.285 ;
        RECT 5.605 1250.025 6.815 1251.115 ;
        RECT 6.295 1249.485 6.815 1250.025 ;
        RECT 2912.805 1250.025 2914.015 1251.115 ;
        RECT 2912.805 1249.485 2913.325 1250.025 ;
        RECT 6.295 1246.935 6.815 1247.475 ;
        RECT 5.605 1245.845 6.815 1246.935 ;
        RECT 2906.365 1245.845 2906.655 1247.010 ;
        RECT 2912.805 1246.935 2913.325 1247.475 ;
        RECT 2912.805 1245.845 2914.015 1246.935 ;
        RECT 5.520 1245.675 6.900 1245.845 ;
        RECT 2906.300 1245.675 2906.740 1245.845 ;
        RECT 2912.720 1245.675 2914.100 1245.845 ;
        RECT 5.605 1244.585 6.815 1245.675 ;
        RECT 6.295 1244.045 6.815 1244.585 ;
        RECT 2912.805 1244.585 2914.015 1245.675 ;
        RECT 2912.805 1244.045 2913.325 1244.585 ;
        RECT 6.295 1241.495 6.815 1242.035 ;
        RECT 5.605 1240.405 6.815 1241.495 ;
        RECT 2912.805 1241.495 2913.325 1242.035 ;
        RECT 2912.805 1240.405 2914.015 1241.495 ;
        RECT 5.520 1240.235 6.900 1240.405 ;
        RECT 2909.960 1240.235 2910.420 1240.405 ;
        RECT 2912.720 1240.235 2914.100 1240.405 ;
        RECT 5.605 1239.145 6.815 1240.235 ;
        RECT 6.295 1238.605 6.815 1239.145 ;
        RECT 2910.045 1239.070 2910.335 1240.235 ;
        RECT 2912.805 1239.145 2914.015 1240.235 ;
        RECT 2912.805 1238.605 2913.325 1239.145 ;
        RECT 6.295 1236.055 6.815 1236.595 ;
        RECT 5.605 1234.965 6.815 1236.055 ;
        RECT 2912.805 1236.055 2913.325 1236.595 ;
        RECT 2912.805 1234.965 2914.015 1236.055 ;
        RECT 5.520 1234.795 6.900 1234.965 ;
        RECT 2909.960 1234.795 2910.420 1234.965 ;
        RECT 2912.720 1234.795 2914.100 1234.965 ;
        RECT 5.605 1233.705 6.815 1234.795 ;
        RECT 6.295 1233.165 6.815 1233.705 ;
        RECT 2910.045 1233.630 2910.335 1234.795 ;
        RECT 2912.805 1233.705 2914.015 1234.795 ;
        RECT 2912.805 1233.165 2913.325 1233.705 ;
        RECT 6.295 1230.615 6.815 1231.155 ;
        RECT 5.605 1229.525 6.815 1230.615 ;
        RECT 2912.805 1230.615 2913.325 1231.155 ;
        RECT 2912.805 1229.525 2914.015 1230.615 ;
        RECT 5.520 1229.355 6.900 1229.525 ;
        RECT 2909.960 1229.355 2910.420 1229.525 ;
        RECT 2912.720 1229.355 2914.100 1229.525 ;
        RECT 5.605 1228.265 6.815 1229.355 ;
        RECT 6.295 1227.725 6.815 1228.265 ;
        RECT 2910.045 1228.190 2910.335 1229.355 ;
        RECT 2912.805 1228.265 2914.015 1229.355 ;
        RECT 2912.805 1227.725 2913.325 1228.265 ;
        RECT 6.295 1225.175 6.815 1225.715 ;
        RECT 5.605 1224.085 6.815 1225.175 ;
        RECT 2912.805 1225.175 2913.325 1225.715 ;
        RECT 2912.805 1224.085 2914.015 1225.175 ;
        RECT 5.520 1223.915 6.900 1224.085 ;
        RECT 2909.960 1223.915 2910.420 1224.085 ;
        RECT 2912.720 1223.915 2914.100 1224.085 ;
        RECT 5.605 1222.825 6.815 1223.915 ;
        RECT 6.295 1222.285 6.815 1222.825 ;
        RECT 2910.045 1222.750 2910.335 1223.915 ;
        RECT 2912.805 1222.825 2914.015 1223.915 ;
        RECT 2912.805 1222.285 2913.325 1222.825 ;
        RECT 6.295 1219.735 6.815 1220.275 ;
        RECT 5.605 1218.645 6.815 1219.735 ;
        RECT 2912.805 1219.735 2913.325 1220.275 ;
        RECT 2912.805 1218.645 2914.015 1219.735 ;
        RECT 5.520 1218.475 6.900 1218.645 ;
        RECT 8.740 1218.475 10.120 1218.645 ;
        RECT 2909.960 1218.475 2910.420 1218.645 ;
        RECT 2912.720 1218.475 2914.100 1218.645 ;
        RECT 5.605 1217.385 6.815 1218.475 ;
        RECT 9.015 1217.750 9.345 1218.475 ;
        RECT 6.295 1216.845 6.815 1217.385 ;
        RECT 2910.045 1217.310 2910.335 1218.475 ;
        RECT 2912.805 1217.385 2914.015 1218.475 ;
        RECT 2912.805 1216.845 2913.325 1217.385 ;
        RECT 6.295 1214.295 6.815 1214.835 ;
        RECT 5.605 1213.205 6.815 1214.295 ;
        RECT 2912.805 1214.295 2913.325 1214.835 ;
        RECT 2912.805 1213.205 2914.015 1214.295 ;
        RECT 5.520 1213.035 6.900 1213.205 ;
        RECT 2909.960 1213.035 2910.420 1213.205 ;
        RECT 2912.720 1213.035 2914.100 1213.205 ;
        RECT 5.605 1211.945 6.815 1213.035 ;
        RECT 6.295 1211.405 6.815 1211.945 ;
        RECT 2910.045 1211.870 2910.335 1213.035 ;
        RECT 2912.805 1211.945 2914.015 1213.035 ;
        RECT 2912.805 1211.405 2913.325 1211.945 ;
        RECT 6.295 1208.855 6.815 1209.395 ;
        RECT 5.605 1207.765 6.815 1208.855 ;
        RECT 2912.805 1208.855 2913.325 1209.395 ;
        RECT 2912.805 1207.765 2914.015 1208.855 ;
        RECT 5.520 1207.595 6.900 1207.765 ;
        RECT 2909.960 1207.595 2910.420 1207.765 ;
        RECT 2912.720 1207.595 2914.100 1207.765 ;
        RECT 5.605 1206.505 6.815 1207.595 ;
        RECT 6.295 1205.965 6.815 1206.505 ;
        RECT 2910.045 1206.430 2910.335 1207.595 ;
        RECT 2912.805 1206.505 2914.015 1207.595 ;
        RECT 2912.805 1205.965 2913.325 1206.505 ;
        RECT 6.295 1203.415 6.815 1203.955 ;
        RECT 5.605 1202.325 6.815 1203.415 ;
        RECT 2912.805 1203.415 2913.325 1203.955 ;
        RECT 2912.805 1202.325 2914.015 1203.415 ;
        RECT 5.520 1202.155 6.900 1202.325 ;
        RECT 2909.960 1202.155 2910.420 1202.325 ;
        RECT 2912.720 1202.155 2914.100 1202.325 ;
        RECT 5.605 1201.065 6.815 1202.155 ;
        RECT 6.295 1200.525 6.815 1201.065 ;
        RECT 2910.045 1200.990 2910.335 1202.155 ;
        RECT 2912.805 1201.065 2914.015 1202.155 ;
        RECT 2912.805 1200.525 2913.325 1201.065 ;
        RECT 6.295 1197.975 6.815 1198.515 ;
        RECT 5.605 1196.885 6.815 1197.975 ;
        RECT 2912.805 1197.975 2913.325 1198.515 ;
        RECT 2912.805 1196.885 2914.015 1197.975 ;
        RECT 5.520 1196.715 6.900 1196.885 ;
        RECT 2909.960 1196.715 2910.420 1196.885 ;
        RECT 2912.720 1196.715 2914.100 1196.885 ;
        RECT 5.605 1195.625 6.815 1196.715 ;
        RECT 6.295 1195.085 6.815 1195.625 ;
        RECT 2910.045 1195.550 2910.335 1196.715 ;
        RECT 2912.805 1195.625 2914.015 1196.715 ;
        RECT 2912.805 1195.085 2913.325 1195.625 ;
        RECT 6.295 1192.535 6.815 1193.075 ;
        RECT 5.605 1191.445 6.815 1192.535 ;
        RECT 2912.805 1192.535 2913.325 1193.075 ;
        RECT 2912.805 1191.445 2914.015 1192.535 ;
        RECT 5.520 1191.275 6.900 1191.445 ;
        RECT 2909.960 1191.275 2910.420 1191.445 ;
        RECT 2912.720 1191.275 2914.100 1191.445 ;
        RECT 5.605 1190.185 6.815 1191.275 ;
        RECT 6.295 1189.645 6.815 1190.185 ;
        RECT 2910.045 1190.110 2910.335 1191.275 ;
        RECT 2912.805 1190.185 2914.015 1191.275 ;
        RECT 2912.805 1189.645 2913.325 1190.185 ;
        RECT 6.295 1187.095 6.815 1187.635 ;
        RECT 5.605 1186.005 6.815 1187.095 ;
        RECT 2912.805 1187.095 2913.325 1187.635 ;
        RECT 2912.805 1186.005 2914.015 1187.095 ;
        RECT 5.520 1185.835 6.900 1186.005 ;
        RECT 2909.960 1185.835 2910.420 1186.005 ;
        RECT 2912.720 1185.835 2914.100 1186.005 ;
        RECT 5.605 1184.745 6.815 1185.835 ;
        RECT 6.295 1184.205 6.815 1184.745 ;
        RECT 2910.045 1184.670 2910.335 1185.835 ;
        RECT 2912.805 1184.745 2914.015 1185.835 ;
        RECT 2912.805 1184.205 2913.325 1184.745 ;
        RECT 6.295 1181.655 6.815 1182.195 ;
        RECT 5.605 1180.565 6.815 1181.655 ;
        RECT 2912.805 1181.655 2913.325 1182.195 ;
        RECT 2912.805 1180.565 2914.015 1181.655 ;
        RECT 5.520 1180.395 6.900 1180.565 ;
        RECT 2909.960 1180.395 2910.420 1180.565 ;
        RECT 2912.720 1180.395 2914.100 1180.565 ;
        RECT 5.605 1179.305 6.815 1180.395 ;
        RECT 6.295 1178.765 6.815 1179.305 ;
        RECT 2910.045 1179.230 2910.335 1180.395 ;
        RECT 2912.805 1179.305 2914.015 1180.395 ;
        RECT 2912.805 1178.765 2913.325 1179.305 ;
        RECT 6.295 1176.215 6.815 1176.755 ;
        RECT 5.605 1175.125 6.815 1176.215 ;
        RECT 2912.805 1176.215 2913.325 1176.755 ;
        RECT 2912.805 1175.125 2914.015 1176.215 ;
        RECT 5.520 1174.955 6.900 1175.125 ;
        RECT 2909.960 1174.955 2910.420 1175.125 ;
        RECT 2912.720 1174.955 2914.100 1175.125 ;
        RECT 5.605 1173.865 6.815 1174.955 ;
        RECT 6.295 1173.325 6.815 1173.865 ;
        RECT 2910.045 1173.790 2910.335 1174.955 ;
        RECT 2912.805 1173.865 2914.015 1174.955 ;
        RECT 2912.805 1173.325 2913.325 1173.865 ;
        RECT 6.295 1170.775 6.815 1171.315 ;
        RECT 5.605 1169.685 6.815 1170.775 ;
        RECT 2912.805 1170.775 2913.325 1171.315 ;
        RECT 2912.805 1169.685 2914.015 1170.775 ;
        RECT 5.520 1169.515 6.900 1169.685 ;
        RECT 2909.960 1169.515 2910.420 1169.685 ;
        RECT 2912.720 1169.515 2914.100 1169.685 ;
        RECT 5.605 1168.425 6.815 1169.515 ;
        RECT 6.295 1167.885 6.815 1168.425 ;
        RECT 2910.045 1168.350 2910.335 1169.515 ;
        RECT 2912.805 1168.425 2914.015 1169.515 ;
        RECT 2912.805 1167.885 2913.325 1168.425 ;
        RECT 6.295 1165.335 6.815 1165.875 ;
        RECT 5.605 1164.245 6.815 1165.335 ;
        RECT 2912.805 1165.335 2913.325 1165.875 ;
        RECT 2912.805 1164.245 2914.015 1165.335 ;
        RECT 5.520 1164.075 6.900 1164.245 ;
        RECT 2909.960 1164.075 2910.420 1164.245 ;
        RECT 2912.720 1164.075 2914.100 1164.245 ;
        RECT 5.605 1162.985 6.815 1164.075 ;
        RECT 6.295 1162.445 6.815 1162.985 ;
        RECT 2910.045 1162.910 2910.335 1164.075 ;
        RECT 2912.805 1162.985 2914.015 1164.075 ;
        RECT 2912.805 1162.445 2913.325 1162.985 ;
        RECT 6.295 1159.895 6.815 1160.435 ;
        RECT 5.605 1158.805 6.815 1159.895 ;
        RECT 2912.805 1159.895 2913.325 1160.435 ;
        RECT 2912.805 1158.805 2914.015 1159.895 ;
        RECT 5.520 1158.635 6.900 1158.805 ;
        RECT 2909.960 1158.635 2910.420 1158.805 ;
        RECT 2912.720 1158.635 2914.100 1158.805 ;
        RECT 5.605 1157.545 6.815 1158.635 ;
        RECT 6.295 1157.005 6.815 1157.545 ;
        RECT 2910.045 1157.470 2910.335 1158.635 ;
        RECT 2912.805 1157.545 2914.015 1158.635 ;
        RECT 2912.805 1157.005 2913.325 1157.545 ;
        RECT 6.295 1154.455 6.815 1154.995 ;
        RECT 5.605 1153.365 6.815 1154.455 ;
        RECT 2912.805 1154.455 2913.325 1154.995 ;
        RECT 2912.805 1153.365 2914.015 1154.455 ;
        RECT 5.520 1153.195 6.900 1153.365 ;
        RECT 2909.960 1153.195 2910.420 1153.365 ;
        RECT 2912.720 1153.195 2914.100 1153.365 ;
        RECT 5.605 1152.105 6.815 1153.195 ;
        RECT 6.295 1151.565 6.815 1152.105 ;
        RECT 2910.045 1152.030 2910.335 1153.195 ;
        RECT 2912.805 1152.105 2914.015 1153.195 ;
        RECT 2912.805 1151.565 2913.325 1152.105 ;
        RECT 6.295 1149.015 6.815 1149.555 ;
        RECT 5.605 1147.925 6.815 1149.015 ;
        RECT 2912.805 1149.015 2913.325 1149.555 ;
        RECT 2912.805 1147.925 2914.015 1149.015 ;
        RECT 5.520 1147.755 6.900 1147.925 ;
        RECT 2909.960 1147.755 2910.420 1147.925 ;
        RECT 2912.720 1147.755 2914.100 1147.925 ;
        RECT 5.605 1146.665 6.815 1147.755 ;
        RECT 6.295 1146.125 6.815 1146.665 ;
        RECT 2910.045 1146.590 2910.335 1147.755 ;
        RECT 2912.805 1146.665 2914.015 1147.755 ;
        RECT 2912.805 1146.125 2913.325 1146.665 ;
        RECT 6.295 1143.575 6.815 1144.115 ;
        RECT 5.605 1142.485 6.815 1143.575 ;
        RECT 2912.805 1143.575 2913.325 1144.115 ;
        RECT 2912.805 1142.485 2914.015 1143.575 ;
        RECT 5.520 1142.315 6.900 1142.485 ;
        RECT 2909.960 1142.315 2910.420 1142.485 ;
        RECT 2912.720 1142.315 2914.100 1142.485 ;
        RECT 5.605 1141.225 6.815 1142.315 ;
        RECT 6.295 1140.685 6.815 1141.225 ;
        RECT 2910.045 1141.150 2910.335 1142.315 ;
        RECT 2912.805 1141.225 2914.015 1142.315 ;
        RECT 2912.805 1140.685 2913.325 1141.225 ;
        RECT 6.295 1138.135 6.815 1138.675 ;
        RECT 5.605 1137.045 6.815 1138.135 ;
        RECT 2912.805 1138.135 2913.325 1138.675 ;
        RECT 2912.805 1137.045 2914.015 1138.135 ;
        RECT 5.520 1136.875 6.900 1137.045 ;
        RECT 2909.960 1136.875 2910.420 1137.045 ;
        RECT 2912.720 1136.875 2914.100 1137.045 ;
        RECT 5.605 1135.785 6.815 1136.875 ;
        RECT 6.295 1135.245 6.815 1135.785 ;
        RECT 2910.045 1135.710 2910.335 1136.875 ;
        RECT 2912.805 1135.785 2914.015 1136.875 ;
        RECT 2912.805 1135.245 2913.325 1135.785 ;
        RECT 6.295 1132.695 6.815 1133.235 ;
        RECT 5.605 1131.605 6.815 1132.695 ;
        RECT 2912.805 1132.695 2913.325 1133.235 ;
        RECT 2912.805 1131.605 2914.015 1132.695 ;
        RECT 5.520 1131.435 6.900 1131.605 ;
        RECT 2909.960 1131.435 2910.420 1131.605 ;
        RECT 2912.720 1131.435 2914.100 1131.605 ;
        RECT 5.605 1130.345 6.815 1131.435 ;
        RECT 6.295 1129.805 6.815 1130.345 ;
        RECT 2910.045 1130.270 2910.335 1131.435 ;
        RECT 2912.805 1130.345 2914.015 1131.435 ;
        RECT 2912.805 1129.805 2913.325 1130.345 ;
        RECT 6.295 1127.255 6.815 1127.795 ;
        RECT 5.605 1126.165 6.815 1127.255 ;
        RECT 2912.805 1127.255 2913.325 1127.795 ;
        RECT 2912.805 1126.165 2914.015 1127.255 ;
        RECT 5.520 1125.995 6.900 1126.165 ;
        RECT 2909.960 1125.995 2910.420 1126.165 ;
        RECT 2912.720 1125.995 2914.100 1126.165 ;
        RECT 5.605 1124.905 6.815 1125.995 ;
        RECT 6.295 1124.365 6.815 1124.905 ;
        RECT 2910.045 1124.830 2910.335 1125.995 ;
        RECT 2912.805 1124.905 2914.015 1125.995 ;
        RECT 2912.805 1124.365 2913.325 1124.905 ;
        RECT 6.295 1121.815 6.815 1122.355 ;
        RECT 5.605 1120.725 6.815 1121.815 ;
        RECT 2912.805 1121.815 2913.325 1122.355 ;
        RECT 2912.805 1120.725 2914.015 1121.815 ;
        RECT 5.520 1120.555 6.900 1120.725 ;
        RECT 2909.960 1120.555 2910.420 1120.725 ;
        RECT 2912.720 1120.555 2914.100 1120.725 ;
        RECT 5.605 1119.465 6.815 1120.555 ;
        RECT 6.295 1118.925 6.815 1119.465 ;
        RECT 2910.045 1119.390 2910.335 1120.555 ;
        RECT 2912.805 1119.465 2914.015 1120.555 ;
        RECT 2912.805 1118.925 2913.325 1119.465 ;
        RECT 6.295 1116.375 6.815 1116.915 ;
        RECT 5.605 1115.285 6.815 1116.375 ;
        RECT 2912.805 1116.375 2913.325 1116.915 ;
        RECT 2912.805 1115.285 2914.015 1116.375 ;
        RECT 5.520 1115.115 6.900 1115.285 ;
        RECT 2909.960 1115.115 2910.420 1115.285 ;
        RECT 2912.720 1115.115 2914.100 1115.285 ;
        RECT 5.605 1114.025 6.815 1115.115 ;
        RECT 6.295 1113.485 6.815 1114.025 ;
        RECT 2910.045 1113.950 2910.335 1115.115 ;
        RECT 2912.805 1114.025 2914.015 1115.115 ;
        RECT 2912.805 1113.485 2913.325 1114.025 ;
        RECT 6.295 1110.935 6.815 1111.475 ;
        RECT 5.605 1109.845 6.815 1110.935 ;
        RECT 2912.805 1110.935 2913.325 1111.475 ;
        RECT 9.015 1109.845 9.345 1110.570 ;
        RECT 2912.805 1109.845 2914.015 1110.935 ;
        RECT 5.520 1109.675 6.900 1109.845 ;
        RECT 8.740 1109.675 10.120 1109.845 ;
        RECT 2909.960 1109.675 2910.420 1109.845 ;
        RECT 2912.720 1109.675 2914.100 1109.845 ;
        RECT 5.605 1108.585 6.815 1109.675 ;
        RECT 6.295 1108.045 6.815 1108.585 ;
        RECT 2910.045 1108.510 2910.335 1109.675 ;
        RECT 2912.805 1108.585 2914.015 1109.675 ;
        RECT 2912.805 1108.045 2913.325 1108.585 ;
        RECT 6.295 1105.495 6.815 1106.035 ;
        RECT 5.605 1104.405 6.815 1105.495 ;
        RECT 2912.805 1105.495 2913.325 1106.035 ;
        RECT 2912.805 1104.405 2914.015 1105.495 ;
        RECT 5.520 1104.235 6.900 1104.405 ;
        RECT 2909.960 1104.235 2910.420 1104.405 ;
        RECT 2912.720 1104.235 2914.100 1104.405 ;
        RECT 5.605 1103.145 6.815 1104.235 ;
        RECT 6.295 1102.605 6.815 1103.145 ;
        RECT 2910.045 1103.070 2910.335 1104.235 ;
        RECT 2912.805 1103.145 2914.015 1104.235 ;
        RECT 2912.805 1102.605 2913.325 1103.145 ;
        RECT 6.295 1100.055 6.815 1100.595 ;
        RECT 5.605 1098.965 6.815 1100.055 ;
        RECT 2912.805 1100.055 2913.325 1100.595 ;
        RECT 2912.805 1098.965 2914.015 1100.055 ;
        RECT 5.520 1098.795 6.900 1098.965 ;
        RECT 2909.960 1098.795 2910.420 1098.965 ;
        RECT 2912.720 1098.795 2914.100 1098.965 ;
        RECT 5.605 1097.705 6.815 1098.795 ;
        RECT 6.295 1097.165 6.815 1097.705 ;
        RECT 2910.045 1097.630 2910.335 1098.795 ;
        RECT 2912.805 1097.705 2914.015 1098.795 ;
        RECT 2912.805 1097.165 2913.325 1097.705 ;
        RECT 6.295 1094.615 6.815 1095.155 ;
        RECT 5.605 1093.525 6.815 1094.615 ;
        RECT 2912.805 1094.615 2913.325 1095.155 ;
        RECT 2912.805 1093.525 2914.015 1094.615 ;
        RECT 5.520 1093.355 6.900 1093.525 ;
        RECT 2909.960 1093.355 2910.420 1093.525 ;
        RECT 2912.720 1093.355 2914.100 1093.525 ;
        RECT 5.605 1092.265 6.815 1093.355 ;
        RECT 6.295 1091.725 6.815 1092.265 ;
        RECT 2910.045 1092.190 2910.335 1093.355 ;
        RECT 2912.805 1092.265 2914.015 1093.355 ;
        RECT 2912.805 1091.725 2913.325 1092.265 ;
        RECT 6.295 1089.175 6.815 1089.715 ;
        RECT 5.605 1088.085 6.815 1089.175 ;
        RECT 2912.805 1089.175 2913.325 1089.715 ;
        RECT 2912.805 1088.085 2914.015 1089.175 ;
        RECT 5.520 1087.915 6.900 1088.085 ;
        RECT 2909.960 1087.915 2910.420 1088.085 ;
        RECT 2912.720 1087.915 2914.100 1088.085 ;
        RECT 5.605 1086.825 6.815 1087.915 ;
        RECT 6.295 1086.285 6.815 1086.825 ;
        RECT 2910.045 1086.750 2910.335 1087.915 ;
        RECT 2912.805 1086.825 2914.015 1087.915 ;
        RECT 2912.805 1086.285 2913.325 1086.825 ;
        RECT 6.295 1083.735 6.815 1084.275 ;
        RECT 5.605 1082.645 6.815 1083.735 ;
        RECT 2912.805 1083.735 2913.325 1084.275 ;
        RECT 2912.805 1082.645 2914.015 1083.735 ;
        RECT 5.520 1082.475 6.900 1082.645 ;
        RECT 2909.960 1082.475 2910.420 1082.645 ;
        RECT 2912.720 1082.475 2914.100 1082.645 ;
        RECT 5.605 1081.385 6.815 1082.475 ;
        RECT 6.295 1080.845 6.815 1081.385 ;
        RECT 2910.045 1081.310 2910.335 1082.475 ;
        RECT 2912.805 1081.385 2914.015 1082.475 ;
        RECT 2912.805 1080.845 2913.325 1081.385 ;
        RECT 6.295 1078.295 6.815 1078.835 ;
        RECT 5.605 1077.205 6.815 1078.295 ;
        RECT 2912.805 1078.295 2913.325 1078.835 ;
        RECT 2912.805 1077.205 2914.015 1078.295 ;
        RECT 5.520 1077.035 6.900 1077.205 ;
        RECT 2909.960 1077.035 2910.420 1077.205 ;
        RECT 2912.720 1077.035 2914.100 1077.205 ;
        RECT 5.605 1075.945 6.815 1077.035 ;
        RECT 6.295 1075.405 6.815 1075.945 ;
        RECT 2910.045 1075.870 2910.335 1077.035 ;
        RECT 2912.805 1075.945 2914.015 1077.035 ;
        RECT 2912.805 1075.405 2913.325 1075.945 ;
        RECT 6.295 1072.855 6.815 1073.395 ;
        RECT 5.605 1071.765 6.815 1072.855 ;
        RECT 2912.805 1072.855 2913.325 1073.395 ;
        RECT 2912.805 1071.765 2914.015 1072.855 ;
        RECT 5.520 1071.595 6.900 1071.765 ;
        RECT 2909.960 1071.595 2910.420 1071.765 ;
        RECT 2912.720 1071.595 2914.100 1071.765 ;
        RECT 5.605 1070.505 6.815 1071.595 ;
        RECT 6.295 1069.965 6.815 1070.505 ;
        RECT 2910.045 1070.430 2910.335 1071.595 ;
        RECT 2912.805 1070.505 2914.015 1071.595 ;
        RECT 2912.805 1069.965 2913.325 1070.505 ;
        RECT 6.295 1067.415 6.815 1067.955 ;
        RECT 5.605 1066.325 6.815 1067.415 ;
        RECT 2912.805 1067.415 2913.325 1067.955 ;
        RECT 2912.805 1066.325 2914.015 1067.415 ;
        RECT 5.520 1066.155 6.900 1066.325 ;
        RECT 2909.960 1066.155 2910.420 1066.325 ;
        RECT 2912.720 1066.155 2914.100 1066.325 ;
        RECT 5.605 1065.065 6.815 1066.155 ;
        RECT 6.295 1064.525 6.815 1065.065 ;
        RECT 2910.045 1064.990 2910.335 1066.155 ;
        RECT 2912.805 1065.065 2914.015 1066.155 ;
        RECT 2912.805 1064.525 2913.325 1065.065 ;
        RECT 6.295 1061.975 6.815 1062.515 ;
        RECT 5.605 1060.885 6.815 1061.975 ;
        RECT 2912.805 1061.975 2913.325 1062.515 ;
        RECT 2912.805 1060.885 2914.015 1061.975 ;
        RECT 5.520 1060.715 6.900 1060.885 ;
        RECT 2909.960 1060.715 2910.420 1060.885 ;
        RECT 2912.720 1060.715 2914.100 1060.885 ;
        RECT 5.605 1059.625 6.815 1060.715 ;
        RECT 6.295 1059.085 6.815 1059.625 ;
        RECT 2910.045 1059.550 2910.335 1060.715 ;
        RECT 2912.805 1059.625 2914.015 1060.715 ;
        RECT 2912.805 1059.085 2913.325 1059.625 ;
        RECT 6.295 1056.535 6.815 1057.075 ;
        RECT 5.605 1055.445 6.815 1056.535 ;
        RECT 2912.805 1056.535 2913.325 1057.075 ;
        RECT 2912.805 1055.445 2914.015 1056.535 ;
        RECT 5.520 1055.275 6.900 1055.445 ;
        RECT 2909.960 1055.275 2910.420 1055.445 ;
        RECT 2912.720 1055.275 2914.100 1055.445 ;
        RECT 5.605 1054.185 6.815 1055.275 ;
        RECT 6.295 1053.645 6.815 1054.185 ;
        RECT 2910.045 1054.110 2910.335 1055.275 ;
        RECT 2912.805 1054.185 2914.015 1055.275 ;
        RECT 2912.805 1053.645 2913.325 1054.185 ;
        RECT 6.295 1051.095 6.815 1051.635 ;
        RECT 5.605 1050.005 6.815 1051.095 ;
        RECT 2912.805 1051.095 2913.325 1051.635 ;
        RECT 2912.805 1050.005 2914.015 1051.095 ;
        RECT 5.520 1049.835 6.900 1050.005 ;
        RECT 2909.960 1049.835 2910.420 1050.005 ;
        RECT 2912.720 1049.835 2914.100 1050.005 ;
        RECT 5.605 1048.745 6.815 1049.835 ;
        RECT 6.295 1048.205 6.815 1048.745 ;
        RECT 2910.045 1048.670 2910.335 1049.835 ;
        RECT 2912.805 1048.745 2914.015 1049.835 ;
        RECT 2912.805 1048.205 2913.325 1048.745 ;
        RECT 6.295 1045.655 6.815 1046.195 ;
        RECT 5.605 1044.565 6.815 1045.655 ;
        RECT 2912.805 1045.655 2913.325 1046.195 ;
        RECT 2912.805 1044.565 2914.015 1045.655 ;
        RECT 5.520 1044.395 6.900 1044.565 ;
        RECT 2909.960 1044.395 2910.420 1044.565 ;
        RECT 2912.720 1044.395 2914.100 1044.565 ;
        RECT 5.605 1043.305 6.815 1044.395 ;
        RECT 6.295 1042.765 6.815 1043.305 ;
        RECT 2910.045 1043.230 2910.335 1044.395 ;
        RECT 2912.805 1043.305 2914.015 1044.395 ;
        RECT 2912.805 1042.765 2913.325 1043.305 ;
        RECT 6.295 1040.215 6.815 1040.755 ;
        RECT 5.605 1039.125 6.815 1040.215 ;
        RECT 2912.805 1040.215 2913.325 1040.755 ;
        RECT 2912.805 1039.125 2914.015 1040.215 ;
        RECT 5.520 1038.955 6.900 1039.125 ;
        RECT 2909.960 1038.955 2910.420 1039.125 ;
        RECT 2912.720 1038.955 2914.100 1039.125 ;
        RECT 5.605 1037.865 6.815 1038.955 ;
        RECT 6.295 1037.325 6.815 1037.865 ;
        RECT 2910.045 1037.790 2910.335 1038.955 ;
        RECT 2912.805 1037.865 2914.015 1038.955 ;
        RECT 2912.805 1037.325 2913.325 1037.865 ;
        RECT 6.295 1034.775 6.815 1035.315 ;
        RECT 5.605 1033.685 6.815 1034.775 ;
        RECT 2912.805 1034.775 2913.325 1035.315 ;
        RECT 9.015 1033.685 9.345 1034.410 ;
        RECT 2912.805 1033.685 2914.015 1034.775 ;
        RECT 5.520 1033.515 6.900 1033.685 ;
        RECT 8.740 1033.515 10.120 1033.685 ;
        RECT 2909.960 1033.515 2910.420 1033.685 ;
        RECT 2912.720 1033.515 2914.100 1033.685 ;
        RECT 5.605 1032.425 6.815 1033.515 ;
        RECT 6.295 1031.885 6.815 1032.425 ;
        RECT 2910.045 1032.350 2910.335 1033.515 ;
        RECT 2912.805 1032.425 2914.015 1033.515 ;
        RECT 2912.805 1031.885 2913.325 1032.425 ;
        RECT 6.295 1029.335 6.815 1029.875 ;
        RECT 5.605 1028.245 6.815 1029.335 ;
        RECT 2912.805 1029.335 2913.325 1029.875 ;
        RECT 2912.805 1028.245 2914.015 1029.335 ;
        RECT 5.520 1028.075 6.900 1028.245 ;
        RECT 2909.960 1028.075 2910.420 1028.245 ;
        RECT 2912.720 1028.075 2914.100 1028.245 ;
        RECT 5.605 1026.985 6.815 1028.075 ;
        RECT 6.295 1026.445 6.815 1026.985 ;
        RECT 2910.045 1026.910 2910.335 1028.075 ;
        RECT 2912.805 1026.985 2914.015 1028.075 ;
        RECT 2912.805 1026.445 2913.325 1026.985 ;
        RECT 6.295 1023.895 6.815 1024.435 ;
        RECT 5.605 1022.805 6.815 1023.895 ;
        RECT 2912.805 1023.895 2913.325 1024.435 ;
        RECT 2912.805 1022.805 2914.015 1023.895 ;
        RECT 5.520 1022.635 6.900 1022.805 ;
        RECT 2909.960 1022.635 2910.420 1022.805 ;
        RECT 2912.720 1022.635 2914.100 1022.805 ;
        RECT 5.605 1021.545 6.815 1022.635 ;
        RECT 6.295 1021.005 6.815 1021.545 ;
        RECT 2910.045 1021.470 2910.335 1022.635 ;
        RECT 2912.805 1021.545 2914.015 1022.635 ;
        RECT 2912.805 1021.005 2913.325 1021.545 ;
        RECT 6.295 1018.455 6.815 1018.995 ;
        RECT 5.605 1017.365 6.815 1018.455 ;
        RECT 2912.805 1018.455 2913.325 1018.995 ;
        RECT 2912.805 1017.365 2914.015 1018.455 ;
        RECT 5.520 1017.195 6.900 1017.365 ;
        RECT 2909.960 1017.195 2910.420 1017.365 ;
        RECT 2912.720 1017.195 2914.100 1017.365 ;
        RECT 5.605 1016.105 6.815 1017.195 ;
        RECT 6.295 1015.565 6.815 1016.105 ;
        RECT 2910.045 1016.030 2910.335 1017.195 ;
        RECT 2912.805 1016.105 2914.015 1017.195 ;
        RECT 2912.805 1015.565 2913.325 1016.105 ;
        RECT 6.295 1013.015 6.815 1013.555 ;
        RECT 5.605 1011.925 6.815 1013.015 ;
        RECT 2912.805 1013.015 2913.325 1013.555 ;
        RECT 2912.805 1011.925 2914.015 1013.015 ;
        RECT 5.520 1011.755 6.900 1011.925 ;
        RECT 2909.960 1011.755 2910.420 1011.925 ;
        RECT 2912.720 1011.755 2914.100 1011.925 ;
        RECT 5.605 1010.665 6.815 1011.755 ;
        RECT 6.295 1010.125 6.815 1010.665 ;
        RECT 2910.045 1010.590 2910.335 1011.755 ;
        RECT 2912.805 1010.665 2914.015 1011.755 ;
        RECT 2912.805 1010.125 2913.325 1010.665 ;
        RECT 6.295 1007.575 6.815 1008.115 ;
        RECT 5.605 1006.485 6.815 1007.575 ;
        RECT 2912.805 1007.575 2913.325 1008.115 ;
        RECT 2909.315 1006.485 2909.645 1007.210 ;
        RECT 2912.805 1006.485 2914.015 1007.575 ;
        RECT 5.520 1006.315 6.900 1006.485 ;
        RECT 2909.040 1006.315 2910.420 1006.485 ;
        RECT 2912.720 1006.315 2914.100 1006.485 ;
        RECT 5.605 1005.225 6.815 1006.315 ;
        RECT 6.295 1004.685 6.815 1005.225 ;
        RECT 2910.045 1005.150 2910.335 1006.315 ;
        RECT 2912.805 1005.225 2914.015 1006.315 ;
        RECT 2912.805 1004.685 2913.325 1005.225 ;
        RECT 6.295 1002.135 6.815 1002.675 ;
        RECT 5.605 1001.045 6.815 1002.135 ;
        RECT 2912.805 1002.135 2913.325 1002.675 ;
        RECT 2912.805 1001.045 2914.015 1002.135 ;
        RECT 5.520 1000.875 6.900 1001.045 ;
        RECT 2909.960 1000.875 2910.420 1001.045 ;
        RECT 2912.720 1000.875 2914.100 1001.045 ;
        RECT 5.605 999.785 6.815 1000.875 ;
        RECT 6.295 999.245 6.815 999.785 ;
        RECT 2910.045 999.710 2910.335 1000.875 ;
        RECT 2912.805 999.785 2914.015 1000.875 ;
        RECT 2912.805 999.245 2913.325 999.785 ;
        RECT 6.295 996.695 6.815 997.235 ;
        RECT 5.605 995.605 6.815 996.695 ;
        RECT 2912.805 996.695 2913.325 997.235 ;
        RECT 2909.315 995.605 2909.645 996.330 ;
        RECT 2912.805 995.605 2914.015 996.695 ;
        RECT 5.520 995.435 6.900 995.605 ;
        RECT 2909.040 995.435 2910.420 995.605 ;
        RECT 2912.720 995.435 2914.100 995.605 ;
        RECT 5.605 994.345 6.815 995.435 ;
        RECT 6.295 993.805 6.815 994.345 ;
        RECT 2910.045 994.270 2910.335 995.435 ;
        RECT 2912.805 994.345 2914.015 995.435 ;
        RECT 2912.805 993.805 2913.325 994.345 ;
        RECT 6.295 991.255 6.815 991.795 ;
        RECT 5.605 990.165 6.815 991.255 ;
        RECT 2912.805 991.255 2913.325 991.795 ;
        RECT 2912.805 990.165 2914.015 991.255 ;
        RECT 5.520 989.995 6.900 990.165 ;
        RECT 2909.960 989.995 2910.420 990.165 ;
        RECT 2912.720 989.995 2914.100 990.165 ;
        RECT 5.605 988.905 6.815 989.995 ;
        RECT 6.295 988.365 6.815 988.905 ;
        RECT 2910.045 988.830 2910.335 989.995 ;
        RECT 2912.805 988.905 2914.015 989.995 ;
        RECT 2912.805 988.365 2913.325 988.905 ;
        RECT 6.295 985.815 6.815 986.355 ;
        RECT 5.605 984.725 6.815 985.815 ;
        RECT 2912.805 985.815 2913.325 986.355 ;
        RECT 2912.805 984.725 2914.015 985.815 ;
        RECT 5.520 984.555 6.900 984.725 ;
        RECT 2909.960 984.555 2910.420 984.725 ;
        RECT 2912.720 984.555 2914.100 984.725 ;
        RECT 5.605 983.465 6.815 984.555 ;
        RECT 6.295 982.925 6.815 983.465 ;
        RECT 2910.045 983.390 2910.335 984.555 ;
        RECT 2912.805 983.465 2914.015 984.555 ;
        RECT 2912.805 982.925 2913.325 983.465 ;
        RECT 6.295 980.375 6.815 980.915 ;
        RECT 5.605 979.285 6.815 980.375 ;
        RECT 2912.805 980.375 2913.325 980.915 ;
        RECT 2912.805 979.285 2914.015 980.375 ;
        RECT 5.520 979.115 6.900 979.285 ;
        RECT 2909.960 979.115 2910.420 979.285 ;
        RECT 2912.720 979.115 2914.100 979.285 ;
        RECT 5.605 978.025 6.815 979.115 ;
        RECT 6.295 977.485 6.815 978.025 ;
        RECT 2910.045 977.950 2910.335 979.115 ;
        RECT 2912.805 978.025 2914.015 979.115 ;
        RECT 2912.805 977.485 2913.325 978.025 ;
        RECT 6.295 974.935 6.815 975.475 ;
        RECT 5.605 973.845 6.815 974.935 ;
        RECT 2912.805 974.935 2913.325 975.475 ;
        RECT 2912.805 973.845 2914.015 974.935 ;
        RECT 5.520 973.675 6.900 973.845 ;
        RECT 2909.960 973.675 2910.420 973.845 ;
        RECT 2912.720 973.675 2914.100 973.845 ;
        RECT 5.605 972.585 6.815 973.675 ;
        RECT 6.295 972.045 6.815 972.585 ;
        RECT 2910.045 972.510 2910.335 973.675 ;
        RECT 2912.805 972.585 2914.015 973.675 ;
        RECT 2912.805 972.045 2913.325 972.585 ;
        RECT 6.295 969.495 6.815 970.035 ;
        RECT 5.605 968.405 6.815 969.495 ;
        RECT 2912.805 969.495 2913.325 970.035 ;
        RECT 2912.805 968.405 2914.015 969.495 ;
        RECT 5.520 968.235 6.900 968.405 ;
        RECT 2909.960 968.235 2910.420 968.405 ;
        RECT 2912.720 968.235 2914.100 968.405 ;
        RECT 5.605 967.145 6.815 968.235 ;
        RECT 6.295 966.605 6.815 967.145 ;
        RECT 2910.045 967.070 2910.335 968.235 ;
        RECT 2912.805 967.145 2914.015 968.235 ;
        RECT 2912.805 966.605 2913.325 967.145 ;
        RECT 6.295 964.055 6.815 964.595 ;
        RECT 5.605 962.965 6.815 964.055 ;
        RECT 2912.805 964.055 2913.325 964.595 ;
        RECT 2912.805 962.965 2914.015 964.055 ;
        RECT 5.520 962.795 6.900 962.965 ;
        RECT 2909.960 962.795 2910.420 962.965 ;
        RECT 2912.720 962.795 2914.100 962.965 ;
        RECT 5.605 961.705 6.815 962.795 ;
        RECT 6.295 961.165 6.815 961.705 ;
        RECT 2910.045 961.630 2910.335 962.795 ;
        RECT 2912.805 961.705 2914.015 962.795 ;
        RECT 2912.805 961.165 2913.325 961.705 ;
        RECT 6.295 958.615 6.815 959.155 ;
        RECT 5.605 957.525 6.815 958.615 ;
        RECT 2912.805 958.615 2913.325 959.155 ;
        RECT 2912.805 957.525 2914.015 958.615 ;
        RECT 5.520 957.355 6.900 957.525 ;
        RECT 2909.960 957.355 2910.420 957.525 ;
        RECT 2912.720 957.355 2914.100 957.525 ;
        RECT 5.605 956.265 6.815 957.355 ;
        RECT 6.295 955.725 6.815 956.265 ;
        RECT 2910.045 956.190 2910.335 957.355 ;
        RECT 2912.805 956.265 2914.015 957.355 ;
        RECT 2912.805 955.725 2913.325 956.265 ;
        RECT 6.295 953.175 6.815 953.715 ;
        RECT 5.605 952.085 6.815 953.175 ;
        RECT 2912.805 953.175 2913.325 953.715 ;
        RECT 2912.805 952.085 2914.015 953.175 ;
        RECT 5.520 951.915 6.900 952.085 ;
        RECT 2909.960 951.915 2910.420 952.085 ;
        RECT 2912.720 951.915 2914.100 952.085 ;
        RECT 5.605 950.825 6.815 951.915 ;
        RECT 6.295 950.285 6.815 950.825 ;
        RECT 2910.045 950.750 2910.335 951.915 ;
        RECT 2912.805 950.825 2914.015 951.915 ;
        RECT 2912.805 950.285 2913.325 950.825 ;
        RECT 6.295 947.735 6.815 948.275 ;
        RECT 5.605 946.645 6.815 947.735 ;
        RECT 2912.805 947.735 2913.325 948.275 ;
        RECT 2912.805 946.645 2914.015 947.735 ;
        RECT 5.520 946.475 6.900 946.645 ;
        RECT 2909.960 946.475 2910.420 946.645 ;
        RECT 2912.720 946.475 2914.100 946.645 ;
        RECT 5.605 945.385 6.815 946.475 ;
        RECT 6.295 944.845 6.815 945.385 ;
        RECT 2910.045 945.310 2910.335 946.475 ;
        RECT 2912.805 945.385 2914.015 946.475 ;
        RECT 2912.805 944.845 2913.325 945.385 ;
        RECT 6.295 942.295 6.815 942.835 ;
        RECT 5.605 941.205 6.815 942.295 ;
        RECT 2912.805 942.295 2913.325 942.835 ;
        RECT 2912.805 941.205 2914.015 942.295 ;
        RECT 5.520 941.035 6.900 941.205 ;
        RECT 2909.960 941.035 2910.420 941.205 ;
        RECT 2912.720 941.035 2914.100 941.205 ;
        RECT 5.605 939.945 6.815 941.035 ;
        RECT 6.295 939.405 6.815 939.945 ;
        RECT 2910.045 939.870 2910.335 941.035 ;
        RECT 2912.805 939.945 2914.015 941.035 ;
        RECT 2912.805 939.405 2913.325 939.945 ;
        RECT 6.295 936.855 6.815 937.395 ;
        RECT 5.605 935.765 6.815 936.855 ;
        RECT 2912.805 936.855 2913.325 937.395 ;
        RECT 2912.805 935.765 2914.015 936.855 ;
        RECT 5.520 935.595 6.900 935.765 ;
        RECT 2909.960 935.595 2910.420 935.765 ;
        RECT 2912.720 935.595 2914.100 935.765 ;
        RECT 5.605 934.505 6.815 935.595 ;
        RECT 6.295 933.965 6.815 934.505 ;
        RECT 2910.045 934.430 2910.335 935.595 ;
        RECT 2912.805 934.505 2914.015 935.595 ;
        RECT 2912.805 933.965 2913.325 934.505 ;
        RECT 6.295 931.415 6.815 931.955 ;
        RECT 5.605 930.325 6.815 931.415 ;
        RECT 2912.805 931.415 2913.325 931.955 ;
        RECT 2912.805 930.325 2914.015 931.415 ;
        RECT 5.520 930.155 6.900 930.325 ;
        RECT 2909.960 930.155 2910.420 930.325 ;
        RECT 2912.720 930.155 2914.100 930.325 ;
        RECT 5.605 929.065 6.815 930.155 ;
        RECT 6.295 928.525 6.815 929.065 ;
        RECT 2910.045 928.990 2910.335 930.155 ;
        RECT 2912.805 929.065 2914.015 930.155 ;
        RECT 2912.805 928.525 2913.325 929.065 ;
        RECT 6.295 925.975 6.815 926.515 ;
        RECT 5.605 924.885 6.815 925.975 ;
        RECT 2912.805 925.975 2913.325 926.515 ;
        RECT 2912.805 924.885 2914.015 925.975 ;
        RECT 5.520 924.715 6.900 924.885 ;
        RECT 2909.960 924.715 2910.420 924.885 ;
        RECT 2912.720 924.715 2914.100 924.885 ;
        RECT 5.605 923.625 6.815 924.715 ;
        RECT 6.295 923.085 6.815 923.625 ;
        RECT 2910.045 923.550 2910.335 924.715 ;
        RECT 2912.805 923.625 2914.015 924.715 ;
        RECT 2912.805 923.085 2913.325 923.625 ;
        RECT 6.295 920.535 6.815 921.075 ;
        RECT 5.605 919.445 6.815 920.535 ;
        RECT 2912.805 920.535 2913.325 921.075 ;
        RECT 2912.805 919.445 2914.015 920.535 ;
        RECT 5.520 919.275 6.900 919.445 ;
        RECT 2909.960 919.275 2910.420 919.445 ;
        RECT 2912.720 919.275 2914.100 919.445 ;
        RECT 5.605 918.185 6.815 919.275 ;
        RECT 6.295 917.645 6.815 918.185 ;
        RECT 2910.045 918.110 2910.335 919.275 ;
        RECT 2912.805 918.185 2914.015 919.275 ;
        RECT 2912.805 917.645 2913.325 918.185 ;
        RECT 6.295 915.095 6.815 915.635 ;
        RECT 5.605 914.005 6.815 915.095 ;
        RECT 2912.805 915.095 2913.325 915.635 ;
        RECT 2912.805 914.005 2914.015 915.095 ;
        RECT 5.520 913.835 6.900 914.005 ;
        RECT 2909.960 913.835 2910.420 914.005 ;
        RECT 2912.720 913.835 2914.100 914.005 ;
        RECT 5.605 912.745 6.815 913.835 ;
        RECT 6.295 912.205 6.815 912.745 ;
        RECT 2910.045 912.670 2910.335 913.835 ;
        RECT 2912.805 912.745 2914.015 913.835 ;
        RECT 2912.805 912.205 2913.325 912.745 ;
        RECT 6.295 909.655 6.815 910.195 ;
        RECT 5.605 908.565 6.815 909.655 ;
        RECT 2912.805 909.655 2913.325 910.195 ;
        RECT 2912.805 908.565 2914.015 909.655 ;
        RECT 5.520 908.395 6.900 908.565 ;
        RECT 2909.960 908.395 2910.420 908.565 ;
        RECT 2912.720 908.395 2914.100 908.565 ;
        RECT 5.605 907.305 6.815 908.395 ;
        RECT 6.295 906.765 6.815 907.305 ;
        RECT 2910.045 907.230 2910.335 908.395 ;
        RECT 2912.805 907.305 2914.015 908.395 ;
        RECT 2912.805 906.765 2913.325 907.305 ;
        RECT 6.295 904.215 6.815 904.755 ;
        RECT 5.605 903.125 6.815 904.215 ;
        RECT 2912.805 904.215 2913.325 904.755 ;
        RECT 2912.805 903.125 2914.015 904.215 ;
        RECT 5.520 902.955 6.900 903.125 ;
        RECT 2909.960 902.955 2910.420 903.125 ;
        RECT 2912.720 902.955 2914.100 903.125 ;
        RECT 5.605 901.865 6.815 902.955 ;
        RECT 6.295 901.325 6.815 901.865 ;
        RECT 2910.045 901.790 2910.335 902.955 ;
        RECT 2912.805 901.865 2914.015 902.955 ;
        RECT 2912.805 901.325 2913.325 901.865 ;
        RECT 6.295 898.775 6.815 899.315 ;
        RECT 5.605 897.685 6.815 898.775 ;
        RECT 2912.805 898.775 2913.325 899.315 ;
        RECT 2912.805 897.685 2914.015 898.775 ;
        RECT 5.520 897.515 6.900 897.685 ;
        RECT 2909.960 897.515 2910.420 897.685 ;
        RECT 2912.720 897.515 2914.100 897.685 ;
        RECT 5.605 896.425 6.815 897.515 ;
        RECT 6.295 895.885 6.815 896.425 ;
        RECT 2910.045 896.350 2910.335 897.515 ;
        RECT 2912.805 896.425 2914.015 897.515 ;
        RECT 2912.805 895.885 2913.325 896.425 ;
        RECT 6.295 893.335 6.815 893.875 ;
        RECT 5.605 892.245 6.815 893.335 ;
        RECT 2912.805 893.335 2913.325 893.875 ;
        RECT 2912.805 892.245 2914.015 893.335 ;
        RECT 5.520 892.075 6.900 892.245 ;
        RECT 2909.960 892.075 2910.420 892.245 ;
        RECT 2912.720 892.075 2914.100 892.245 ;
        RECT 5.605 890.985 6.815 892.075 ;
        RECT 6.295 890.445 6.815 890.985 ;
        RECT 2910.045 890.910 2910.335 892.075 ;
        RECT 2912.805 890.985 2914.015 892.075 ;
        RECT 2912.805 890.445 2913.325 890.985 ;
        RECT 6.295 887.895 6.815 888.435 ;
        RECT 5.605 886.805 6.815 887.895 ;
        RECT 2912.805 887.895 2913.325 888.435 ;
        RECT 2912.805 886.805 2914.015 887.895 ;
        RECT 5.520 886.635 6.900 886.805 ;
        RECT 2909.960 886.635 2910.420 886.805 ;
        RECT 2912.720 886.635 2914.100 886.805 ;
        RECT 5.605 885.545 6.815 886.635 ;
        RECT 6.295 885.005 6.815 885.545 ;
        RECT 2910.045 885.470 2910.335 886.635 ;
        RECT 2912.805 885.545 2914.015 886.635 ;
        RECT 2912.805 885.005 2913.325 885.545 ;
        RECT 6.295 882.455 6.815 882.995 ;
        RECT 5.605 881.365 6.815 882.455 ;
        RECT 2912.805 882.455 2913.325 882.995 ;
        RECT 2912.805 881.365 2914.015 882.455 ;
        RECT 5.520 881.195 6.900 881.365 ;
        RECT 2909.960 881.195 2910.420 881.365 ;
        RECT 2912.720 881.195 2914.100 881.365 ;
        RECT 5.605 880.105 6.815 881.195 ;
        RECT 6.295 879.565 6.815 880.105 ;
        RECT 2910.045 880.030 2910.335 881.195 ;
        RECT 2912.805 880.105 2914.015 881.195 ;
        RECT 2912.805 879.565 2913.325 880.105 ;
        RECT 6.295 877.015 6.815 877.555 ;
        RECT 5.605 875.925 6.815 877.015 ;
        RECT 2912.805 877.015 2913.325 877.555 ;
        RECT 2912.805 875.925 2914.015 877.015 ;
        RECT 5.520 875.755 6.900 875.925 ;
        RECT 2909.960 875.755 2910.420 875.925 ;
        RECT 2912.720 875.755 2914.100 875.925 ;
        RECT 5.605 874.665 6.815 875.755 ;
        RECT 6.295 874.125 6.815 874.665 ;
        RECT 2910.045 874.590 2910.335 875.755 ;
        RECT 2912.805 874.665 2914.015 875.755 ;
        RECT 2912.805 874.125 2913.325 874.665 ;
        RECT 6.295 871.575 6.815 872.115 ;
        RECT 5.605 870.485 6.815 871.575 ;
        RECT 2912.805 871.575 2913.325 872.115 ;
        RECT 2912.805 870.485 2914.015 871.575 ;
        RECT 5.520 870.315 6.900 870.485 ;
        RECT 2909.960 870.315 2910.420 870.485 ;
        RECT 2912.720 870.315 2914.100 870.485 ;
        RECT 5.605 869.225 6.815 870.315 ;
        RECT 6.295 868.685 6.815 869.225 ;
        RECT 2910.045 869.150 2910.335 870.315 ;
        RECT 2912.805 869.225 2914.015 870.315 ;
        RECT 2912.805 868.685 2913.325 869.225 ;
        RECT 6.295 866.135 6.815 866.675 ;
        RECT 5.605 865.045 6.815 866.135 ;
        RECT 2912.805 866.135 2913.325 866.675 ;
        RECT 2912.805 865.045 2914.015 866.135 ;
        RECT 5.520 864.875 6.900 865.045 ;
        RECT 2909.960 864.875 2910.420 865.045 ;
        RECT 2912.720 864.875 2914.100 865.045 ;
        RECT 5.605 863.785 6.815 864.875 ;
        RECT 6.295 863.245 6.815 863.785 ;
        RECT 2910.045 863.710 2910.335 864.875 ;
        RECT 2912.805 863.785 2914.015 864.875 ;
        RECT 2912.805 863.245 2913.325 863.785 ;
        RECT 6.295 860.695 6.815 861.235 ;
        RECT 5.605 859.605 6.815 860.695 ;
        RECT 2912.805 860.695 2913.325 861.235 ;
        RECT 2912.805 859.605 2914.015 860.695 ;
        RECT 5.520 859.435 6.900 859.605 ;
        RECT 2909.960 859.435 2910.420 859.605 ;
        RECT 2912.720 859.435 2914.100 859.605 ;
        RECT 5.605 858.345 6.815 859.435 ;
        RECT 6.295 857.805 6.815 858.345 ;
        RECT 2910.045 858.270 2910.335 859.435 ;
        RECT 2912.805 858.345 2914.015 859.435 ;
        RECT 2912.805 857.805 2913.325 858.345 ;
        RECT 6.295 855.255 6.815 855.795 ;
        RECT 5.605 854.165 6.815 855.255 ;
        RECT 2912.805 855.255 2913.325 855.795 ;
        RECT 2912.805 854.165 2914.015 855.255 ;
        RECT 5.520 853.995 6.900 854.165 ;
        RECT 2909.960 853.995 2910.420 854.165 ;
        RECT 2912.720 853.995 2914.100 854.165 ;
        RECT 5.605 852.905 6.815 853.995 ;
        RECT 6.295 852.365 6.815 852.905 ;
        RECT 2910.045 852.830 2910.335 853.995 ;
        RECT 2912.805 852.905 2914.015 853.995 ;
        RECT 2912.805 852.365 2913.325 852.905 ;
        RECT 6.295 849.815 6.815 850.355 ;
        RECT 5.605 848.725 6.815 849.815 ;
        RECT 2912.805 849.815 2913.325 850.355 ;
        RECT 2912.805 848.725 2914.015 849.815 ;
        RECT 5.520 848.555 6.900 848.725 ;
        RECT 2909.960 848.555 2910.420 848.725 ;
        RECT 2912.720 848.555 2914.100 848.725 ;
        RECT 5.605 847.465 6.815 848.555 ;
        RECT 6.295 846.925 6.815 847.465 ;
        RECT 2910.045 847.390 2910.335 848.555 ;
        RECT 2912.805 847.465 2914.015 848.555 ;
        RECT 2912.805 846.925 2913.325 847.465 ;
        RECT 6.295 844.375 6.815 844.915 ;
        RECT 5.605 843.285 6.815 844.375 ;
        RECT 2912.805 844.375 2913.325 844.915 ;
        RECT 2912.805 843.285 2914.015 844.375 ;
        RECT 5.520 843.115 6.900 843.285 ;
        RECT 2909.960 843.115 2910.420 843.285 ;
        RECT 2912.720 843.115 2914.100 843.285 ;
        RECT 5.605 842.025 6.815 843.115 ;
        RECT 6.295 841.485 6.815 842.025 ;
        RECT 2910.045 841.950 2910.335 843.115 ;
        RECT 2912.805 842.025 2914.015 843.115 ;
        RECT 2912.805 841.485 2913.325 842.025 ;
        RECT 6.295 838.935 6.815 839.475 ;
        RECT 5.605 837.845 6.815 838.935 ;
        RECT 2912.805 838.935 2913.325 839.475 ;
        RECT 2912.805 837.845 2914.015 838.935 ;
        RECT 5.520 837.675 6.900 837.845 ;
        RECT 2909.960 837.675 2910.420 837.845 ;
        RECT 2912.720 837.675 2914.100 837.845 ;
        RECT 5.605 836.585 6.815 837.675 ;
        RECT 6.295 836.045 6.815 836.585 ;
        RECT 2910.045 836.510 2910.335 837.675 ;
        RECT 2912.805 836.585 2914.015 837.675 ;
        RECT 2912.805 836.045 2913.325 836.585 ;
        RECT 6.295 833.495 6.815 834.035 ;
        RECT 5.605 832.405 6.815 833.495 ;
        RECT 2912.805 833.495 2913.325 834.035 ;
        RECT 2912.805 832.405 2914.015 833.495 ;
        RECT 5.520 832.235 6.900 832.405 ;
        RECT 2909.960 832.235 2910.420 832.405 ;
        RECT 2912.720 832.235 2914.100 832.405 ;
        RECT 5.605 831.145 6.815 832.235 ;
        RECT 6.295 830.605 6.815 831.145 ;
        RECT 2910.045 831.070 2910.335 832.235 ;
        RECT 2912.805 831.145 2914.015 832.235 ;
        RECT 2912.805 830.605 2913.325 831.145 ;
        RECT 6.295 828.055 6.815 828.595 ;
        RECT 5.605 826.965 6.815 828.055 ;
        RECT 2912.805 828.055 2913.325 828.595 ;
        RECT 2912.805 826.965 2914.015 828.055 ;
        RECT 5.520 826.795 6.900 826.965 ;
        RECT 2909.960 826.795 2910.420 826.965 ;
        RECT 2912.720 826.795 2914.100 826.965 ;
        RECT 5.605 825.705 6.815 826.795 ;
        RECT 6.295 825.165 6.815 825.705 ;
        RECT 2910.045 825.630 2910.335 826.795 ;
        RECT 2912.805 825.705 2914.015 826.795 ;
        RECT 2912.805 825.165 2913.325 825.705 ;
        RECT 6.295 822.615 6.815 823.155 ;
        RECT 5.605 821.525 6.815 822.615 ;
        RECT 2912.805 822.615 2913.325 823.155 ;
        RECT 2912.805 821.525 2914.015 822.615 ;
        RECT 5.520 821.355 6.900 821.525 ;
        RECT 2909.960 821.355 2910.420 821.525 ;
        RECT 2912.720 821.355 2914.100 821.525 ;
        RECT 5.605 820.265 6.815 821.355 ;
        RECT 6.295 819.725 6.815 820.265 ;
        RECT 2910.045 820.190 2910.335 821.355 ;
        RECT 2912.805 820.265 2914.015 821.355 ;
        RECT 2912.805 819.725 2913.325 820.265 ;
        RECT 6.295 817.175 6.815 817.715 ;
        RECT 5.605 816.085 6.815 817.175 ;
        RECT 2912.805 817.175 2913.325 817.715 ;
        RECT 2912.805 816.085 2914.015 817.175 ;
        RECT 5.520 815.915 6.900 816.085 ;
        RECT 2909.960 815.915 2910.420 816.085 ;
        RECT 2912.720 815.915 2914.100 816.085 ;
        RECT 5.605 814.825 6.815 815.915 ;
        RECT 6.295 814.285 6.815 814.825 ;
        RECT 2910.045 814.750 2910.335 815.915 ;
        RECT 2912.805 814.825 2914.015 815.915 ;
        RECT 2912.805 814.285 2913.325 814.825 ;
        RECT 6.295 811.735 6.815 812.275 ;
        RECT 5.605 810.645 6.815 811.735 ;
        RECT 2912.805 811.735 2913.325 812.275 ;
        RECT 2909.315 810.645 2909.645 811.370 ;
        RECT 2912.805 810.645 2914.015 811.735 ;
        RECT 5.520 810.475 6.900 810.645 ;
        RECT 2909.040 810.475 2910.420 810.645 ;
        RECT 2912.720 810.475 2914.100 810.645 ;
        RECT 5.605 809.385 6.815 810.475 ;
        RECT 6.295 808.845 6.815 809.385 ;
        RECT 2910.045 809.310 2910.335 810.475 ;
        RECT 2912.805 809.385 2914.015 810.475 ;
        RECT 2912.805 808.845 2913.325 809.385 ;
        RECT 6.295 806.295 6.815 806.835 ;
        RECT 5.605 805.205 6.815 806.295 ;
        RECT 2912.805 806.295 2913.325 806.835 ;
        RECT 2912.805 805.205 2914.015 806.295 ;
        RECT 5.520 805.035 6.900 805.205 ;
        RECT 2909.960 805.035 2910.420 805.205 ;
        RECT 2912.720 805.035 2914.100 805.205 ;
        RECT 5.605 803.945 6.815 805.035 ;
        RECT 6.295 803.405 6.815 803.945 ;
        RECT 2910.045 803.870 2910.335 805.035 ;
        RECT 2912.805 803.945 2914.015 805.035 ;
        RECT 2912.805 803.405 2913.325 803.945 ;
        RECT 6.295 800.855 6.815 801.395 ;
        RECT 5.605 799.765 6.815 800.855 ;
        RECT 2912.805 800.855 2913.325 801.395 ;
        RECT 2912.805 799.765 2914.015 800.855 ;
        RECT 5.520 799.595 6.900 799.765 ;
        RECT 2909.960 799.595 2910.420 799.765 ;
        RECT 2912.720 799.595 2914.100 799.765 ;
        RECT 5.605 798.505 6.815 799.595 ;
        RECT 6.295 797.965 6.815 798.505 ;
        RECT 2910.045 798.430 2910.335 799.595 ;
        RECT 2912.805 798.505 2914.015 799.595 ;
        RECT 2912.805 797.965 2913.325 798.505 ;
        RECT 6.295 795.415 6.815 795.955 ;
        RECT 5.605 794.325 6.815 795.415 ;
        RECT 2912.805 795.415 2913.325 795.955 ;
        RECT 2912.805 794.325 2914.015 795.415 ;
        RECT 5.520 794.155 6.900 794.325 ;
        RECT 2909.960 794.155 2910.420 794.325 ;
        RECT 2912.720 794.155 2914.100 794.325 ;
        RECT 5.605 793.065 6.815 794.155 ;
        RECT 6.295 792.525 6.815 793.065 ;
        RECT 2910.045 792.990 2910.335 794.155 ;
        RECT 2912.805 793.065 2914.015 794.155 ;
        RECT 2912.805 792.525 2913.325 793.065 ;
        RECT 6.295 789.975 6.815 790.515 ;
        RECT 5.605 788.885 6.815 789.975 ;
        RECT 2912.805 789.975 2913.325 790.515 ;
        RECT 2912.805 788.885 2914.015 789.975 ;
        RECT 5.520 788.715 6.900 788.885 ;
        RECT 2909.960 788.715 2910.420 788.885 ;
        RECT 2912.720 788.715 2914.100 788.885 ;
        RECT 5.605 787.625 6.815 788.715 ;
        RECT 6.295 787.085 6.815 787.625 ;
        RECT 2910.045 787.550 2910.335 788.715 ;
        RECT 2912.805 787.625 2914.015 788.715 ;
        RECT 2912.805 787.085 2913.325 787.625 ;
        RECT 6.295 784.535 6.815 785.075 ;
        RECT 5.605 783.445 6.815 784.535 ;
        RECT 2912.805 784.535 2913.325 785.075 ;
        RECT 2912.805 783.445 2914.015 784.535 ;
        RECT 5.520 783.275 6.900 783.445 ;
        RECT 2909.960 783.275 2910.420 783.445 ;
        RECT 2912.720 783.275 2914.100 783.445 ;
        RECT 5.605 782.185 6.815 783.275 ;
        RECT 6.295 781.645 6.815 782.185 ;
        RECT 2910.045 782.110 2910.335 783.275 ;
        RECT 2912.805 782.185 2914.015 783.275 ;
        RECT 2912.805 781.645 2913.325 782.185 ;
        RECT 6.295 779.095 6.815 779.635 ;
        RECT 5.605 778.005 6.815 779.095 ;
        RECT 2912.805 779.095 2913.325 779.635 ;
        RECT 2912.805 778.005 2914.015 779.095 ;
        RECT 5.520 777.835 6.900 778.005 ;
        RECT 2909.960 777.835 2910.420 778.005 ;
        RECT 2912.720 777.835 2914.100 778.005 ;
        RECT 5.605 776.745 6.815 777.835 ;
        RECT 6.295 776.205 6.815 776.745 ;
        RECT 2910.045 776.670 2910.335 777.835 ;
        RECT 2912.805 776.745 2914.015 777.835 ;
        RECT 2912.805 776.205 2913.325 776.745 ;
        RECT 6.295 773.655 6.815 774.195 ;
        RECT 5.605 772.565 6.815 773.655 ;
        RECT 2912.805 773.655 2913.325 774.195 ;
        RECT 2912.805 772.565 2914.015 773.655 ;
        RECT 5.520 772.395 6.900 772.565 ;
        RECT 2909.960 772.395 2910.420 772.565 ;
        RECT 2912.720 772.395 2914.100 772.565 ;
        RECT 5.605 771.305 6.815 772.395 ;
        RECT 6.295 770.765 6.815 771.305 ;
        RECT 2910.045 771.230 2910.335 772.395 ;
        RECT 2912.805 771.305 2914.015 772.395 ;
        RECT 2912.805 770.765 2913.325 771.305 ;
        RECT 6.295 768.215 6.815 768.755 ;
        RECT 5.605 767.125 6.815 768.215 ;
        RECT 2912.805 768.215 2913.325 768.755 ;
        RECT 2912.805 767.125 2914.015 768.215 ;
        RECT 5.520 766.955 6.900 767.125 ;
        RECT 2909.960 766.955 2910.420 767.125 ;
        RECT 2912.720 766.955 2914.100 767.125 ;
        RECT 5.605 765.865 6.815 766.955 ;
        RECT 6.295 765.325 6.815 765.865 ;
        RECT 2910.045 765.790 2910.335 766.955 ;
        RECT 2912.805 765.865 2914.015 766.955 ;
        RECT 2912.805 765.325 2913.325 765.865 ;
        RECT 6.295 762.775 6.815 763.315 ;
        RECT 5.605 761.685 6.815 762.775 ;
        RECT 2912.805 762.775 2913.325 763.315 ;
        RECT 2912.805 761.685 2914.015 762.775 ;
        RECT 5.520 761.515 6.900 761.685 ;
        RECT 2909.960 761.515 2910.420 761.685 ;
        RECT 2912.720 761.515 2914.100 761.685 ;
        RECT 5.605 760.425 6.815 761.515 ;
        RECT 6.295 759.885 6.815 760.425 ;
        RECT 2910.045 760.350 2910.335 761.515 ;
        RECT 2912.805 760.425 2914.015 761.515 ;
        RECT 2912.805 759.885 2913.325 760.425 ;
        RECT 6.295 757.335 6.815 757.875 ;
        RECT 5.605 756.245 6.815 757.335 ;
        RECT 2912.805 757.335 2913.325 757.875 ;
        RECT 2912.805 756.245 2914.015 757.335 ;
        RECT 5.520 756.075 6.900 756.245 ;
        RECT 2909.960 756.075 2910.420 756.245 ;
        RECT 2912.720 756.075 2914.100 756.245 ;
        RECT 5.605 754.985 6.815 756.075 ;
        RECT 6.295 754.445 6.815 754.985 ;
        RECT 2910.045 754.910 2910.335 756.075 ;
        RECT 2912.805 754.985 2914.015 756.075 ;
        RECT 2912.805 754.445 2913.325 754.985 ;
        RECT 6.295 751.895 6.815 752.435 ;
        RECT 5.605 750.805 6.815 751.895 ;
        RECT 2912.805 751.895 2913.325 752.435 ;
        RECT 2912.805 750.805 2914.015 751.895 ;
        RECT 5.520 750.635 6.900 750.805 ;
        RECT 2909.960 750.635 2910.420 750.805 ;
        RECT 2912.720 750.635 2914.100 750.805 ;
        RECT 5.605 749.545 6.815 750.635 ;
        RECT 6.295 749.005 6.815 749.545 ;
        RECT 2910.045 749.470 2910.335 750.635 ;
        RECT 2912.805 749.545 2914.015 750.635 ;
        RECT 2912.805 749.005 2913.325 749.545 ;
        RECT 6.295 746.455 6.815 746.995 ;
        RECT 5.605 745.365 6.815 746.455 ;
        RECT 2912.805 746.455 2913.325 746.995 ;
        RECT 2912.805 745.365 2914.015 746.455 ;
        RECT 5.520 745.195 6.900 745.365 ;
        RECT 2909.960 745.195 2910.420 745.365 ;
        RECT 2912.720 745.195 2914.100 745.365 ;
        RECT 5.605 744.105 6.815 745.195 ;
        RECT 6.295 743.565 6.815 744.105 ;
        RECT 2910.045 744.030 2910.335 745.195 ;
        RECT 2912.805 744.105 2914.015 745.195 ;
        RECT 2912.805 743.565 2913.325 744.105 ;
        RECT 6.295 741.015 6.815 741.555 ;
        RECT 5.605 739.925 6.815 741.015 ;
        RECT 2912.805 741.015 2913.325 741.555 ;
        RECT 2912.805 739.925 2914.015 741.015 ;
        RECT 5.520 739.755 6.900 739.925 ;
        RECT 2909.960 739.755 2910.420 739.925 ;
        RECT 2912.720 739.755 2914.100 739.925 ;
        RECT 5.605 738.665 6.815 739.755 ;
        RECT 6.295 738.125 6.815 738.665 ;
        RECT 2910.045 738.590 2910.335 739.755 ;
        RECT 2912.805 738.665 2914.015 739.755 ;
        RECT 2912.805 738.125 2913.325 738.665 ;
        RECT 6.295 735.575 6.815 736.115 ;
        RECT 5.605 734.485 6.815 735.575 ;
        RECT 2912.805 735.575 2913.325 736.115 ;
        RECT 2909.315 734.485 2909.645 735.210 ;
        RECT 2912.805 734.485 2914.015 735.575 ;
        RECT 5.520 734.315 6.900 734.485 ;
        RECT 2909.040 734.315 2910.420 734.485 ;
        RECT 2912.720 734.315 2914.100 734.485 ;
        RECT 5.605 733.225 6.815 734.315 ;
        RECT 6.295 732.685 6.815 733.225 ;
        RECT 2910.045 733.150 2910.335 734.315 ;
        RECT 2912.805 733.225 2914.015 734.315 ;
        RECT 2912.805 732.685 2913.325 733.225 ;
        RECT 6.295 730.135 6.815 730.675 ;
        RECT 5.605 729.045 6.815 730.135 ;
        RECT 2912.805 730.135 2913.325 730.675 ;
        RECT 2912.805 729.045 2914.015 730.135 ;
        RECT 5.520 728.875 6.900 729.045 ;
        RECT 2909.960 728.875 2910.420 729.045 ;
        RECT 2912.720 728.875 2914.100 729.045 ;
        RECT 5.605 727.785 6.815 728.875 ;
        RECT 6.295 727.245 6.815 727.785 ;
        RECT 2910.045 727.710 2910.335 728.875 ;
        RECT 2912.805 727.785 2914.015 728.875 ;
        RECT 2912.805 727.245 2913.325 727.785 ;
        RECT 6.295 724.695 6.815 725.235 ;
        RECT 5.605 723.605 6.815 724.695 ;
        RECT 2912.805 724.695 2913.325 725.235 ;
        RECT 2912.805 723.605 2914.015 724.695 ;
        RECT 5.520 723.435 6.900 723.605 ;
        RECT 8.740 723.435 10.120 723.605 ;
        RECT 2909.960 723.435 2910.420 723.605 ;
        RECT 2912.720 723.435 2914.100 723.605 ;
        RECT 5.605 722.345 6.815 723.435 ;
        RECT 9.015 722.710 9.345 723.435 ;
        RECT 6.295 721.805 6.815 722.345 ;
        RECT 2910.045 722.270 2910.335 723.435 ;
        RECT 2912.805 722.345 2914.015 723.435 ;
        RECT 2912.805 721.805 2913.325 722.345 ;
        RECT 6.295 719.255 6.815 719.795 ;
        RECT 5.605 718.165 6.815 719.255 ;
        RECT 2912.805 719.255 2913.325 719.795 ;
        RECT 2912.805 718.165 2914.015 719.255 ;
        RECT 5.520 717.995 6.900 718.165 ;
        RECT 2909.960 717.995 2910.420 718.165 ;
        RECT 2912.720 717.995 2914.100 718.165 ;
        RECT 5.605 716.905 6.815 717.995 ;
        RECT 6.295 716.365 6.815 716.905 ;
        RECT 2910.045 716.830 2910.335 717.995 ;
        RECT 2912.805 716.905 2914.015 717.995 ;
        RECT 2912.805 716.365 2913.325 716.905 ;
        RECT 6.295 713.815 6.815 714.355 ;
        RECT 5.605 712.725 6.815 713.815 ;
        RECT 2912.805 713.815 2913.325 714.355 ;
        RECT 2912.805 712.725 2914.015 713.815 ;
        RECT 5.520 712.555 6.900 712.725 ;
        RECT 2909.960 712.555 2910.420 712.725 ;
        RECT 2912.720 712.555 2914.100 712.725 ;
        RECT 5.605 711.465 6.815 712.555 ;
        RECT 6.295 710.925 6.815 711.465 ;
        RECT 2910.045 711.390 2910.335 712.555 ;
        RECT 2912.805 711.465 2914.015 712.555 ;
        RECT 2912.805 710.925 2913.325 711.465 ;
        RECT 6.295 708.375 6.815 708.915 ;
        RECT 5.605 707.285 6.815 708.375 ;
        RECT 2912.805 708.375 2913.325 708.915 ;
        RECT 2912.805 707.285 2914.015 708.375 ;
        RECT 5.520 707.115 6.900 707.285 ;
        RECT 2909.960 707.115 2910.420 707.285 ;
        RECT 2912.720 707.115 2914.100 707.285 ;
        RECT 5.605 706.025 6.815 707.115 ;
        RECT 6.295 705.485 6.815 706.025 ;
        RECT 2910.045 705.950 2910.335 707.115 ;
        RECT 2912.805 706.025 2914.015 707.115 ;
        RECT 2912.805 705.485 2913.325 706.025 ;
        RECT 6.295 702.935 6.815 703.475 ;
        RECT 5.605 701.845 6.815 702.935 ;
        RECT 2912.805 702.935 2913.325 703.475 ;
        RECT 2912.805 701.845 2914.015 702.935 ;
        RECT 5.520 701.675 6.900 701.845 ;
        RECT 2909.960 701.675 2910.420 701.845 ;
        RECT 2912.720 701.675 2914.100 701.845 ;
        RECT 5.605 700.585 6.815 701.675 ;
        RECT 6.295 700.045 6.815 700.585 ;
        RECT 2910.045 700.510 2910.335 701.675 ;
        RECT 2912.805 700.585 2914.015 701.675 ;
        RECT 2912.805 700.045 2913.325 700.585 ;
        RECT 6.295 697.495 6.815 698.035 ;
        RECT 5.605 696.405 6.815 697.495 ;
        RECT 2912.805 697.495 2913.325 698.035 ;
        RECT 2912.805 696.405 2914.015 697.495 ;
        RECT 5.520 696.235 6.900 696.405 ;
        RECT 2909.960 696.235 2910.420 696.405 ;
        RECT 2912.720 696.235 2914.100 696.405 ;
        RECT 5.605 695.145 6.815 696.235 ;
        RECT 6.295 694.605 6.815 695.145 ;
        RECT 2910.045 695.070 2910.335 696.235 ;
        RECT 2912.805 695.145 2914.015 696.235 ;
        RECT 2912.805 694.605 2913.325 695.145 ;
        RECT 6.295 692.055 6.815 692.595 ;
        RECT 5.605 690.965 6.815 692.055 ;
        RECT 2912.805 692.055 2913.325 692.595 ;
        RECT 2912.805 690.965 2914.015 692.055 ;
        RECT 5.520 690.795 6.900 690.965 ;
        RECT 2909.960 690.795 2910.420 690.965 ;
        RECT 2912.720 690.795 2914.100 690.965 ;
        RECT 5.605 689.705 6.815 690.795 ;
        RECT 6.295 689.165 6.815 689.705 ;
        RECT 2910.045 689.630 2910.335 690.795 ;
        RECT 2912.805 689.705 2914.015 690.795 ;
        RECT 2912.805 689.165 2913.325 689.705 ;
        RECT 6.295 686.615 6.815 687.155 ;
        RECT 5.605 685.525 6.815 686.615 ;
        RECT 2912.805 686.615 2913.325 687.155 ;
        RECT 2912.805 685.525 2914.015 686.615 ;
        RECT 5.520 685.355 6.900 685.525 ;
        RECT 2909.960 685.355 2910.420 685.525 ;
        RECT 2912.720 685.355 2914.100 685.525 ;
        RECT 5.605 684.265 6.815 685.355 ;
        RECT 6.295 683.725 6.815 684.265 ;
        RECT 2910.045 684.190 2910.335 685.355 ;
        RECT 2912.805 684.265 2914.015 685.355 ;
        RECT 2912.805 683.725 2913.325 684.265 ;
        RECT 6.295 681.175 6.815 681.715 ;
        RECT 5.605 680.085 6.815 681.175 ;
        RECT 2912.805 681.175 2913.325 681.715 ;
        RECT 2912.805 680.085 2914.015 681.175 ;
        RECT 5.520 679.915 6.900 680.085 ;
        RECT 2909.960 679.915 2910.420 680.085 ;
        RECT 2912.720 679.915 2914.100 680.085 ;
        RECT 5.605 678.825 6.815 679.915 ;
        RECT 6.295 678.285 6.815 678.825 ;
        RECT 2910.045 678.750 2910.335 679.915 ;
        RECT 2912.805 678.825 2914.015 679.915 ;
        RECT 2912.805 678.285 2913.325 678.825 ;
        RECT 6.295 675.735 6.815 676.275 ;
        RECT 5.605 674.645 6.815 675.735 ;
        RECT 2912.805 675.735 2913.325 676.275 ;
        RECT 2912.805 674.645 2914.015 675.735 ;
        RECT 5.520 674.475 6.900 674.645 ;
        RECT 2909.960 674.475 2910.420 674.645 ;
        RECT 2912.720 674.475 2914.100 674.645 ;
        RECT 5.605 673.385 6.815 674.475 ;
        RECT 6.295 672.845 6.815 673.385 ;
        RECT 2910.045 673.310 2910.335 674.475 ;
        RECT 2912.805 673.385 2914.015 674.475 ;
        RECT 2912.805 672.845 2913.325 673.385 ;
        RECT 6.295 670.295 6.815 670.835 ;
        RECT 5.605 669.205 6.815 670.295 ;
        RECT 2912.805 670.295 2913.325 670.835 ;
        RECT 2912.805 669.205 2914.015 670.295 ;
        RECT 5.520 669.035 6.900 669.205 ;
        RECT 2909.960 669.035 2910.420 669.205 ;
        RECT 2912.720 669.035 2914.100 669.205 ;
        RECT 5.605 667.945 6.815 669.035 ;
        RECT 6.295 667.405 6.815 667.945 ;
        RECT 2910.045 667.870 2910.335 669.035 ;
        RECT 2912.805 667.945 2914.015 669.035 ;
        RECT 2912.805 667.405 2913.325 667.945 ;
        RECT 6.295 664.855 6.815 665.395 ;
        RECT 5.605 663.765 6.815 664.855 ;
        RECT 2912.805 664.855 2913.325 665.395 ;
        RECT 2912.805 663.765 2914.015 664.855 ;
        RECT 5.520 663.595 6.900 663.765 ;
        RECT 2909.960 663.595 2910.420 663.765 ;
        RECT 2912.720 663.595 2914.100 663.765 ;
        RECT 5.605 662.505 6.815 663.595 ;
        RECT 6.295 661.965 6.815 662.505 ;
        RECT 2910.045 662.430 2910.335 663.595 ;
        RECT 2912.805 662.505 2914.015 663.595 ;
        RECT 2912.805 661.965 2913.325 662.505 ;
        RECT 6.295 659.415 6.815 659.955 ;
        RECT 5.605 658.325 6.815 659.415 ;
        RECT 2912.805 659.415 2913.325 659.955 ;
        RECT 2912.805 658.325 2914.015 659.415 ;
        RECT 5.520 658.155 6.900 658.325 ;
        RECT 2909.960 658.155 2910.420 658.325 ;
        RECT 2912.720 658.155 2914.100 658.325 ;
        RECT 5.605 657.065 6.815 658.155 ;
        RECT 6.295 656.525 6.815 657.065 ;
        RECT 2910.045 656.990 2910.335 658.155 ;
        RECT 2912.805 657.065 2914.015 658.155 ;
        RECT 2912.805 656.525 2913.325 657.065 ;
        RECT 6.295 653.975 6.815 654.515 ;
        RECT 5.605 652.885 6.815 653.975 ;
        RECT 2912.805 653.975 2913.325 654.515 ;
        RECT 2912.805 652.885 2914.015 653.975 ;
        RECT 5.520 652.715 6.900 652.885 ;
        RECT 2909.960 652.715 2910.420 652.885 ;
        RECT 2912.720 652.715 2914.100 652.885 ;
        RECT 5.605 651.625 6.815 652.715 ;
        RECT 6.295 651.085 6.815 651.625 ;
        RECT 2910.045 651.550 2910.335 652.715 ;
        RECT 2912.805 651.625 2914.015 652.715 ;
        RECT 2912.805 651.085 2913.325 651.625 ;
        RECT 6.295 648.535 6.815 649.075 ;
        RECT 5.605 647.445 6.815 648.535 ;
        RECT 2912.805 648.535 2913.325 649.075 ;
        RECT 2912.805 647.445 2914.015 648.535 ;
        RECT 5.520 647.275 6.900 647.445 ;
        RECT 2909.960 647.275 2910.420 647.445 ;
        RECT 2912.720 647.275 2914.100 647.445 ;
        RECT 5.605 646.185 6.815 647.275 ;
        RECT 6.295 645.645 6.815 646.185 ;
        RECT 2910.045 646.110 2910.335 647.275 ;
        RECT 2912.805 646.185 2914.015 647.275 ;
        RECT 2912.805 645.645 2913.325 646.185 ;
        RECT 6.295 643.095 6.815 643.635 ;
        RECT 5.605 642.005 6.815 643.095 ;
        RECT 2912.805 643.095 2913.325 643.635 ;
        RECT 2912.805 642.005 2914.015 643.095 ;
        RECT 5.520 641.835 6.900 642.005 ;
        RECT 2909.960 641.835 2910.420 642.005 ;
        RECT 2912.720 641.835 2914.100 642.005 ;
        RECT 5.605 640.745 6.815 641.835 ;
        RECT 6.295 640.205 6.815 640.745 ;
        RECT 2910.045 640.670 2910.335 641.835 ;
        RECT 2912.805 640.745 2914.015 641.835 ;
        RECT 2912.805 640.205 2913.325 640.745 ;
        RECT 6.295 637.655 6.815 638.195 ;
        RECT 5.605 636.565 6.815 637.655 ;
        RECT 2912.805 637.655 2913.325 638.195 ;
        RECT 2912.805 636.565 2914.015 637.655 ;
        RECT 5.520 636.395 6.900 636.565 ;
        RECT 2909.960 636.395 2910.420 636.565 ;
        RECT 2912.720 636.395 2914.100 636.565 ;
        RECT 5.605 635.305 6.815 636.395 ;
        RECT 6.295 634.765 6.815 635.305 ;
        RECT 2910.045 635.230 2910.335 636.395 ;
        RECT 2912.805 635.305 2914.015 636.395 ;
        RECT 2912.805 634.765 2913.325 635.305 ;
        RECT 6.295 632.215 6.815 632.755 ;
        RECT 5.605 631.125 6.815 632.215 ;
        RECT 2912.805 632.215 2913.325 632.755 ;
        RECT 2912.805 631.125 2914.015 632.215 ;
        RECT 5.520 630.955 6.900 631.125 ;
        RECT 8.740 630.955 10.120 631.125 ;
        RECT 2909.960 630.955 2910.420 631.125 ;
        RECT 2912.720 630.955 2914.100 631.125 ;
        RECT 5.605 629.865 6.815 630.955 ;
        RECT 9.015 630.230 9.345 630.955 ;
        RECT 6.295 629.325 6.815 629.865 ;
        RECT 2910.045 629.790 2910.335 630.955 ;
        RECT 2912.805 629.865 2914.015 630.955 ;
        RECT 2912.805 629.325 2913.325 629.865 ;
        RECT 6.295 626.775 6.815 627.315 ;
        RECT 5.605 625.685 6.815 626.775 ;
        RECT 2912.805 626.775 2913.325 627.315 ;
        RECT 2912.805 625.685 2914.015 626.775 ;
        RECT 5.520 625.515 6.900 625.685 ;
        RECT 2909.960 625.515 2910.420 625.685 ;
        RECT 2912.720 625.515 2914.100 625.685 ;
        RECT 5.605 624.425 6.815 625.515 ;
        RECT 6.295 623.885 6.815 624.425 ;
        RECT 2910.045 624.350 2910.335 625.515 ;
        RECT 2912.805 624.425 2914.015 625.515 ;
        RECT 2912.805 623.885 2913.325 624.425 ;
        RECT 6.295 621.335 6.815 621.875 ;
        RECT 5.605 620.245 6.815 621.335 ;
        RECT 2912.805 621.335 2913.325 621.875 ;
        RECT 2912.805 620.245 2914.015 621.335 ;
        RECT 5.520 620.075 6.900 620.245 ;
        RECT 2909.960 620.075 2910.420 620.245 ;
        RECT 2912.720 620.075 2914.100 620.245 ;
        RECT 5.605 618.985 6.815 620.075 ;
        RECT 6.295 618.445 6.815 618.985 ;
        RECT 2910.045 618.910 2910.335 620.075 ;
        RECT 2912.805 618.985 2914.015 620.075 ;
        RECT 2912.805 618.445 2913.325 618.985 ;
        RECT 6.295 615.895 6.815 616.435 ;
        RECT 5.605 614.805 6.815 615.895 ;
        RECT 2912.805 615.895 2913.325 616.435 ;
        RECT 2912.805 614.805 2914.015 615.895 ;
        RECT 5.520 614.635 6.900 614.805 ;
        RECT 2909.960 614.635 2910.420 614.805 ;
        RECT 2912.720 614.635 2914.100 614.805 ;
        RECT 5.605 613.545 6.815 614.635 ;
        RECT 6.295 613.005 6.815 613.545 ;
        RECT 2910.045 613.470 2910.335 614.635 ;
        RECT 2912.805 613.545 2914.015 614.635 ;
        RECT 2912.805 613.005 2913.325 613.545 ;
        RECT 6.295 610.455 6.815 610.995 ;
        RECT 5.605 609.365 6.815 610.455 ;
        RECT 2912.805 610.455 2913.325 610.995 ;
        RECT 2912.805 609.365 2914.015 610.455 ;
        RECT 5.520 609.195 6.900 609.365 ;
        RECT 2909.960 609.195 2910.420 609.365 ;
        RECT 2912.720 609.195 2914.100 609.365 ;
        RECT 5.605 608.105 6.815 609.195 ;
        RECT 6.295 607.565 6.815 608.105 ;
        RECT 2910.045 608.030 2910.335 609.195 ;
        RECT 2912.805 608.105 2914.015 609.195 ;
        RECT 2912.805 607.565 2913.325 608.105 ;
        RECT 6.295 605.015 6.815 605.555 ;
        RECT 5.605 603.925 6.815 605.015 ;
        RECT 2912.805 605.015 2913.325 605.555 ;
        RECT 2912.805 603.925 2914.015 605.015 ;
        RECT 5.520 603.755 6.900 603.925 ;
        RECT 8.740 603.755 10.120 603.925 ;
        RECT 2909.960 603.755 2910.420 603.925 ;
        RECT 2912.720 603.755 2914.100 603.925 ;
        RECT 5.605 602.665 6.815 603.755 ;
        RECT 9.015 603.030 9.345 603.755 ;
        RECT 6.295 602.125 6.815 602.665 ;
        RECT 2910.045 602.590 2910.335 603.755 ;
        RECT 2912.805 602.665 2914.015 603.755 ;
        RECT 2912.805 602.125 2913.325 602.665 ;
        RECT 6.295 599.575 6.815 600.115 ;
        RECT 5.605 598.485 6.815 599.575 ;
        RECT 2912.805 599.575 2913.325 600.115 ;
        RECT 2912.805 598.485 2914.015 599.575 ;
        RECT 5.520 598.315 6.900 598.485 ;
        RECT 2909.960 598.315 2910.420 598.485 ;
        RECT 2912.720 598.315 2914.100 598.485 ;
        RECT 5.605 597.225 6.815 598.315 ;
        RECT 6.295 596.685 6.815 597.225 ;
        RECT 2910.045 597.150 2910.335 598.315 ;
        RECT 2912.805 597.225 2914.015 598.315 ;
        RECT 2912.805 596.685 2913.325 597.225 ;
        RECT 6.295 594.135 6.815 594.675 ;
        RECT 5.605 593.045 6.815 594.135 ;
        RECT 2912.805 594.135 2913.325 594.675 ;
        RECT 2912.805 593.045 2914.015 594.135 ;
        RECT 5.520 592.875 6.900 593.045 ;
        RECT 2909.960 592.875 2910.420 593.045 ;
        RECT 2912.720 592.875 2914.100 593.045 ;
        RECT 5.605 591.785 6.815 592.875 ;
        RECT 6.295 591.245 6.815 591.785 ;
        RECT 2910.045 591.710 2910.335 592.875 ;
        RECT 2912.805 591.785 2914.015 592.875 ;
        RECT 2912.805 591.245 2913.325 591.785 ;
        RECT 6.295 588.695 6.815 589.235 ;
        RECT 5.605 587.605 6.815 588.695 ;
        RECT 2912.805 588.695 2913.325 589.235 ;
        RECT 2912.805 587.605 2914.015 588.695 ;
        RECT 5.520 587.435 6.900 587.605 ;
        RECT 2909.960 587.435 2910.420 587.605 ;
        RECT 2912.720 587.435 2914.100 587.605 ;
        RECT 5.605 586.345 6.815 587.435 ;
        RECT 6.295 585.805 6.815 586.345 ;
        RECT 2910.045 586.270 2910.335 587.435 ;
        RECT 2912.805 586.345 2914.015 587.435 ;
        RECT 2912.805 585.805 2913.325 586.345 ;
        RECT 6.295 583.255 6.815 583.795 ;
        RECT 5.605 582.165 6.815 583.255 ;
        RECT 2912.805 583.255 2913.325 583.795 ;
        RECT 2912.805 582.165 2914.015 583.255 ;
        RECT 5.520 581.995 6.900 582.165 ;
        RECT 2909.960 581.995 2910.420 582.165 ;
        RECT 2912.720 581.995 2914.100 582.165 ;
        RECT 5.605 580.905 6.815 581.995 ;
        RECT 6.295 580.365 6.815 580.905 ;
        RECT 2910.045 580.830 2910.335 581.995 ;
        RECT 2912.805 580.905 2914.015 581.995 ;
        RECT 2912.805 580.365 2913.325 580.905 ;
        RECT 6.295 577.815 6.815 578.355 ;
        RECT 5.605 576.725 6.815 577.815 ;
        RECT 2912.805 577.815 2913.325 578.355 ;
        RECT 2912.805 576.725 2914.015 577.815 ;
        RECT 5.520 576.555 6.900 576.725 ;
        RECT 2909.960 576.555 2910.420 576.725 ;
        RECT 2912.720 576.555 2914.100 576.725 ;
        RECT 5.605 575.465 6.815 576.555 ;
        RECT 6.295 574.925 6.815 575.465 ;
        RECT 2910.045 575.390 2910.335 576.555 ;
        RECT 2912.805 575.465 2914.015 576.555 ;
        RECT 2912.805 574.925 2913.325 575.465 ;
        RECT 6.295 572.375 6.815 572.915 ;
        RECT 5.605 571.285 6.815 572.375 ;
        RECT 2912.805 572.375 2913.325 572.915 ;
        RECT 2912.805 571.285 2914.015 572.375 ;
        RECT 5.520 571.115 6.900 571.285 ;
        RECT 2909.960 571.115 2910.420 571.285 ;
        RECT 2912.720 571.115 2914.100 571.285 ;
        RECT 5.605 570.025 6.815 571.115 ;
        RECT 6.295 569.485 6.815 570.025 ;
        RECT 2910.045 569.950 2910.335 571.115 ;
        RECT 2912.805 570.025 2914.015 571.115 ;
        RECT 2912.805 569.485 2913.325 570.025 ;
        RECT 6.295 566.935 6.815 567.475 ;
        RECT 5.605 565.845 6.815 566.935 ;
        RECT 2912.805 566.935 2913.325 567.475 ;
        RECT 2912.805 565.845 2914.015 566.935 ;
        RECT 5.520 565.675 6.900 565.845 ;
        RECT 2909.960 565.675 2910.420 565.845 ;
        RECT 2912.720 565.675 2914.100 565.845 ;
        RECT 5.605 564.585 6.815 565.675 ;
        RECT 6.295 564.045 6.815 564.585 ;
        RECT 2910.045 564.510 2910.335 565.675 ;
        RECT 2912.805 564.585 2914.015 565.675 ;
        RECT 2912.805 564.045 2913.325 564.585 ;
        RECT 6.295 561.495 6.815 562.035 ;
        RECT 5.605 560.405 6.815 561.495 ;
        RECT 2912.805 561.495 2913.325 562.035 ;
        RECT 2912.805 560.405 2914.015 561.495 ;
        RECT 5.520 560.235 6.900 560.405 ;
        RECT 2909.960 560.235 2910.420 560.405 ;
        RECT 2912.720 560.235 2914.100 560.405 ;
        RECT 5.605 559.145 6.815 560.235 ;
        RECT 6.295 558.605 6.815 559.145 ;
        RECT 2910.045 559.070 2910.335 560.235 ;
        RECT 2912.805 559.145 2914.015 560.235 ;
        RECT 2912.805 558.605 2913.325 559.145 ;
        RECT 6.295 556.055 6.815 556.595 ;
        RECT 5.605 554.965 6.815 556.055 ;
        RECT 2912.805 556.055 2913.325 556.595 ;
        RECT 2912.805 554.965 2914.015 556.055 ;
        RECT 5.520 554.795 6.900 554.965 ;
        RECT 2909.960 554.795 2910.420 554.965 ;
        RECT 2912.720 554.795 2914.100 554.965 ;
        RECT 5.605 553.705 6.815 554.795 ;
        RECT 6.295 553.165 6.815 553.705 ;
        RECT 2910.045 553.630 2910.335 554.795 ;
        RECT 2912.805 553.705 2914.015 554.795 ;
        RECT 2912.805 553.165 2913.325 553.705 ;
        RECT 6.295 550.615 6.815 551.155 ;
        RECT 5.605 549.525 6.815 550.615 ;
        RECT 2912.805 550.615 2913.325 551.155 ;
        RECT 2912.805 549.525 2914.015 550.615 ;
        RECT 5.520 549.355 6.900 549.525 ;
        RECT 2909.960 549.355 2910.420 549.525 ;
        RECT 2912.720 549.355 2914.100 549.525 ;
        RECT 5.605 548.265 6.815 549.355 ;
        RECT 6.295 547.725 6.815 548.265 ;
        RECT 2910.045 548.190 2910.335 549.355 ;
        RECT 2912.805 548.265 2914.015 549.355 ;
        RECT 2912.805 547.725 2913.325 548.265 ;
        RECT 6.295 545.175 6.815 545.715 ;
        RECT 5.605 544.085 6.815 545.175 ;
        RECT 2912.805 545.175 2913.325 545.715 ;
        RECT 2912.805 544.085 2914.015 545.175 ;
        RECT 5.520 543.915 6.900 544.085 ;
        RECT 2909.960 543.915 2910.420 544.085 ;
        RECT 2912.720 543.915 2914.100 544.085 ;
        RECT 5.605 542.825 6.815 543.915 ;
        RECT 6.295 542.285 6.815 542.825 ;
        RECT 2910.045 542.750 2910.335 543.915 ;
        RECT 2912.805 542.825 2914.015 543.915 ;
        RECT 2912.805 542.285 2913.325 542.825 ;
        RECT 6.295 539.735 6.815 540.275 ;
        RECT 5.605 538.645 6.815 539.735 ;
        RECT 2912.805 539.735 2913.325 540.275 ;
        RECT 2912.805 538.645 2914.015 539.735 ;
        RECT 5.520 538.475 6.900 538.645 ;
        RECT 2909.960 538.475 2910.420 538.645 ;
        RECT 2912.720 538.475 2914.100 538.645 ;
        RECT 5.605 537.385 6.815 538.475 ;
        RECT 6.295 536.845 6.815 537.385 ;
        RECT 2910.045 537.310 2910.335 538.475 ;
        RECT 2912.805 537.385 2914.015 538.475 ;
        RECT 2912.805 536.845 2913.325 537.385 ;
        RECT 6.295 534.295 6.815 534.835 ;
        RECT 5.605 533.205 6.815 534.295 ;
        RECT 2912.805 534.295 2913.325 534.835 ;
        RECT 2912.805 533.205 2914.015 534.295 ;
        RECT 5.520 533.035 6.900 533.205 ;
        RECT 2909.960 533.035 2910.420 533.205 ;
        RECT 2912.720 533.035 2914.100 533.205 ;
        RECT 5.605 531.945 6.815 533.035 ;
        RECT 6.295 531.405 6.815 531.945 ;
        RECT 2910.045 531.870 2910.335 533.035 ;
        RECT 2912.805 531.945 2914.015 533.035 ;
        RECT 2912.805 531.405 2913.325 531.945 ;
        RECT 6.295 528.855 6.815 529.395 ;
        RECT 5.605 527.765 6.815 528.855 ;
        RECT 2912.805 528.855 2913.325 529.395 ;
        RECT 2912.805 527.765 2914.015 528.855 ;
        RECT 5.520 527.595 6.900 527.765 ;
        RECT 2909.960 527.595 2910.420 527.765 ;
        RECT 2912.720 527.595 2914.100 527.765 ;
        RECT 5.605 526.505 6.815 527.595 ;
        RECT 6.295 525.965 6.815 526.505 ;
        RECT 2910.045 526.430 2910.335 527.595 ;
        RECT 2912.805 526.505 2914.015 527.595 ;
        RECT 2912.805 525.965 2913.325 526.505 ;
        RECT 6.295 523.415 6.815 523.955 ;
        RECT 5.605 522.325 6.815 523.415 ;
        RECT 2912.805 523.415 2913.325 523.955 ;
        RECT 2912.805 522.325 2914.015 523.415 ;
        RECT 5.520 522.155 6.900 522.325 ;
        RECT 2909.960 522.155 2910.420 522.325 ;
        RECT 2912.720 522.155 2914.100 522.325 ;
        RECT 5.605 521.065 6.815 522.155 ;
        RECT 6.295 520.525 6.815 521.065 ;
        RECT 2910.045 520.990 2910.335 522.155 ;
        RECT 2912.805 521.065 2914.015 522.155 ;
        RECT 2912.805 520.525 2913.325 521.065 ;
        RECT 6.295 517.975 6.815 518.515 ;
        RECT 5.605 516.885 6.815 517.975 ;
        RECT 2912.805 517.975 2913.325 518.515 ;
        RECT 2912.805 516.885 2914.015 517.975 ;
        RECT 5.520 516.715 6.900 516.885 ;
        RECT 2909.960 516.715 2910.420 516.885 ;
        RECT 2912.720 516.715 2914.100 516.885 ;
        RECT 5.605 515.625 6.815 516.715 ;
        RECT 6.295 515.085 6.815 515.625 ;
        RECT 2910.045 515.550 2910.335 516.715 ;
        RECT 2912.805 515.625 2914.015 516.715 ;
        RECT 2912.805 515.085 2913.325 515.625 ;
        RECT 6.295 512.535 6.815 513.075 ;
        RECT 5.605 511.445 6.815 512.535 ;
        RECT 2912.805 512.535 2913.325 513.075 ;
        RECT 2912.805 511.445 2914.015 512.535 ;
        RECT 5.520 511.275 6.900 511.445 ;
        RECT 2909.960 511.275 2910.420 511.445 ;
        RECT 2912.720 511.275 2914.100 511.445 ;
        RECT 5.605 510.185 6.815 511.275 ;
        RECT 6.295 509.645 6.815 510.185 ;
        RECT 2910.045 510.110 2910.335 511.275 ;
        RECT 2912.805 510.185 2914.015 511.275 ;
        RECT 2912.805 509.645 2913.325 510.185 ;
        RECT 6.295 507.095 6.815 507.635 ;
        RECT 5.605 506.005 6.815 507.095 ;
        RECT 2912.805 507.095 2913.325 507.635 ;
        RECT 2912.805 506.005 2914.015 507.095 ;
        RECT 5.520 505.835 6.900 506.005 ;
        RECT 2909.960 505.835 2910.420 506.005 ;
        RECT 2912.720 505.835 2914.100 506.005 ;
        RECT 5.605 504.745 6.815 505.835 ;
        RECT 6.295 504.205 6.815 504.745 ;
        RECT 2910.045 504.670 2910.335 505.835 ;
        RECT 2912.805 504.745 2914.015 505.835 ;
        RECT 2912.805 504.205 2913.325 504.745 ;
        RECT 6.295 501.655 6.815 502.195 ;
        RECT 5.605 500.565 6.815 501.655 ;
        RECT 2912.805 501.655 2913.325 502.195 ;
        RECT 2912.805 500.565 2914.015 501.655 ;
        RECT 5.520 500.395 6.900 500.565 ;
        RECT 2909.960 500.395 2910.420 500.565 ;
        RECT 2912.720 500.395 2914.100 500.565 ;
        RECT 5.605 499.305 6.815 500.395 ;
        RECT 6.295 498.765 6.815 499.305 ;
        RECT 2910.045 499.230 2910.335 500.395 ;
        RECT 2912.805 499.305 2914.015 500.395 ;
        RECT 2912.805 498.765 2913.325 499.305 ;
        RECT 6.295 496.215 6.815 496.755 ;
        RECT 5.605 495.125 6.815 496.215 ;
        RECT 2912.805 496.215 2913.325 496.755 ;
        RECT 2912.805 495.125 2914.015 496.215 ;
        RECT 5.520 494.955 6.900 495.125 ;
        RECT 2909.960 494.955 2910.420 495.125 ;
        RECT 2912.720 494.955 2914.100 495.125 ;
        RECT 5.605 493.865 6.815 494.955 ;
        RECT 6.295 493.325 6.815 493.865 ;
        RECT 2910.045 493.790 2910.335 494.955 ;
        RECT 2912.805 493.865 2914.015 494.955 ;
        RECT 2912.805 493.325 2913.325 493.865 ;
        RECT 6.295 490.775 6.815 491.315 ;
        RECT 5.605 489.685 6.815 490.775 ;
        RECT 2912.805 490.775 2913.325 491.315 ;
        RECT 2912.805 489.685 2914.015 490.775 ;
        RECT 5.520 489.515 6.900 489.685 ;
        RECT 2909.960 489.515 2910.420 489.685 ;
        RECT 2912.720 489.515 2914.100 489.685 ;
        RECT 5.605 488.425 6.815 489.515 ;
        RECT 6.295 487.885 6.815 488.425 ;
        RECT 2910.045 488.350 2910.335 489.515 ;
        RECT 2912.805 488.425 2914.015 489.515 ;
        RECT 2912.805 487.885 2913.325 488.425 ;
        RECT 6.295 485.335 6.815 485.875 ;
        RECT 5.605 484.245 6.815 485.335 ;
        RECT 2912.805 485.335 2913.325 485.875 ;
        RECT 2912.805 484.245 2914.015 485.335 ;
        RECT 5.520 484.075 6.900 484.245 ;
        RECT 2909.960 484.075 2910.420 484.245 ;
        RECT 2912.720 484.075 2914.100 484.245 ;
        RECT 5.605 482.985 6.815 484.075 ;
        RECT 6.295 482.445 6.815 482.985 ;
        RECT 2910.045 482.910 2910.335 484.075 ;
        RECT 2912.805 482.985 2914.015 484.075 ;
        RECT 2912.805 482.445 2913.325 482.985 ;
        RECT 6.295 479.895 6.815 480.435 ;
        RECT 5.605 478.805 6.815 479.895 ;
        RECT 2912.805 479.895 2913.325 480.435 ;
        RECT 2912.805 478.805 2914.015 479.895 ;
        RECT 5.520 478.635 6.900 478.805 ;
        RECT 2909.960 478.635 2910.420 478.805 ;
        RECT 2912.720 478.635 2914.100 478.805 ;
        RECT 5.605 477.545 6.815 478.635 ;
        RECT 6.295 477.005 6.815 477.545 ;
        RECT 2910.045 477.470 2910.335 478.635 ;
        RECT 2912.805 477.545 2914.015 478.635 ;
        RECT 2912.805 477.005 2913.325 477.545 ;
        RECT 6.295 474.455 6.815 474.995 ;
        RECT 5.605 473.365 6.815 474.455 ;
        RECT 2912.805 474.455 2913.325 474.995 ;
        RECT 2912.805 473.365 2914.015 474.455 ;
        RECT 5.520 473.195 6.900 473.365 ;
        RECT 2909.960 473.195 2910.420 473.365 ;
        RECT 2912.720 473.195 2914.100 473.365 ;
        RECT 5.605 472.105 6.815 473.195 ;
        RECT 6.295 471.565 6.815 472.105 ;
        RECT 2910.045 472.030 2910.335 473.195 ;
        RECT 2912.805 472.105 2914.015 473.195 ;
        RECT 2912.805 471.565 2913.325 472.105 ;
        RECT 6.295 469.015 6.815 469.555 ;
        RECT 5.605 467.925 6.815 469.015 ;
        RECT 2912.805 469.015 2913.325 469.555 ;
        RECT 2909.315 467.925 2909.645 468.650 ;
        RECT 2912.805 467.925 2914.015 469.015 ;
        RECT 5.520 467.755 6.900 467.925 ;
        RECT 2909.040 467.755 2910.420 467.925 ;
        RECT 2912.720 467.755 2914.100 467.925 ;
        RECT 5.605 466.665 6.815 467.755 ;
        RECT 6.295 466.125 6.815 466.665 ;
        RECT 2910.045 466.590 2910.335 467.755 ;
        RECT 2912.805 466.665 2914.015 467.755 ;
        RECT 2912.805 466.125 2913.325 466.665 ;
        RECT 6.295 463.575 6.815 464.115 ;
        RECT 5.605 462.485 6.815 463.575 ;
        RECT 2912.805 463.575 2913.325 464.115 ;
        RECT 2912.805 462.485 2914.015 463.575 ;
        RECT 5.520 462.315 6.900 462.485 ;
        RECT 2909.960 462.315 2910.420 462.485 ;
        RECT 2912.720 462.315 2914.100 462.485 ;
        RECT 5.605 461.225 6.815 462.315 ;
        RECT 6.295 460.685 6.815 461.225 ;
        RECT 2910.045 461.150 2910.335 462.315 ;
        RECT 2912.805 461.225 2914.015 462.315 ;
        RECT 2912.805 460.685 2913.325 461.225 ;
        RECT 6.295 458.135 6.815 458.675 ;
        RECT 5.605 457.045 6.815 458.135 ;
        RECT 2912.805 458.135 2913.325 458.675 ;
        RECT 2912.805 457.045 2914.015 458.135 ;
        RECT 5.520 456.875 6.900 457.045 ;
        RECT 2909.960 456.875 2910.420 457.045 ;
        RECT 2912.720 456.875 2914.100 457.045 ;
        RECT 5.605 455.785 6.815 456.875 ;
        RECT 6.295 455.245 6.815 455.785 ;
        RECT 2910.045 455.710 2910.335 456.875 ;
        RECT 2912.805 455.785 2914.015 456.875 ;
        RECT 2912.805 455.245 2913.325 455.785 ;
        RECT 6.295 452.695 6.815 453.235 ;
        RECT 5.605 451.605 6.815 452.695 ;
        RECT 2912.805 452.695 2913.325 453.235 ;
        RECT 2912.805 451.605 2914.015 452.695 ;
        RECT 5.520 451.435 6.900 451.605 ;
        RECT 2909.960 451.435 2911.800 451.605 ;
        RECT 2912.720 451.435 2914.100 451.605 ;
        RECT 5.605 450.345 6.815 451.435 ;
        RECT 6.295 449.805 6.815 450.345 ;
        RECT 2910.045 450.270 2910.335 451.435 ;
        RECT 2910.695 450.710 2911.025 451.435 ;
        RECT 2912.805 450.345 2914.015 451.435 ;
        RECT 2912.805 449.805 2913.325 450.345 ;
        RECT 6.295 447.255 6.815 447.795 ;
        RECT 5.605 446.165 6.815 447.255 ;
        RECT 2912.805 447.255 2913.325 447.795 ;
        RECT 2912.805 446.165 2914.015 447.255 ;
        RECT 5.520 445.995 6.900 446.165 ;
        RECT 2909.960 445.995 2910.420 446.165 ;
        RECT 2912.720 445.995 2914.100 446.165 ;
        RECT 5.605 444.905 6.815 445.995 ;
        RECT 6.295 444.365 6.815 444.905 ;
        RECT 2910.045 444.830 2910.335 445.995 ;
        RECT 2912.805 444.905 2914.015 445.995 ;
        RECT 2912.805 444.365 2913.325 444.905 ;
        RECT 6.295 441.815 6.815 442.355 ;
        RECT 5.605 440.725 6.815 441.815 ;
        RECT 2912.805 441.815 2913.325 442.355 ;
        RECT 9.015 440.725 9.345 441.450 ;
        RECT 2912.805 440.725 2914.015 441.815 ;
        RECT 5.520 440.555 6.900 440.725 ;
        RECT 8.740 440.555 10.120 440.725 ;
        RECT 2909.960 440.555 2910.420 440.725 ;
        RECT 2912.720 440.555 2914.100 440.725 ;
        RECT 5.605 439.465 6.815 440.555 ;
        RECT 9.015 439.830 9.345 440.555 ;
        RECT 6.295 438.925 6.815 439.465 ;
        RECT 2910.045 439.390 2910.335 440.555 ;
        RECT 2912.805 439.465 2914.015 440.555 ;
        RECT 2912.805 438.925 2913.325 439.465 ;
        RECT 6.295 436.375 6.815 436.915 ;
        RECT 5.605 435.285 6.815 436.375 ;
        RECT 2912.805 436.375 2913.325 436.915 ;
        RECT 2912.805 435.285 2914.015 436.375 ;
        RECT 5.520 435.115 6.900 435.285 ;
        RECT 2909.960 435.115 2910.420 435.285 ;
        RECT 2912.720 435.115 2914.100 435.285 ;
        RECT 5.605 434.025 6.815 435.115 ;
        RECT 6.295 433.485 6.815 434.025 ;
        RECT 2910.045 433.950 2910.335 435.115 ;
        RECT 2912.805 434.025 2914.015 435.115 ;
        RECT 2912.805 433.485 2913.325 434.025 ;
        RECT 6.295 430.935 6.815 431.475 ;
        RECT 5.605 429.845 6.815 430.935 ;
        RECT 2912.805 430.935 2913.325 431.475 ;
        RECT 2912.805 429.845 2914.015 430.935 ;
        RECT 5.520 429.675 6.900 429.845 ;
        RECT 2909.960 429.675 2910.420 429.845 ;
        RECT 2912.720 429.675 2914.100 429.845 ;
        RECT 5.605 428.585 6.815 429.675 ;
        RECT 6.295 428.045 6.815 428.585 ;
        RECT 2910.045 428.510 2910.335 429.675 ;
        RECT 2912.805 428.585 2914.015 429.675 ;
        RECT 2912.805 428.045 2913.325 428.585 ;
        RECT 6.295 425.495 6.815 426.035 ;
        RECT 5.605 424.405 6.815 425.495 ;
        RECT 2912.805 425.495 2913.325 426.035 ;
        RECT 2912.805 424.405 2914.015 425.495 ;
        RECT 5.520 424.235 6.900 424.405 ;
        RECT 2909.960 424.235 2910.420 424.405 ;
        RECT 2912.720 424.235 2914.100 424.405 ;
        RECT 5.605 423.145 6.815 424.235 ;
        RECT 6.295 422.605 6.815 423.145 ;
        RECT 2910.045 423.070 2910.335 424.235 ;
        RECT 2912.805 423.145 2914.015 424.235 ;
        RECT 2912.805 422.605 2913.325 423.145 ;
        RECT 6.295 420.055 6.815 420.595 ;
        RECT 5.605 418.965 6.815 420.055 ;
        RECT 2912.805 420.055 2913.325 420.595 ;
        RECT 2912.805 418.965 2914.015 420.055 ;
        RECT 5.520 418.795 6.900 418.965 ;
        RECT 2909.960 418.795 2910.420 418.965 ;
        RECT 2912.720 418.795 2914.100 418.965 ;
        RECT 5.605 417.705 6.815 418.795 ;
        RECT 6.295 417.165 6.815 417.705 ;
        RECT 2910.045 417.630 2910.335 418.795 ;
        RECT 2912.805 417.705 2914.015 418.795 ;
        RECT 2912.805 417.165 2913.325 417.705 ;
        RECT 6.295 414.615 6.815 415.155 ;
        RECT 5.605 413.525 6.815 414.615 ;
        RECT 2912.805 414.615 2913.325 415.155 ;
        RECT 2912.805 413.525 2914.015 414.615 ;
        RECT 5.520 413.355 6.900 413.525 ;
        RECT 2909.960 413.355 2910.420 413.525 ;
        RECT 2912.720 413.355 2914.100 413.525 ;
        RECT 5.605 412.265 6.815 413.355 ;
        RECT 6.295 411.725 6.815 412.265 ;
        RECT 2910.045 412.190 2910.335 413.355 ;
        RECT 2912.805 412.265 2914.015 413.355 ;
        RECT 2912.805 411.725 2913.325 412.265 ;
        RECT 6.295 409.175 6.815 409.715 ;
        RECT 5.605 408.085 6.815 409.175 ;
        RECT 2912.805 409.175 2913.325 409.715 ;
        RECT 2912.805 408.085 2914.015 409.175 ;
        RECT 5.520 407.915 6.900 408.085 ;
        RECT 2909.960 407.915 2910.420 408.085 ;
        RECT 2912.720 407.915 2914.100 408.085 ;
        RECT 5.605 406.825 6.815 407.915 ;
        RECT 6.295 406.285 6.815 406.825 ;
        RECT 2910.045 406.750 2910.335 407.915 ;
        RECT 2912.805 406.825 2914.015 407.915 ;
        RECT 2912.805 406.285 2913.325 406.825 ;
        RECT 6.295 403.735 6.815 404.275 ;
        RECT 5.605 402.645 6.815 403.735 ;
        RECT 2912.805 403.735 2913.325 404.275 ;
        RECT 2912.805 402.645 2914.015 403.735 ;
        RECT 5.520 402.475 6.900 402.645 ;
        RECT 8.740 402.475 10.120 402.645 ;
        RECT 2909.960 402.475 2910.420 402.645 ;
        RECT 2912.720 402.475 2914.100 402.645 ;
        RECT 5.605 401.385 6.815 402.475 ;
        RECT 9.015 401.750 9.345 402.475 ;
        RECT 6.295 400.845 6.815 401.385 ;
        RECT 2910.045 401.310 2910.335 402.475 ;
        RECT 2912.805 401.385 2914.015 402.475 ;
        RECT 2912.805 400.845 2913.325 401.385 ;
        RECT 6.295 398.295 6.815 398.835 ;
        RECT 5.605 397.205 6.815 398.295 ;
        RECT 2912.805 398.295 2913.325 398.835 ;
        RECT 2912.805 397.205 2914.015 398.295 ;
        RECT 5.520 397.035 6.900 397.205 ;
        RECT 2909.960 397.035 2910.420 397.205 ;
        RECT 2912.720 397.035 2914.100 397.205 ;
        RECT 5.605 395.945 6.815 397.035 ;
        RECT 6.295 395.405 6.815 395.945 ;
        RECT 2910.045 395.870 2910.335 397.035 ;
        RECT 2912.805 395.945 2914.015 397.035 ;
        RECT 2912.805 395.405 2913.325 395.945 ;
        RECT 6.295 392.855 6.815 393.395 ;
        RECT 5.605 391.765 6.815 392.855 ;
        RECT 2912.805 392.855 2913.325 393.395 ;
        RECT 9.015 391.765 9.345 392.490 ;
        RECT 2912.805 391.765 2914.015 392.855 ;
        RECT 5.520 391.595 6.900 391.765 ;
        RECT 8.740 391.595 10.120 391.765 ;
        RECT 2909.960 391.595 2910.420 391.765 ;
        RECT 2912.720 391.595 2914.100 391.765 ;
        RECT 5.605 390.505 6.815 391.595 ;
        RECT 6.295 389.965 6.815 390.505 ;
        RECT 2910.045 390.430 2910.335 391.595 ;
        RECT 2912.805 390.505 2914.015 391.595 ;
        RECT 2912.805 389.965 2913.325 390.505 ;
        RECT 6.295 387.415 6.815 387.955 ;
        RECT 5.605 386.325 6.815 387.415 ;
        RECT 2912.805 387.415 2913.325 387.955 ;
        RECT 2912.805 386.325 2914.015 387.415 ;
        RECT 5.520 386.155 6.900 386.325 ;
        RECT 2909.960 386.155 2910.420 386.325 ;
        RECT 2912.720 386.155 2914.100 386.325 ;
        RECT 5.605 385.065 6.815 386.155 ;
        RECT 6.295 384.525 6.815 385.065 ;
        RECT 2910.045 384.990 2910.335 386.155 ;
        RECT 2912.805 385.065 2914.015 386.155 ;
        RECT 2912.805 384.525 2913.325 385.065 ;
        RECT 6.295 381.975 6.815 382.515 ;
        RECT 5.605 380.885 6.815 381.975 ;
        RECT 2912.805 381.975 2913.325 382.515 ;
        RECT 2912.805 380.885 2914.015 381.975 ;
        RECT 5.520 380.715 6.900 380.885 ;
        RECT 2909.960 380.715 2910.420 380.885 ;
        RECT 2912.720 380.715 2914.100 380.885 ;
        RECT 5.605 379.625 6.815 380.715 ;
        RECT 6.295 379.085 6.815 379.625 ;
        RECT 2910.045 379.550 2910.335 380.715 ;
        RECT 2912.805 379.625 2914.015 380.715 ;
        RECT 2912.805 379.085 2913.325 379.625 ;
        RECT 6.295 376.535 6.815 377.075 ;
        RECT 5.605 375.445 6.815 376.535 ;
        RECT 2912.805 376.535 2913.325 377.075 ;
        RECT 2912.805 375.445 2914.015 376.535 ;
        RECT 5.520 375.275 6.900 375.445 ;
        RECT 2909.960 375.275 2910.420 375.445 ;
        RECT 2912.720 375.275 2914.100 375.445 ;
        RECT 5.605 374.185 6.815 375.275 ;
        RECT 6.295 373.645 6.815 374.185 ;
        RECT 2910.045 374.110 2910.335 375.275 ;
        RECT 2912.805 374.185 2914.015 375.275 ;
        RECT 2912.805 373.645 2913.325 374.185 ;
        RECT 6.295 371.095 6.815 371.635 ;
        RECT 5.605 370.005 6.815 371.095 ;
        RECT 2912.805 371.095 2913.325 371.635 ;
        RECT 2912.805 370.005 2914.015 371.095 ;
        RECT 5.520 369.835 6.900 370.005 ;
        RECT 2909.960 369.835 2910.420 370.005 ;
        RECT 2912.720 369.835 2914.100 370.005 ;
        RECT 5.605 368.745 6.815 369.835 ;
        RECT 6.295 368.205 6.815 368.745 ;
        RECT 2910.045 368.670 2910.335 369.835 ;
        RECT 2912.805 368.745 2914.015 369.835 ;
        RECT 2912.805 368.205 2913.325 368.745 ;
        RECT 6.295 365.655 6.815 366.195 ;
        RECT 5.605 364.565 6.815 365.655 ;
        RECT 2912.805 365.655 2913.325 366.195 ;
        RECT 2912.805 364.565 2914.015 365.655 ;
        RECT 5.520 364.395 6.900 364.565 ;
        RECT 2909.960 364.395 2910.420 364.565 ;
        RECT 2912.720 364.395 2914.100 364.565 ;
        RECT 5.605 363.305 6.815 364.395 ;
        RECT 6.295 362.765 6.815 363.305 ;
        RECT 2910.045 363.230 2910.335 364.395 ;
        RECT 2912.805 363.305 2914.015 364.395 ;
        RECT 2912.805 362.765 2913.325 363.305 ;
        RECT 6.295 360.215 6.815 360.755 ;
        RECT 5.605 359.125 6.815 360.215 ;
        RECT 2912.805 360.215 2913.325 360.755 ;
        RECT 2912.805 359.125 2914.015 360.215 ;
        RECT 5.520 358.955 6.900 359.125 ;
        RECT 2909.960 358.955 2910.420 359.125 ;
        RECT 2912.720 358.955 2914.100 359.125 ;
        RECT 5.605 357.865 6.815 358.955 ;
        RECT 6.295 357.325 6.815 357.865 ;
        RECT 2910.045 357.790 2910.335 358.955 ;
        RECT 2912.805 357.865 2914.015 358.955 ;
        RECT 2912.805 357.325 2913.325 357.865 ;
        RECT 6.295 354.775 6.815 355.315 ;
        RECT 5.605 353.685 6.815 354.775 ;
        RECT 2912.805 354.775 2913.325 355.315 ;
        RECT 2912.805 353.685 2914.015 354.775 ;
        RECT 5.520 353.515 6.900 353.685 ;
        RECT 2909.960 353.515 2910.420 353.685 ;
        RECT 2912.720 353.515 2914.100 353.685 ;
        RECT 5.605 352.425 6.815 353.515 ;
        RECT 6.295 351.885 6.815 352.425 ;
        RECT 2910.045 352.350 2910.335 353.515 ;
        RECT 2912.805 352.425 2914.015 353.515 ;
        RECT 2912.805 351.885 2913.325 352.425 ;
        RECT 6.295 349.335 6.815 349.875 ;
        RECT 5.605 348.245 6.815 349.335 ;
        RECT 2912.805 349.335 2913.325 349.875 ;
        RECT 2912.805 348.245 2914.015 349.335 ;
        RECT 5.520 348.075 6.900 348.245 ;
        RECT 2909.960 348.075 2910.420 348.245 ;
        RECT 2912.720 348.075 2914.100 348.245 ;
        RECT 5.605 346.985 6.815 348.075 ;
        RECT 6.295 346.445 6.815 346.985 ;
        RECT 2910.045 346.910 2910.335 348.075 ;
        RECT 2912.805 346.985 2914.015 348.075 ;
        RECT 2912.805 346.445 2913.325 346.985 ;
        RECT 6.295 343.895 6.815 344.435 ;
        RECT 5.605 342.805 6.815 343.895 ;
        RECT 2912.805 343.895 2913.325 344.435 ;
        RECT 2912.805 342.805 2914.015 343.895 ;
        RECT 5.520 342.635 6.900 342.805 ;
        RECT 2909.960 342.635 2910.420 342.805 ;
        RECT 2912.720 342.635 2914.100 342.805 ;
        RECT 5.605 341.545 6.815 342.635 ;
        RECT 6.295 341.005 6.815 341.545 ;
        RECT 2910.045 341.470 2910.335 342.635 ;
        RECT 2912.805 341.545 2914.015 342.635 ;
        RECT 2912.805 341.005 2913.325 341.545 ;
        RECT 6.295 338.455 6.815 338.995 ;
        RECT 5.605 337.365 6.815 338.455 ;
        RECT 2912.805 338.455 2913.325 338.995 ;
        RECT 2912.805 337.365 2914.015 338.455 ;
        RECT 5.520 337.195 6.900 337.365 ;
        RECT 2909.960 337.195 2910.420 337.365 ;
        RECT 2912.720 337.195 2914.100 337.365 ;
        RECT 5.605 336.105 6.815 337.195 ;
        RECT 6.295 335.565 6.815 336.105 ;
        RECT 2910.045 336.030 2910.335 337.195 ;
        RECT 2912.805 336.105 2914.015 337.195 ;
        RECT 2912.805 335.565 2913.325 336.105 ;
        RECT 6.295 333.015 6.815 333.555 ;
        RECT 5.605 331.925 6.815 333.015 ;
        RECT 2912.805 333.015 2913.325 333.555 ;
        RECT 2912.805 331.925 2914.015 333.015 ;
        RECT 5.520 331.755 6.900 331.925 ;
        RECT 2909.960 331.755 2910.420 331.925 ;
        RECT 2912.720 331.755 2914.100 331.925 ;
        RECT 5.605 330.665 6.815 331.755 ;
        RECT 6.295 330.125 6.815 330.665 ;
        RECT 2910.045 330.590 2910.335 331.755 ;
        RECT 2912.805 330.665 2914.015 331.755 ;
        RECT 2912.805 330.125 2913.325 330.665 ;
        RECT 6.295 327.575 6.815 328.115 ;
        RECT 5.605 326.485 6.815 327.575 ;
        RECT 2912.805 327.575 2913.325 328.115 ;
        RECT 2912.805 326.485 2914.015 327.575 ;
        RECT 5.520 326.315 6.900 326.485 ;
        RECT 2909.960 326.315 2910.420 326.485 ;
        RECT 2912.720 326.315 2914.100 326.485 ;
        RECT 5.605 325.225 6.815 326.315 ;
        RECT 6.295 324.685 6.815 325.225 ;
        RECT 2910.045 325.150 2910.335 326.315 ;
        RECT 2912.805 325.225 2914.015 326.315 ;
        RECT 2912.805 324.685 2913.325 325.225 ;
        RECT 6.295 322.135 6.815 322.675 ;
        RECT 5.605 321.045 6.815 322.135 ;
        RECT 2912.805 322.135 2913.325 322.675 ;
        RECT 2912.805 321.045 2914.015 322.135 ;
        RECT 5.520 320.875 6.900 321.045 ;
        RECT 2909.960 320.875 2910.420 321.045 ;
        RECT 2912.720 320.875 2914.100 321.045 ;
        RECT 5.605 319.785 6.815 320.875 ;
        RECT 6.295 319.245 6.815 319.785 ;
        RECT 2910.045 319.710 2910.335 320.875 ;
        RECT 2912.805 319.785 2914.015 320.875 ;
        RECT 2912.805 319.245 2913.325 319.785 ;
        RECT 6.295 316.695 6.815 317.235 ;
        RECT 5.605 315.605 6.815 316.695 ;
        RECT 2912.805 316.695 2913.325 317.235 ;
        RECT 2912.805 315.605 2914.015 316.695 ;
        RECT 5.520 315.435 6.900 315.605 ;
        RECT 8.740 315.435 10.120 315.605 ;
        RECT 2909.960 315.435 2910.420 315.605 ;
        RECT 2912.720 315.435 2914.100 315.605 ;
        RECT 5.605 314.345 6.815 315.435 ;
        RECT 9.015 314.710 9.345 315.435 ;
        RECT 6.295 313.805 6.815 314.345 ;
        RECT 2910.045 314.270 2910.335 315.435 ;
        RECT 2912.805 314.345 2914.015 315.435 ;
        RECT 2912.805 313.805 2913.325 314.345 ;
        RECT 6.295 311.255 6.815 311.795 ;
        RECT 5.605 310.165 6.815 311.255 ;
        RECT 2912.805 311.255 2913.325 311.795 ;
        RECT 2912.805 310.165 2914.015 311.255 ;
        RECT 5.520 309.995 6.900 310.165 ;
        RECT 2909.960 309.995 2910.420 310.165 ;
        RECT 2912.720 309.995 2914.100 310.165 ;
        RECT 5.605 308.905 6.815 309.995 ;
        RECT 6.295 308.365 6.815 308.905 ;
        RECT 2910.045 308.830 2910.335 309.995 ;
        RECT 2912.805 308.905 2914.015 309.995 ;
        RECT 2912.805 308.365 2913.325 308.905 ;
        RECT 6.295 305.815 6.815 306.355 ;
        RECT 5.605 304.725 6.815 305.815 ;
        RECT 2912.805 305.815 2913.325 306.355 ;
        RECT 2912.805 304.725 2914.015 305.815 ;
        RECT 5.520 304.555 6.900 304.725 ;
        RECT 2909.960 304.555 2910.420 304.725 ;
        RECT 2912.720 304.555 2914.100 304.725 ;
        RECT 5.605 303.465 6.815 304.555 ;
        RECT 6.295 302.925 6.815 303.465 ;
        RECT 2910.045 303.390 2910.335 304.555 ;
        RECT 2912.805 303.465 2914.015 304.555 ;
        RECT 2912.805 302.925 2913.325 303.465 ;
        RECT 6.295 300.375 6.815 300.915 ;
        RECT 5.605 299.285 6.815 300.375 ;
        RECT 2912.805 300.375 2913.325 300.915 ;
        RECT 2912.805 299.285 2914.015 300.375 ;
        RECT 5.520 299.115 6.900 299.285 ;
        RECT 2909.960 299.115 2910.420 299.285 ;
        RECT 2912.720 299.115 2914.100 299.285 ;
        RECT 5.605 298.025 6.815 299.115 ;
        RECT 6.295 297.485 6.815 298.025 ;
        RECT 2910.045 297.950 2910.335 299.115 ;
        RECT 2912.805 298.025 2914.015 299.115 ;
        RECT 2912.805 297.485 2913.325 298.025 ;
        RECT 6.295 294.935 6.815 295.475 ;
        RECT 5.605 293.845 6.815 294.935 ;
        RECT 2912.805 294.935 2913.325 295.475 ;
        RECT 2912.805 293.845 2914.015 294.935 ;
        RECT 5.520 293.675 6.900 293.845 ;
        RECT 2909.960 293.675 2910.420 293.845 ;
        RECT 2912.720 293.675 2914.100 293.845 ;
        RECT 5.605 292.585 6.815 293.675 ;
        RECT 6.295 292.045 6.815 292.585 ;
        RECT 2910.045 292.510 2910.335 293.675 ;
        RECT 2912.805 292.585 2914.015 293.675 ;
        RECT 2912.805 292.045 2913.325 292.585 ;
        RECT 6.295 289.495 6.815 290.035 ;
        RECT 5.605 288.405 6.815 289.495 ;
        RECT 2912.805 289.495 2913.325 290.035 ;
        RECT 2909.315 288.405 2909.645 289.130 ;
        RECT 2912.805 288.405 2914.015 289.495 ;
        RECT 5.520 288.235 6.900 288.405 ;
        RECT 2909.040 288.235 2910.420 288.405 ;
        RECT 2912.720 288.235 2914.100 288.405 ;
        RECT 5.605 287.145 6.815 288.235 ;
        RECT 6.295 286.605 6.815 287.145 ;
        RECT 2910.045 287.070 2910.335 288.235 ;
        RECT 2912.805 287.145 2914.015 288.235 ;
        RECT 2912.805 286.605 2913.325 287.145 ;
        RECT 6.295 284.055 6.815 284.595 ;
        RECT 5.605 282.965 6.815 284.055 ;
        RECT 2912.805 284.055 2913.325 284.595 ;
        RECT 2912.805 282.965 2914.015 284.055 ;
        RECT 5.520 282.795 6.900 282.965 ;
        RECT 2909.960 282.795 2910.420 282.965 ;
        RECT 2912.720 282.795 2914.100 282.965 ;
        RECT 5.605 281.705 6.815 282.795 ;
        RECT 6.295 281.165 6.815 281.705 ;
        RECT 2910.045 281.630 2910.335 282.795 ;
        RECT 2912.805 281.705 2914.015 282.795 ;
        RECT 2912.805 281.165 2913.325 281.705 ;
        RECT 6.295 278.615 6.815 279.155 ;
        RECT 5.605 277.525 6.815 278.615 ;
        RECT 2912.805 278.615 2913.325 279.155 ;
        RECT 2912.805 277.525 2914.015 278.615 ;
        RECT 5.520 277.355 6.900 277.525 ;
        RECT 2909.960 277.355 2910.420 277.525 ;
        RECT 2912.720 277.355 2914.100 277.525 ;
        RECT 5.605 276.265 6.815 277.355 ;
        RECT 6.295 275.725 6.815 276.265 ;
        RECT 2910.045 276.190 2910.335 277.355 ;
        RECT 2912.805 276.265 2914.015 277.355 ;
        RECT 2912.805 275.725 2913.325 276.265 ;
        RECT 6.295 273.175 6.815 273.715 ;
        RECT 5.605 272.085 6.815 273.175 ;
        RECT 2912.805 273.175 2913.325 273.715 ;
        RECT 2912.805 272.085 2914.015 273.175 ;
        RECT 5.520 271.915 6.900 272.085 ;
        RECT 2909.960 271.915 2910.420 272.085 ;
        RECT 2912.720 271.915 2914.100 272.085 ;
        RECT 5.605 270.825 6.815 271.915 ;
        RECT 6.295 270.285 6.815 270.825 ;
        RECT 2910.045 270.750 2910.335 271.915 ;
        RECT 2912.805 270.825 2914.015 271.915 ;
        RECT 2912.805 270.285 2913.325 270.825 ;
        RECT 6.295 267.735 6.815 268.275 ;
        RECT 5.605 266.645 6.815 267.735 ;
        RECT 2912.805 267.735 2913.325 268.275 ;
        RECT 2912.805 266.645 2914.015 267.735 ;
        RECT 5.520 266.475 6.900 266.645 ;
        RECT 2909.960 266.475 2910.420 266.645 ;
        RECT 2912.720 266.475 2914.100 266.645 ;
        RECT 5.605 265.385 6.815 266.475 ;
        RECT 6.295 264.845 6.815 265.385 ;
        RECT 2910.045 265.310 2910.335 266.475 ;
        RECT 2912.805 265.385 2914.015 266.475 ;
        RECT 2912.805 264.845 2913.325 265.385 ;
        RECT 6.295 262.295 6.815 262.835 ;
        RECT 5.605 261.205 6.815 262.295 ;
        RECT 2912.805 262.295 2913.325 262.835 ;
        RECT 2912.805 261.205 2914.015 262.295 ;
        RECT 5.520 261.035 6.900 261.205 ;
        RECT 2909.960 261.035 2910.420 261.205 ;
        RECT 2912.720 261.035 2914.100 261.205 ;
        RECT 5.605 259.945 6.815 261.035 ;
        RECT 6.295 259.405 6.815 259.945 ;
        RECT 2910.045 259.870 2910.335 261.035 ;
        RECT 2912.805 259.945 2914.015 261.035 ;
        RECT 2912.805 259.405 2913.325 259.945 ;
        RECT 6.295 256.855 6.815 257.395 ;
        RECT 5.605 255.765 6.815 256.855 ;
        RECT 2912.805 256.855 2913.325 257.395 ;
        RECT 2912.805 255.765 2914.015 256.855 ;
        RECT 5.520 255.595 6.900 255.765 ;
        RECT 2909.960 255.595 2910.420 255.765 ;
        RECT 2912.720 255.595 2914.100 255.765 ;
        RECT 5.605 254.505 6.815 255.595 ;
        RECT 6.295 253.965 6.815 254.505 ;
        RECT 2910.045 254.430 2910.335 255.595 ;
        RECT 2912.805 254.505 2914.015 255.595 ;
        RECT 2912.805 253.965 2913.325 254.505 ;
        RECT 6.295 251.415 6.815 251.955 ;
        RECT 5.605 250.325 6.815 251.415 ;
        RECT 2912.805 251.415 2913.325 251.955 ;
        RECT 2912.805 250.325 2914.015 251.415 ;
        RECT 5.520 250.155 6.900 250.325 ;
        RECT 2909.960 250.155 2910.420 250.325 ;
        RECT 2912.720 250.155 2914.100 250.325 ;
        RECT 5.605 249.065 6.815 250.155 ;
        RECT 6.295 248.525 6.815 249.065 ;
        RECT 2910.045 248.990 2910.335 250.155 ;
        RECT 2912.805 249.065 2914.015 250.155 ;
        RECT 2912.805 248.525 2913.325 249.065 ;
        RECT 6.295 245.975 6.815 246.515 ;
        RECT 5.605 244.885 6.815 245.975 ;
        RECT 2912.805 245.975 2913.325 246.515 ;
        RECT 2912.805 244.885 2914.015 245.975 ;
        RECT 5.520 244.715 6.900 244.885 ;
        RECT 2909.960 244.715 2910.420 244.885 ;
        RECT 2912.720 244.715 2914.100 244.885 ;
        RECT 5.605 243.625 6.815 244.715 ;
        RECT 6.295 243.085 6.815 243.625 ;
        RECT 2910.045 243.550 2910.335 244.715 ;
        RECT 2912.805 243.625 2914.015 244.715 ;
        RECT 2912.805 243.085 2913.325 243.625 ;
        RECT 6.295 240.535 6.815 241.075 ;
        RECT 5.605 239.445 6.815 240.535 ;
        RECT 2912.805 240.535 2913.325 241.075 ;
        RECT 2912.805 239.445 2914.015 240.535 ;
        RECT 5.520 239.275 6.900 239.445 ;
        RECT 2909.960 239.275 2910.420 239.445 ;
        RECT 2912.720 239.275 2914.100 239.445 ;
        RECT 5.605 238.185 6.815 239.275 ;
        RECT 6.295 237.645 6.815 238.185 ;
        RECT 2910.045 238.110 2910.335 239.275 ;
        RECT 2912.805 238.185 2914.015 239.275 ;
        RECT 2912.805 237.645 2913.325 238.185 ;
        RECT 6.295 235.095 6.815 235.635 ;
        RECT 5.605 234.005 6.815 235.095 ;
        RECT 2912.805 235.095 2913.325 235.635 ;
        RECT 2912.805 234.005 2914.015 235.095 ;
        RECT 5.520 233.835 6.900 234.005 ;
        RECT 2909.960 233.835 2911.800 234.005 ;
        RECT 2912.720 233.835 2914.100 234.005 ;
        RECT 5.605 232.745 6.815 233.835 ;
        RECT 6.295 232.205 6.815 232.745 ;
        RECT 2910.045 232.670 2910.335 233.835 ;
        RECT 2910.695 233.110 2911.025 233.835 ;
        RECT 2912.805 232.745 2914.015 233.835 ;
        RECT 2912.805 232.205 2913.325 232.745 ;
        RECT 6.295 229.655 6.815 230.195 ;
        RECT 5.605 228.565 6.815 229.655 ;
        RECT 2912.805 229.655 2913.325 230.195 ;
        RECT 2912.805 228.565 2914.015 229.655 ;
        RECT 5.520 228.395 6.900 228.565 ;
        RECT 2909.960 228.395 2910.420 228.565 ;
        RECT 2912.720 228.395 2914.100 228.565 ;
        RECT 5.605 227.305 6.815 228.395 ;
        RECT 6.295 226.765 6.815 227.305 ;
        RECT 2910.045 227.230 2910.335 228.395 ;
        RECT 2912.805 227.305 2914.015 228.395 ;
        RECT 2912.805 226.765 2913.325 227.305 ;
        RECT 6.295 224.215 6.815 224.755 ;
        RECT 5.605 223.125 6.815 224.215 ;
        RECT 2912.805 224.215 2913.325 224.755 ;
        RECT 2912.805 223.125 2914.015 224.215 ;
        RECT 5.520 222.955 6.900 223.125 ;
        RECT 2909.960 222.955 2910.420 223.125 ;
        RECT 2912.720 222.955 2914.100 223.125 ;
        RECT 5.605 221.865 6.815 222.955 ;
        RECT 6.295 221.325 6.815 221.865 ;
        RECT 2910.045 221.790 2910.335 222.955 ;
        RECT 2912.805 221.865 2914.015 222.955 ;
        RECT 2912.805 221.325 2913.325 221.865 ;
        RECT 6.295 218.775 6.815 219.315 ;
        RECT 5.605 217.685 6.815 218.775 ;
        RECT 2912.805 218.775 2913.325 219.315 ;
        RECT 2912.805 217.685 2914.015 218.775 ;
        RECT 5.520 217.515 6.900 217.685 ;
        RECT 2909.960 217.515 2910.420 217.685 ;
        RECT 2912.720 217.515 2914.100 217.685 ;
        RECT 5.605 216.425 6.815 217.515 ;
        RECT 6.295 215.885 6.815 216.425 ;
        RECT 2910.045 216.350 2910.335 217.515 ;
        RECT 2912.805 216.425 2914.015 217.515 ;
        RECT 2912.805 215.885 2913.325 216.425 ;
        RECT 6.295 213.335 6.815 213.875 ;
        RECT 5.605 212.245 6.815 213.335 ;
        RECT 2912.805 213.335 2913.325 213.875 ;
        RECT 2912.805 212.245 2914.015 213.335 ;
        RECT 5.520 212.075 6.900 212.245 ;
        RECT 2909.960 212.075 2910.420 212.245 ;
        RECT 2912.720 212.075 2914.100 212.245 ;
        RECT 5.605 210.985 6.815 212.075 ;
        RECT 6.295 210.445 6.815 210.985 ;
        RECT 2910.045 210.910 2910.335 212.075 ;
        RECT 2912.805 210.985 2914.015 212.075 ;
        RECT 2912.805 210.445 2913.325 210.985 ;
        RECT 6.295 207.895 6.815 208.435 ;
        RECT 5.605 206.805 6.815 207.895 ;
        RECT 2912.805 207.895 2913.325 208.435 ;
        RECT 2912.805 206.805 2914.015 207.895 ;
        RECT 5.520 206.635 6.900 206.805 ;
        RECT 2909.960 206.635 2910.420 206.805 ;
        RECT 2912.720 206.635 2914.100 206.805 ;
        RECT 5.605 205.545 6.815 206.635 ;
        RECT 6.295 205.005 6.815 205.545 ;
        RECT 2910.045 205.470 2910.335 206.635 ;
        RECT 2912.805 205.545 2914.015 206.635 ;
        RECT 2912.805 205.005 2913.325 205.545 ;
        RECT 6.295 202.455 6.815 202.995 ;
        RECT 5.605 201.365 6.815 202.455 ;
        RECT 2912.805 202.455 2913.325 202.995 ;
        RECT 2912.805 201.365 2914.015 202.455 ;
        RECT 5.520 201.195 6.900 201.365 ;
        RECT 2909.960 201.195 2910.420 201.365 ;
        RECT 2912.720 201.195 2914.100 201.365 ;
        RECT 5.605 200.105 6.815 201.195 ;
        RECT 6.295 199.565 6.815 200.105 ;
        RECT 2910.045 200.030 2910.335 201.195 ;
        RECT 2912.805 200.105 2914.015 201.195 ;
        RECT 2912.805 199.565 2913.325 200.105 ;
        RECT 6.295 197.015 6.815 197.555 ;
        RECT 5.605 195.925 6.815 197.015 ;
        RECT 2912.805 197.015 2913.325 197.555 ;
        RECT 2912.805 195.925 2914.015 197.015 ;
        RECT 5.520 195.755 6.900 195.925 ;
        RECT 2909.960 195.755 2910.420 195.925 ;
        RECT 2912.720 195.755 2914.100 195.925 ;
        RECT 5.605 194.665 6.815 195.755 ;
        RECT 6.295 194.125 6.815 194.665 ;
        RECT 2910.045 194.590 2910.335 195.755 ;
        RECT 2912.805 194.665 2914.015 195.755 ;
        RECT 2912.805 194.125 2913.325 194.665 ;
        RECT 6.295 191.575 6.815 192.115 ;
        RECT 5.605 190.485 6.815 191.575 ;
        RECT 2912.805 191.575 2913.325 192.115 ;
        RECT 2912.805 190.485 2914.015 191.575 ;
        RECT 5.520 190.315 6.900 190.485 ;
        RECT 2909.960 190.315 2910.420 190.485 ;
        RECT 2912.720 190.315 2914.100 190.485 ;
        RECT 5.605 189.225 6.815 190.315 ;
        RECT 6.295 188.685 6.815 189.225 ;
        RECT 2910.045 189.150 2910.335 190.315 ;
        RECT 2912.805 189.225 2914.015 190.315 ;
        RECT 2912.805 188.685 2913.325 189.225 ;
        RECT 6.295 186.135 6.815 186.675 ;
        RECT 5.605 185.045 6.815 186.135 ;
        RECT 2912.805 186.135 2913.325 186.675 ;
        RECT 2912.805 185.045 2914.015 186.135 ;
        RECT 5.520 184.875 6.900 185.045 ;
        RECT 2909.960 184.875 2910.420 185.045 ;
        RECT 2912.720 184.875 2914.100 185.045 ;
        RECT 5.605 183.785 6.815 184.875 ;
        RECT 6.295 183.245 6.815 183.785 ;
        RECT 2910.045 183.710 2910.335 184.875 ;
        RECT 2912.805 183.785 2914.015 184.875 ;
        RECT 2912.805 183.245 2913.325 183.785 ;
        RECT 6.295 180.695 6.815 181.235 ;
        RECT 5.605 179.605 6.815 180.695 ;
        RECT 2912.805 180.695 2913.325 181.235 ;
        RECT 2912.805 179.605 2914.015 180.695 ;
        RECT 5.520 179.435 6.900 179.605 ;
        RECT 2909.960 179.435 2910.420 179.605 ;
        RECT 2912.720 179.435 2914.100 179.605 ;
        RECT 5.605 178.345 6.815 179.435 ;
        RECT 6.295 177.805 6.815 178.345 ;
        RECT 2910.045 178.270 2910.335 179.435 ;
        RECT 2912.805 178.345 2914.015 179.435 ;
        RECT 2912.805 177.805 2913.325 178.345 ;
        RECT 6.295 175.255 6.815 175.795 ;
        RECT 5.605 174.165 6.815 175.255 ;
        RECT 2912.805 175.255 2913.325 175.795 ;
        RECT 2912.805 174.165 2914.015 175.255 ;
        RECT 5.520 173.995 6.900 174.165 ;
        RECT 2909.960 173.995 2910.420 174.165 ;
        RECT 2912.720 173.995 2914.100 174.165 ;
        RECT 5.605 172.905 6.815 173.995 ;
        RECT 6.295 172.365 6.815 172.905 ;
        RECT 2910.045 172.830 2910.335 173.995 ;
        RECT 2912.805 172.905 2914.015 173.995 ;
        RECT 2912.805 172.365 2913.325 172.905 ;
        RECT 6.295 169.815 6.815 170.355 ;
        RECT 5.605 168.725 6.815 169.815 ;
        RECT 2912.805 169.815 2913.325 170.355 ;
        RECT 2912.805 168.725 2914.015 169.815 ;
        RECT 5.520 168.555 6.900 168.725 ;
        RECT 2909.960 168.555 2910.420 168.725 ;
        RECT 2912.720 168.555 2914.100 168.725 ;
        RECT 5.605 167.465 6.815 168.555 ;
        RECT 6.295 166.925 6.815 167.465 ;
        RECT 2910.045 167.390 2910.335 168.555 ;
        RECT 2912.805 167.465 2914.015 168.555 ;
        RECT 2912.805 166.925 2913.325 167.465 ;
        RECT 6.295 164.375 6.815 164.915 ;
        RECT 5.605 163.285 6.815 164.375 ;
        RECT 2912.805 164.375 2913.325 164.915 ;
        RECT 2912.805 163.285 2914.015 164.375 ;
        RECT 5.520 163.115 6.900 163.285 ;
        RECT 2909.960 163.115 2910.420 163.285 ;
        RECT 2912.720 163.115 2914.100 163.285 ;
        RECT 5.605 162.025 6.815 163.115 ;
        RECT 6.295 161.485 6.815 162.025 ;
        RECT 2910.045 161.950 2910.335 163.115 ;
        RECT 2912.805 162.025 2914.015 163.115 ;
        RECT 2912.805 161.485 2913.325 162.025 ;
        RECT 6.295 158.935 6.815 159.475 ;
        RECT 5.605 157.845 6.815 158.935 ;
        RECT 2912.805 158.935 2913.325 159.475 ;
        RECT 2912.805 157.845 2914.015 158.935 ;
        RECT 5.520 157.675 6.900 157.845 ;
        RECT 2909.960 157.675 2910.420 157.845 ;
        RECT 2912.720 157.675 2914.100 157.845 ;
        RECT 5.605 156.585 6.815 157.675 ;
        RECT 6.295 156.045 6.815 156.585 ;
        RECT 2910.045 156.510 2910.335 157.675 ;
        RECT 2912.805 156.585 2914.015 157.675 ;
        RECT 2912.805 156.045 2913.325 156.585 ;
        RECT 6.295 153.495 6.815 154.035 ;
        RECT 5.605 152.405 6.815 153.495 ;
        RECT 2912.805 153.495 2913.325 154.035 ;
        RECT 2912.805 152.405 2914.015 153.495 ;
        RECT 5.520 152.235 6.900 152.405 ;
        RECT 2909.960 152.235 2910.420 152.405 ;
        RECT 2912.720 152.235 2914.100 152.405 ;
        RECT 5.605 151.145 6.815 152.235 ;
        RECT 6.295 150.605 6.815 151.145 ;
        RECT 2910.045 151.070 2910.335 152.235 ;
        RECT 2912.805 151.145 2914.015 152.235 ;
        RECT 2912.805 150.605 2913.325 151.145 ;
        RECT 6.295 148.055 6.815 148.595 ;
        RECT 5.605 146.965 6.815 148.055 ;
        RECT 2912.805 148.055 2913.325 148.595 ;
        RECT 2912.805 146.965 2914.015 148.055 ;
        RECT 5.520 146.795 6.900 146.965 ;
        RECT 2909.960 146.795 2910.420 146.965 ;
        RECT 2912.720 146.795 2914.100 146.965 ;
        RECT 5.605 145.705 6.815 146.795 ;
        RECT 6.295 145.165 6.815 145.705 ;
        RECT 2910.045 145.630 2910.335 146.795 ;
        RECT 2912.805 145.705 2914.015 146.795 ;
        RECT 2912.805 145.165 2913.325 145.705 ;
        RECT 6.295 142.615 6.815 143.155 ;
        RECT 5.605 141.525 6.815 142.615 ;
        RECT 2912.805 142.615 2913.325 143.155 ;
        RECT 2912.805 141.525 2914.015 142.615 ;
        RECT 5.520 141.355 6.900 141.525 ;
        RECT 2909.960 141.355 2910.420 141.525 ;
        RECT 2912.720 141.355 2914.100 141.525 ;
        RECT 5.605 140.265 6.815 141.355 ;
        RECT 6.295 139.725 6.815 140.265 ;
        RECT 2910.045 140.190 2910.335 141.355 ;
        RECT 2912.805 140.265 2914.015 141.355 ;
        RECT 2912.805 139.725 2913.325 140.265 ;
        RECT 6.295 137.175 6.815 137.715 ;
        RECT 5.605 136.085 6.815 137.175 ;
        RECT 2912.805 137.175 2913.325 137.715 ;
        RECT 2912.805 136.085 2914.015 137.175 ;
        RECT 5.520 135.915 6.900 136.085 ;
        RECT 2909.960 135.915 2910.420 136.085 ;
        RECT 2912.720 135.915 2914.100 136.085 ;
        RECT 5.605 134.825 6.815 135.915 ;
        RECT 6.295 134.285 6.815 134.825 ;
        RECT 2910.045 134.750 2910.335 135.915 ;
        RECT 2912.805 134.825 2914.015 135.915 ;
        RECT 2912.805 134.285 2913.325 134.825 ;
        RECT 6.295 131.735 6.815 132.275 ;
        RECT 5.605 130.645 6.815 131.735 ;
        RECT 2912.805 131.735 2913.325 132.275 ;
        RECT 2912.805 130.645 2914.015 131.735 ;
        RECT 5.520 130.475 6.900 130.645 ;
        RECT 2909.960 130.475 2910.420 130.645 ;
        RECT 2912.720 130.475 2914.100 130.645 ;
        RECT 5.605 129.385 6.815 130.475 ;
        RECT 6.295 128.845 6.815 129.385 ;
        RECT 2910.045 129.310 2910.335 130.475 ;
        RECT 2912.805 129.385 2914.015 130.475 ;
        RECT 2912.805 128.845 2913.325 129.385 ;
        RECT 6.295 126.295 6.815 126.835 ;
        RECT 5.605 125.205 6.815 126.295 ;
        RECT 2912.805 126.295 2913.325 126.835 ;
        RECT 7.415 125.205 7.745 125.705 ;
        RECT 8.340 125.205 8.605 125.665 ;
        RECT 10.510 125.205 10.680 126.005 ;
        RECT 12.390 125.205 12.605 125.705 ;
        RECT 13.525 125.205 13.700 125.985 ;
        RECT 2912.805 125.205 2914.015 126.295 ;
        RECT 5.520 125.035 13.700 125.205 ;
        RECT 2909.960 125.035 2910.420 125.205 ;
        RECT 2912.720 125.035 2914.100 125.205 ;
        RECT 5.605 123.945 6.815 125.035 ;
        RECT 6.295 123.405 6.815 123.945 ;
        RECT 2910.045 123.870 2910.335 125.035 ;
        RECT 2912.805 123.945 2914.015 125.035 ;
        RECT 2912.805 123.405 2913.325 123.945 ;
        RECT 6.295 120.855 6.815 121.395 ;
        RECT 5.605 119.765 6.815 120.855 ;
        RECT 2912.805 120.855 2913.325 121.395 ;
        RECT 2912.805 119.765 2914.015 120.855 ;
        RECT 5.520 119.595 6.900 119.765 ;
        RECT 2909.960 119.595 2910.420 119.765 ;
        RECT 2912.720 119.595 2914.100 119.765 ;
        RECT 5.605 118.505 6.815 119.595 ;
        RECT 6.295 117.965 6.815 118.505 ;
        RECT 2910.045 118.430 2910.335 119.595 ;
        RECT 2912.805 118.505 2914.015 119.595 ;
        RECT 2912.805 117.965 2913.325 118.505 ;
        RECT 6.295 115.415 6.815 115.955 ;
        RECT 5.605 114.325 6.815 115.415 ;
        RECT 2912.805 115.415 2913.325 115.955 ;
        RECT 2912.805 114.325 2914.015 115.415 ;
        RECT 5.520 114.155 6.900 114.325 ;
        RECT 2909.960 114.155 2910.420 114.325 ;
        RECT 2912.720 114.155 2914.100 114.325 ;
        RECT 5.605 113.065 6.815 114.155 ;
        RECT 6.295 112.525 6.815 113.065 ;
        RECT 2910.045 112.990 2910.335 114.155 ;
        RECT 2912.805 113.065 2914.015 114.155 ;
        RECT 2912.805 112.525 2913.325 113.065 ;
        RECT 6.295 109.975 6.815 110.515 ;
        RECT 5.605 108.885 6.815 109.975 ;
        RECT 2912.805 109.975 2913.325 110.515 ;
        RECT 2912.805 108.885 2914.015 109.975 ;
        RECT 5.520 108.715 6.900 108.885 ;
        RECT 2909.960 108.715 2910.420 108.885 ;
        RECT 2912.720 108.715 2914.100 108.885 ;
        RECT 5.605 107.625 6.815 108.715 ;
        RECT 6.295 107.085 6.815 107.625 ;
        RECT 2910.045 107.550 2910.335 108.715 ;
        RECT 2912.805 107.625 2914.015 108.715 ;
        RECT 2912.805 107.085 2913.325 107.625 ;
        RECT 6.295 104.535 6.815 105.075 ;
        RECT 5.605 103.445 6.815 104.535 ;
        RECT 8.865 103.445 9.095 104.585 ;
        RECT 9.765 103.445 9.975 104.585 ;
        RECT 2912.805 104.535 2913.325 105.075 ;
        RECT 2912.805 103.445 2914.015 104.535 ;
        RECT 5.520 103.275 6.900 103.445 ;
        RECT 8.740 103.275 10.120 103.445 ;
        RECT 2909.960 103.275 2910.420 103.445 ;
        RECT 2912.720 103.275 2914.100 103.445 ;
        RECT 5.605 102.185 6.815 103.275 ;
        RECT 6.295 101.645 6.815 102.185 ;
        RECT 2910.045 102.110 2910.335 103.275 ;
        RECT 2912.805 102.185 2914.015 103.275 ;
        RECT 2912.805 101.645 2913.325 102.185 ;
        RECT 6.295 99.095 6.815 99.635 ;
        RECT 5.605 98.005 6.815 99.095 ;
        RECT 2912.805 99.095 2913.325 99.635 ;
        RECT 2912.805 98.005 2914.015 99.095 ;
        RECT 5.520 97.835 6.900 98.005 ;
        RECT 2909.960 97.835 2910.420 98.005 ;
        RECT 2912.720 97.835 2914.100 98.005 ;
        RECT 5.605 96.745 6.815 97.835 ;
        RECT 6.295 96.205 6.815 96.745 ;
        RECT 2910.045 96.670 2910.335 97.835 ;
        RECT 2912.805 96.745 2914.015 97.835 ;
        RECT 2912.805 96.205 2913.325 96.745 ;
        RECT 6.295 93.655 6.815 94.195 ;
        RECT 5.605 92.565 6.815 93.655 ;
        RECT 2912.805 93.655 2913.325 94.195 ;
        RECT 2912.805 92.565 2914.015 93.655 ;
        RECT 5.520 92.395 6.900 92.565 ;
        RECT 2909.960 92.395 2910.420 92.565 ;
        RECT 2912.720 92.395 2914.100 92.565 ;
        RECT 5.605 91.305 6.815 92.395 ;
        RECT 6.295 90.765 6.815 91.305 ;
        RECT 2910.045 91.230 2910.335 92.395 ;
        RECT 2912.805 91.305 2914.015 92.395 ;
        RECT 2912.805 90.765 2913.325 91.305 ;
        RECT 6.295 88.215 6.815 88.755 ;
        RECT 5.605 87.125 6.815 88.215 ;
        RECT 2912.805 88.215 2913.325 88.755 ;
        RECT 2912.805 87.125 2914.015 88.215 ;
        RECT 5.520 86.955 6.900 87.125 ;
        RECT 2909.960 86.955 2910.420 87.125 ;
        RECT 2912.720 86.955 2914.100 87.125 ;
        RECT 5.605 85.865 6.815 86.955 ;
        RECT 6.295 85.325 6.815 85.865 ;
        RECT 2910.045 85.790 2910.335 86.955 ;
        RECT 2912.805 85.865 2914.015 86.955 ;
        RECT 2912.805 85.325 2913.325 85.865 ;
        RECT 6.295 82.775 6.815 83.315 ;
        RECT 5.605 81.685 6.815 82.775 ;
        RECT 2912.805 82.775 2913.325 83.315 ;
        RECT 2912.805 81.685 2914.015 82.775 ;
        RECT 5.520 81.515 6.900 81.685 ;
        RECT 2909.960 81.515 2910.420 81.685 ;
        RECT 2912.720 81.515 2914.100 81.685 ;
        RECT 5.605 80.425 6.815 81.515 ;
        RECT 6.295 79.885 6.815 80.425 ;
        RECT 2910.045 80.350 2910.335 81.515 ;
        RECT 2912.805 80.425 2914.015 81.515 ;
        RECT 2912.805 79.885 2913.325 80.425 ;
        RECT 6.295 77.335 6.815 77.875 ;
        RECT 5.605 76.245 6.815 77.335 ;
        RECT 2912.805 77.335 2913.325 77.875 ;
        RECT 2912.805 76.245 2914.015 77.335 ;
        RECT 5.520 76.075 6.900 76.245 ;
        RECT 2909.960 76.075 2910.420 76.245 ;
        RECT 2912.720 76.075 2914.100 76.245 ;
        RECT 5.605 74.985 6.815 76.075 ;
        RECT 6.295 74.445 6.815 74.985 ;
        RECT 2910.045 74.910 2910.335 76.075 ;
        RECT 2912.805 74.985 2914.015 76.075 ;
        RECT 2912.805 74.445 2913.325 74.985 ;
        RECT 6.295 71.895 6.815 72.435 ;
        RECT 5.605 70.805 6.815 71.895 ;
        RECT 2912.805 71.895 2913.325 72.435 ;
        RECT 2912.805 70.805 2914.015 71.895 ;
        RECT 5.520 70.635 6.900 70.805 ;
        RECT 2909.960 70.635 2910.420 70.805 ;
        RECT 2912.720 70.635 2914.100 70.805 ;
        RECT 5.605 69.545 6.815 70.635 ;
        RECT 6.295 69.005 6.815 69.545 ;
        RECT 2910.045 69.470 2910.335 70.635 ;
        RECT 2912.805 69.545 2914.015 70.635 ;
        RECT 2912.805 69.005 2913.325 69.545 ;
        RECT 6.295 66.455 6.815 66.995 ;
        RECT 5.605 65.365 6.815 66.455 ;
        RECT 2912.805 66.455 2913.325 66.995 ;
        RECT 2912.805 65.365 2914.015 66.455 ;
        RECT 5.520 65.195 6.900 65.365 ;
        RECT 2909.960 65.195 2910.420 65.365 ;
        RECT 2912.720 65.195 2914.100 65.365 ;
        RECT 5.605 64.105 6.815 65.195 ;
        RECT 6.295 63.565 6.815 64.105 ;
        RECT 2910.045 64.030 2910.335 65.195 ;
        RECT 2912.805 64.105 2914.015 65.195 ;
        RECT 2912.805 63.565 2913.325 64.105 ;
        RECT 6.295 61.015 6.815 61.555 ;
        RECT 5.605 59.925 6.815 61.015 ;
        RECT 2912.805 61.015 2913.325 61.555 ;
        RECT 2909.315 59.925 2909.645 60.650 ;
        RECT 2912.805 59.925 2914.015 61.015 ;
        RECT 5.520 59.755 6.900 59.925 ;
        RECT 2909.040 59.755 2910.420 59.925 ;
        RECT 2912.720 59.755 2914.100 59.925 ;
        RECT 5.605 58.665 6.815 59.755 ;
        RECT 6.295 58.125 6.815 58.665 ;
        RECT 2910.045 58.590 2910.335 59.755 ;
        RECT 2912.805 58.665 2914.015 59.755 ;
        RECT 2912.805 58.125 2913.325 58.665 ;
        RECT 6.295 55.575 6.815 56.115 ;
        RECT 5.605 54.485 6.815 55.575 ;
        RECT 2912.805 55.575 2913.325 56.115 ;
        RECT 2912.805 54.485 2914.015 55.575 ;
        RECT 5.520 54.315 6.900 54.485 ;
        RECT 2909.960 54.315 2910.420 54.485 ;
        RECT 2912.720 54.315 2914.100 54.485 ;
        RECT 5.605 53.225 6.815 54.315 ;
        RECT 6.295 52.685 6.815 53.225 ;
        RECT 2910.045 53.150 2910.335 54.315 ;
        RECT 2912.805 53.225 2914.015 54.315 ;
        RECT 2912.805 52.685 2913.325 53.225 ;
        RECT 6.295 50.135 6.815 50.675 ;
        RECT 5.605 49.045 6.815 50.135 ;
        RECT 2912.805 50.135 2913.325 50.675 ;
        RECT 2912.805 49.045 2914.015 50.135 ;
        RECT 5.520 48.875 6.900 49.045 ;
        RECT 2909.960 48.875 2910.420 49.045 ;
        RECT 2912.720 48.875 2914.100 49.045 ;
        RECT 5.605 47.785 6.815 48.875 ;
        RECT 6.295 47.245 6.815 47.785 ;
        RECT 2910.045 47.710 2910.335 48.875 ;
        RECT 2912.805 47.785 2914.015 48.875 ;
        RECT 2912.805 47.245 2913.325 47.785 ;
        RECT 6.295 44.695 6.815 45.235 ;
        RECT 5.605 43.605 6.815 44.695 ;
        RECT 2912.805 44.695 2913.325 45.235 ;
        RECT 2912.805 43.605 2914.015 44.695 ;
        RECT 5.520 43.435 13.700 43.605 ;
        RECT 2909.960 43.435 2910.420 43.605 ;
        RECT 2912.720 43.435 2914.100 43.605 ;
        RECT 5.605 42.345 6.815 43.435 ;
        RECT 7.415 42.935 7.745 43.435 ;
        RECT 8.340 42.975 8.605 43.435 ;
        RECT 10.510 42.635 10.680 43.435 ;
        RECT 12.390 42.935 12.605 43.435 ;
        RECT 13.525 42.655 13.700 43.435 ;
        RECT 6.295 41.805 6.815 42.345 ;
        RECT 2910.045 42.270 2910.335 43.435 ;
        RECT 2912.805 42.345 2914.015 43.435 ;
        RECT 2912.805 41.805 2913.325 42.345 ;
        RECT 6.295 39.255 6.815 39.795 ;
        RECT 5.605 38.165 6.815 39.255 ;
        RECT 2912.805 39.255 2913.325 39.795 ;
        RECT 2912.805 38.165 2914.015 39.255 ;
        RECT 5.520 37.995 6.900 38.165 ;
        RECT 2909.960 37.995 2910.420 38.165 ;
        RECT 2912.720 37.995 2914.100 38.165 ;
        RECT 5.605 36.905 6.815 37.995 ;
        RECT 6.295 36.365 6.815 36.905 ;
        RECT 2910.045 36.830 2910.335 37.995 ;
        RECT 2912.805 36.905 2914.015 37.995 ;
        RECT 2912.805 36.365 2913.325 36.905 ;
        RECT 6.295 33.815 6.815 34.355 ;
        RECT 5.605 32.725 6.815 33.815 ;
        RECT 2912.805 33.815 2913.325 34.355 ;
        RECT 2912.805 32.725 2914.015 33.815 ;
        RECT 5.520 32.555 6.900 32.725 ;
        RECT 2909.960 32.555 2910.420 32.725 ;
        RECT 2912.720 32.555 2914.100 32.725 ;
        RECT 5.605 31.465 6.815 32.555 ;
        RECT 6.295 30.925 6.815 31.465 ;
        RECT 2910.045 31.390 2910.335 32.555 ;
        RECT 2912.805 31.465 2914.015 32.555 ;
        RECT 2912.805 30.925 2913.325 31.465 ;
        RECT 6.295 28.375 6.815 28.915 ;
        RECT 5.605 27.285 6.815 28.375 ;
        RECT 2912.805 28.375 2913.325 28.915 ;
        RECT 2912.805 27.285 2914.015 28.375 ;
        RECT 5.520 27.115 6.900 27.285 ;
        RECT 2909.960 27.115 2910.420 27.285 ;
        RECT 2912.720 27.115 2914.100 27.285 ;
        RECT 5.605 26.025 6.815 27.115 ;
        RECT 6.295 25.485 6.815 26.025 ;
        RECT 2910.045 25.950 2910.335 27.115 ;
        RECT 2912.805 26.025 2914.015 27.115 ;
        RECT 2912.805 25.485 2913.325 26.025 ;
        RECT 6.295 22.935 6.815 23.475 ;
        RECT 5.605 21.845 6.815 22.935 ;
        RECT 2912.805 22.935 2913.325 23.475 ;
        RECT 2912.805 21.845 2914.015 22.935 ;
        RECT 5.520 21.675 13.700 21.845 ;
        RECT 2909.960 21.675 2910.420 21.845 ;
        RECT 2912.720 21.675 2914.100 21.845 ;
        RECT 5.605 20.585 6.815 21.675 ;
        RECT 7.455 21.165 7.705 21.675 ;
        RECT 8.295 21.165 8.545 21.675 ;
        RECT 10.075 21.175 10.325 21.675 ;
        RECT 11.755 20.835 12.005 21.675 ;
        RECT 12.595 21.205 12.845 21.675 ;
        RECT 13.435 20.865 13.685 21.675 ;
        RECT 6.295 20.045 6.815 20.585 ;
        RECT 2910.045 20.510 2910.335 21.675 ;
        RECT 2912.805 20.585 2914.015 21.675 ;
        RECT 2912.805 20.045 2913.325 20.585 ;
        RECT 6.295 17.495 6.815 18.035 ;
        RECT 5.605 16.405 6.815 17.495 ;
        RECT 2912.805 17.495 2913.325 18.035 ;
        RECT 7.415 16.405 7.745 16.905 ;
        RECT 8.340 16.405 8.605 16.865 ;
        RECT 10.510 16.405 10.680 17.205 ;
        RECT 12.390 16.405 12.605 16.905 ;
        RECT 13.525 16.405 13.700 17.185 ;
        RECT 2909.315 16.405 2909.645 17.130 ;
        RECT 2910.695 16.405 2911.025 17.130 ;
        RECT 2912.805 16.405 2914.015 17.495 ;
        RECT 5.520 16.235 13.700 16.405 ;
        RECT 2907.200 16.235 2911.800 16.405 ;
        RECT 2912.720 16.235 2914.100 16.405 ;
        RECT 5.605 15.145 6.815 16.235 ;
        RECT 7.415 15.735 7.745 16.235 ;
        RECT 8.340 15.775 8.605 16.235 ;
        RECT 10.510 15.435 10.680 16.235 ;
        RECT 12.390 15.735 12.605 16.235 ;
        RECT 13.525 15.455 13.700 16.235 ;
        RECT 2907.475 15.510 2907.805 16.235 ;
        RECT 2908.855 15.510 2909.185 16.235 ;
        RECT 6.295 14.605 6.815 15.145 ;
        RECT 2910.045 15.070 2910.335 16.235 ;
        RECT 2910.695 15.510 2911.025 16.235 ;
        RECT 2912.805 15.145 2914.015 16.235 ;
        RECT 2912.805 14.605 2913.325 15.145 ;
        RECT 6.295 12.055 6.815 12.595 ;
        RECT 5.605 10.965 6.815 12.055 ;
        RECT 8.865 10.965 9.095 12.105 ;
        RECT 9.765 10.965 9.975 12.105 ;
        RECT 10.395 10.965 10.725 11.690 ;
        RECT 19.865 10.965 20.155 12.130 ;
        RECT 34.125 10.965 34.415 12.130 ;
        RECT 48.385 10.965 48.675 12.130 ;
        RECT 62.645 10.965 62.935 12.130 ;
        RECT 76.905 10.965 77.195 12.130 ;
        RECT 82.395 10.965 82.725 11.465 ;
        RECT 83.320 10.965 83.585 11.425 ;
        RECT 85.490 10.965 85.660 11.765 ;
        RECT 87.370 10.965 87.585 11.465 ;
        RECT 88.505 10.965 88.685 11.745 ;
        RECT 89.380 10.965 89.550 11.795 ;
        RECT 90.220 10.965 90.390 11.795 ;
        RECT 91.165 10.965 91.455 12.130 ;
        RECT 105.425 10.965 105.715 12.130 ;
        RECT 119.685 10.965 119.975 12.130 ;
        RECT 133.945 10.965 134.235 12.130 ;
        RECT 148.205 10.965 148.495 12.130 ;
        RECT 162.465 10.965 162.755 12.130 ;
        RECT 176.725 10.965 177.015 12.130 ;
        RECT 190.985 10.965 191.275 12.130 ;
        RECT 205.245 10.965 205.535 12.130 ;
        RECT 206.175 10.965 206.425 11.475 ;
        RECT 207.015 10.965 207.265 11.475 ;
        RECT 208.795 10.965 209.045 11.465 ;
        RECT 210.475 10.965 210.725 11.805 ;
        RECT 211.315 10.965 211.565 11.435 ;
        RECT 212.155 10.965 212.405 11.775 ;
        RECT 219.505 10.965 219.795 12.130 ;
        RECT 225.620 10.965 225.870 11.775 ;
        RECT 226.460 10.965 226.710 11.805 ;
        RECT 227.300 10.965 228.070 11.475 ;
        RECT 229.500 10.965 229.830 11.475 ;
        RECT 231.305 10.965 231.510 12.145 ;
        RECT 233.765 10.965 234.055 12.130 ;
        RECT 241.015 10.965 241.465 11.665 ;
        RECT 242.030 10.965 242.360 11.665 ;
        RECT 242.930 10.965 243.260 11.665 ;
        RECT 243.790 10.965 244.120 11.665 ;
        RECT 248.025 10.965 248.315 12.130 ;
        RECT 262.285 10.965 262.575 12.130 ;
        RECT 262.880 10.965 263.130 11.775 ;
        RECT 263.720 10.965 263.970 11.805 ;
        RECT 264.560 10.965 265.330 11.475 ;
        RECT 266.760 10.965 267.090 11.475 ;
        RECT 268.565 10.965 268.770 12.145 ;
        RECT 276.545 10.965 276.835 12.130 ;
        RECT 290.805 10.965 291.095 12.130 ;
        RECT 305.065 10.965 305.355 12.130 ;
        RECT 319.325 10.965 319.615 12.130 ;
        RECT 333.585 10.965 333.875 12.130 ;
        RECT 347.845 10.965 348.135 12.130 ;
        RECT 352.485 10.965 352.715 12.105 ;
        RECT 353.385 10.965 353.595 12.105 ;
        RECT 362.105 10.965 362.395 12.130 ;
        RECT 376.365 10.965 376.655 12.130 ;
        RECT 390.625 10.965 390.915 12.130 ;
        RECT 391.515 10.965 391.845 11.465 ;
        RECT 392.440 10.965 392.705 11.425 ;
        RECT 394.610 10.965 394.780 11.765 ;
        RECT 396.490 10.965 396.705 11.465 ;
        RECT 397.625 10.965 397.805 11.745 ;
        RECT 398.500 10.965 398.670 11.795 ;
        RECT 399.340 10.965 399.510 11.795 ;
        RECT 399.865 10.965 400.095 12.105 ;
        RECT 400.765 10.965 400.975 12.105 ;
        RECT 404.885 10.965 405.175 12.130 ;
        RECT 419.145 10.965 419.435 12.130 ;
        RECT 433.405 10.965 433.695 12.130 ;
        RECT 447.665 10.965 447.955 12.130 ;
        RECT 451.020 10.965 451.270 11.775 ;
        RECT 451.860 10.965 452.110 11.805 ;
        RECT 452.700 10.965 453.470 11.475 ;
        RECT 454.900 10.965 455.230 11.475 ;
        RECT 456.705 10.965 456.910 12.145 ;
        RECT 461.925 10.965 462.215 12.130 ;
        RECT 476.185 10.965 476.475 12.130 ;
        RECT 490.445 10.965 490.735 12.130 ;
        RECT 504.705 10.965 504.995 12.130 ;
        RECT 518.965 10.965 519.255 12.130 ;
        RECT 533.225 10.965 533.515 12.130 ;
        RECT 547.485 10.965 547.775 12.130 ;
        RECT 561.745 10.965 562.035 12.130 ;
        RECT 576.005 10.965 576.295 12.130 ;
        RECT 590.265 10.965 590.555 12.130 ;
        RECT 604.525 10.965 604.815 12.130 ;
        RECT 618.785 10.965 619.075 12.130 ;
        RECT 633.045 10.965 633.335 12.130 ;
        RECT 647.305 10.965 647.595 12.130 ;
        RECT 661.565 10.965 661.855 12.130 ;
        RECT 675.825 10.965 676.115 12.130 ;
        RECT 690.085 10.965 690.375 12.130 ;
        RECT 704.345 10.965 704.635 12.130 ;
        RECT 718.605 10.965 718.895 12.130 ;
        RECT 732.865 10.965 733.155 12.130 ;
        RECT 747.125 10.965 747.415 12.130 ;
        RECT 761.385 10.965 761.675 12.130 ;
        RECT 775.645 10.965 775.935 12.130 ;
        RECT 789.905 10.965 790.195 12.130 ;
        RECT 804.165 10.965 804.455 12.130 ;
        RECT 818.425 10.965 818.715 12.130 ;
        RECT 832.685 10.965 832.975 12.130 ;
        RECT 846.945 10.965 847.235 12.130 ;
        RECT 861.205 10.965 861.495 12.130 ;
        RECT 875.465 10.965 875.755 12.130 ;
        RECT 889.725 10.965 890.015 12.130 ;
        RECT 903.985 10.965 904.275 12.130 ;
        RECT 918.245 10.965 918.535 12.130 ;
        RECT 932.505 10.965 932.795 12.130 ;
        RECT 946.765 10.965 947.055 12.130 ;
        RECT 961.025 10.965 961.315 12.130 ;
        RECT 975.285 10.965 975.575 12.130 ;
        RECT 989.545 10.965 989.835 12.130 ;
        RECT 1003.805 10.965 1004.095 12.130 ;
        RECT 1018.065 10.965 1018.355 12.130 ;
        RECT 1032.325 10.965 1032.615 12.130 ;
        RECT 1046.585 10.965 1046.875 12.130 ;
        RECT 1060.845 10.965 1061.135 12.130 ;
        RECT 1075.105 10.965 1075.395 12.130 ;
        RECT 1089.365 10.965 1089.655 12.130 ;
        RECT 1103.625 10.965 1103.915 12.130 ;
        RECT 1117.885 10.965 1118.175 12.130 ;
        RECT 1132.145 10.965 1132.435 12.130 ;
        RECT 1146.405 10.965 1146.695 12.130 ;
        RECT 1160.665 10.965 1160.955 12.130 ;
        RECT 1174.925 10.965 1175.215 12.130 ;
        RECT 1189.185 10.965 1189.475 12.130 ;
        RECT 1203.445 10.965 1203.735 12.130 ;
        RECT 1217.705 10.965 1217.995 12.130 ;
        RECT 1231.965 10.965 1232.255 12.130 ;
        RECT 1246.225 10.965 1246.515 12.130 ;
        RECT 1260.485 10.965 1260.775 12.130 ;
        RECT 1274.745 10.965 1275.035 12.130 ;
        RECT 1289.005 10.965 1289.295 12.130 ;
        RECT 1303.265 10.965 1303.555 12.130 ;
        RECT 1317.525 10.965 1317.815 12.130 ;
        RECT 1331.785 10.965 1332.075 12.130 ;
        RECT 1346.045 10.965 1346.335 12.130 ;
        RECT 1360.305 10.965 1360.595 12.130 ;
        RECT 1374.565 10.965 1374.855 12.130 ;
        RECT 1388.825 10.965 1389.115 12.130 ;
        RECT 1403.085 10.965 1403.375 12.130 ;
        RECT 1417.345 10.965 1417.635 12.130 ;
        RECT 1431.605 10.965 1431.895 12.130 ;
        RECT 1445.865 10.965 1446.155 12.130 ;
        RECT 1460.125 10.965 1460.415 12.130 ;
        RECT 1474.385 10.965 1474.675 12.130 ;
        RECT 1488.645 10.965 1488.935 12.130 ;
        RECT 1502.905 10.965 1503.195 12.130 ;
        RECT 1517.165 10.965 1517.455 12.130 ;
        RECT 1531.425 10.965 1531.715 12.130 ;
        RECT 1545.685 10.965 1545.975 12.130 ;
        RECT 1559.945 10.965 1560.235 12.130 ;
        RECT 1574.205 10.965 1574.495 12.130 ;
        RECT 1588.465 10.965 1588.755 12.130 ;
        RECT 1602.725 10.965 1603.015 12.130 ;
        RECT 1616.985 10.965 1617.275 12.130 ;
        RECT 1631.245 10.965 1631.535 12.130 ;
        RECT 1645.505 10.965 1645.795 12.130 ;
        RECT 1659.765 10.965 1660.055 12.130 ;
        RECT 1674.025 10.965 1674.315 12.130 ;
        RECT 1688.285 10.965 1688.575 12.130 ;
        RECT 1702.545 10.965 1702.835 12.130 ;
        RECT 1716.805 10.965 1717.095 12.130 ;
        RECT 1731.065 10.965 1731.355 12.130 ;
        RECT 1745.325 10.965 1745.615 12.130 ;
        RECT 1759.585 10.965 1759.875 12.130 ;
        RECT 1773.845 10.965 1774.135 12.130 ;
        RECT 1788.105 10.965 1788.395 12.130 ;
        RECT 1802.365 10.965 1802.655 12.130 ;
        RECT 1816.625 10.965 1816.915 12.130 ;
        RECT 1830.885 10.965 1831.175 12.130 ;
        RECT 1845.145 10.965 1845.435 12.130 ;
        RECT 1859.405 10.965 1859.695 12.130 ;
        RECT 1873.665 10.965 1873.955 12.130 ;
        RECT 1887.925 10.965 1888.215 12.130 ;
        RECT 1902.185 10.965 1902.475 12.130 ;
        RECT 1916.445 10.965 1916.735 12.130 ;
        RECT 1930.705 10.965 1930.995 12.130 ;
        RECT 1944.965 10.965 1945.255 12.130 ;
        RECT 1959.225 10.965 1959.515 12.130 ;
        RECT 1973.485 10.965 1973.775 12.130 ;
        RECT 1987.745 10.965 1988.035 12.130 ;
        RECT 2002.005 10.965 2002.295 12.130 ;
        RECT 2016.265 10.965 2016.555 12.130 ;
        RECT 2030.525 10.965 2030.815 12.130 ;
        RECT 2044.785 10.965 2045.075 12.130 ;
        RECT 2059.045 10.965 2059.335 12.130 ;
        RECT 2073.305 10.965 2073.595 12.130 ;
        RECT 2087.565 10.965 2087.855 12.130 ;
        RECT 2101.825 10.965 2102.115 12.130 ;
        RECT 2116.085 10.965 2116.375 12.130 ;
        RECT 2130.345 10.965 2130.635 12.130 ;
        RECT 2144.605 10.965 2144.895 12.130 ;
        RECT 2158.865 10.965 2159.155 12.130 ;
        RECT 2173.125 10.965 2173.415 12.130 ;
        RECT 2187.385 10.965 2187.675 12.130 ;
        RECT 2201.645 10.965 2201.935 12.130 ;
        RECT 2215.905 10.965 2216.195 12.130 ;
        RECT 2230.165 10.965 2230.455 12.130 ;
        RECT 2244.425 10.965 2244.715 12.130 ;
        RECT 2258.685 10.965 2258.975 12.130 ;
        RECT 2272.945 10.965 2273.235 12.130 ;
        RECT 2287.205 10.965 2287.495 12.130 ;
        RECT 2301.465 10.965 2301.755 12.130 ;
        RECT 2315.725 10.965 2316.015 12.130 ;
        RECT 2329.985 10.965 2330.275 12.130 ;
        RECT 2344.245 10.965 2344.535 12.130 ;
        RECT 2358.505 10.965 2358.795 12.130 ;
        RECT 2372.765 10.965 2373.055 12.130 ;
        RECT 2387.025 10.965 2387.315 12.130 ;
        RECT 2401.285 10.965 2401.575 12.130 ;
        RECT 2415.545 10.965 2415.835 12.130 ;
        RECT 2429.805 10.965 2430.095 12.130 ;
        RECT 2444.065 10.965 2444.355 12.130 ;
        RECT 2458.325 10.965 2458.615 12.130 ;
        RECT 2472.585 10.965 2472.875 12.130 ;
        RECT 2486.845 10.965 2487.135 12.130 ;
        RECT 2501.105 10.965 2501.395 12.130 ;
        RECT 2515.365 10.965 2515.655 12.130 ;
        RECT 2529.625 10.965 2529.915 12.130 ;
        RECT 2543.885 10.965 2544.175 12.130 ;
        RECT 2558.145 10.965 2558.435 12.130 ;
        RECT 2572.405 10.965 2572.695 12.130 ;
        RECT 2586.665 10.965 2586.955 12.130 ;
        RECT 2600.925 10.965 2601.215 12.130 ;
        RECT 2615.185 10.965 2615.475 12.130 ;
        RECT 2629.445 10.965 2629.735 12.130 ;
        RECT 2643.705 10.965 2643.995 12.130 ;
        RECT 2657.965 10.965 2658.255 12.130 ;
        RECT 2672.225 10.965 2672.515 12.130 ;
        RECT 2686.485 10.965 2686.775 12.130 ;
        RECT 2700.745 10.965 2701.035 12.130 ;
        RECT 2715.005 10.965 2715.295 12.130 ;
        RECT 2729.265 10.965 2729.555 12.130 ;
        RECT 2743.525 10.965 2743.815 12.130 ;
        RECT 2757.785 10.965 2758.075 12.130 ;
        RECT 2772.045 10.965 2772.335 12.130 ;
        RECT 2786.305 10.965 2786.595 12.130 ;
        RECT 2800.565 10.965 2800.855 12.130 ;
        RECT 2814.825 10.965 2815.115 12.130 ;
        RECT 2829.085 10.965 2829.375 12.130 ;
        RECT 2843.345 10.965 2843.635 12.130 ;
        RECT 2857.605 10.965 2857.895 12.130 ;
        RECT 2871.865 10.965 2872.155 12.130 ;
        RECT 2886.125 10.965 2886.415 12.130 ;
        RECT 2900.385 10.965 2900.675 12.130 ;
        RECT 2912.805 12.055 2913.325 12.595 ;
        RECT 2909.315 10.965 2909.645 11.690 ;
        RECT 2912.805 10.965 2914.015 12.055 ;
        RECT 5.520 10.795 6.900 10.965 ;
        RECT 8.740 10.795 11.500 10.965 ;
        RECT 19.780 10.795 20.240 10.965 ;
        RECT 34.040 10.795 34.500 10.965 ;
        RECT 48.300 10.795 48.760 10.965 ;
        RECT 62.560 10.795 63.020 10.965 ;
        RECT 76.820 10.795 77.280 10.965 ;
        RECT 81.880 10.795 90.620 10.965 ;
        RECT 91.080 10.795 91.540 10.965 ;
        RECT 105.340 10.795 105.800 10.965 ;
        RECT 119.600 10.795 120.060 10.965 ;
        RECT 133.860 10.795 134.320 10.965 ;
        RECT 148.120 10.795 148.580 10.965 ;
        RECT 162.380 10.795 162.840 10.965 ;
        RECT 176.640 10.795 177.100 10.965 ;
        RECT 190.900 10.795 191.360 10.965 ;
        RECT 205.160 10.795 212.980 10.965 ;
        RECT 219.420 10.795 219.880 10.965 ;
        RECT 225.400 10.795 231.840 10.965 ;
        RECT 233.680 10.795 234.140 10.965 ;
        RECT 240.120 10.795 244.260 10.965 ;
        RECT 247.940 10.795 248.400 10.965 ;
        RECT 262.200 10.795 269.100 10.965 ;
        RECT 276.460 10.795 276.920 10.965 ;
        RECT 290.720 10.795 291.180 10.965 ;
        RECT 304.980 10.795 305.440 10.965 ;
        RECT 319.240 10.795 319.700 10.965 ;
        RECT 333.500 10.795 333.960 10.965 ;
        RECT 347.760 10.795 348.220 10.965 ;
        RECT 352.360 10.795 353.740 10.965 ;
        RECT 362.020 10.795 362.480 10.965 ;
        RECT 376.280 10.795 376.740 10.965 ;
        RECT 390.540 10.795 401.120 10.965 ;
        RECT 404.800 10.795 405.260 10.965 ;
        RECT 419.060 10.795 419.520 10.965 ;
        RECT 433.320 10.795 433.780 10.965 ;
        RECT 447.580 10.795 448.040 10.965 ;
        RECT 450.800 10.795 457.240 10.965 ;
        RECT 461.840 10.795 462.300 10.965 ;
        RECT 476.100 10.795 476.560 10.965 ;
        RECT 490.360 10.795 490.820 10.965 ;
        RECT 504.620 10.795 505.080 10.965 ;
        RECT 518.880 10.795 519.340 10.965 ;
        RECT 533.140 10.795 533.600 10.965 ;
        RECT 547.400 10.795 547.860 10.965 ;
        RECT 561.660 10.795 562.120 10.965 ;
        RECT 575.920 10.795 576.380 10.965 ;
        RECT 590.180 10.795 590.640 10.965 ;
        RECT 604.440 10.795 604.900 10.965 ;
        RECT 618.700 10.795 619.160 10.965 ;
        RECT 632.960 10.795 633.420 10.965 ;
        RECT 647.220 10.795 647.680 10.965 ;
        RECT 661.480 10.795 661.940 10.965 ;
        RECT 675.740 10.795 676.200 10.965 ;
        RECT 690.000 10.795 690.460 10.965 ;
        RECT 704.260 10.795 704.720 10.965 ;
        RECT 718.520 10.795 718.980 10.965 ;
        RECT 732.780 10.795 733.240 10.965 ;
        RECT 747.040 10.795 747.500 10.965 ;
        RECT 761.300 10.795 761.760 10.965 ;
        RECT 775.560 10.795 776.020 10.965 ;
        RECT 789.820 10.795 790.280 10.965 ;
        RECT 804.080 10.795 804.540 10.965 ;
        RECT 818.340 10.795 818.800 10.965 ;
        RECT 832.600 10.795 833.060 10.965 ;
        RECT 846.860 10.795 847.320 10.965 ;
        RECT 861.120 10.795 861.580 10.965 ;
        RECT 875.380 10.795 875.840 10.965 ;
        RECT 889.640 10.795 890.100 10.965 ;
        RECT 903.900 10.795 904.360 10.965 ;
        RECT 918.160 10.795 918.620 10.965 ;
        RECT 932.420 10.795 932.880 10.965 ;
        RECT 946.680 10.795 947.140 10.965 ;
        RECT 960.940 10.795 961.400 10.965 ;
        RECT 975.200 10.795 975.660 10.965 ;
        RECT 989.460 10.795 989.920 10.965 ;
        RECT 1003.720 10.795 1004.180 10.965 ;
        RECT 1017.980 10.795 1018.440 10.965 ;
        RECT 1032.240 10.795 1032.700 10.965 ;
        RECT 1046.500 10.795 1046.960 10.965 ;
        RECT 1060.760 10.795 1061.220 10.965 ;
        RECT 1075.020 10.795 1075.480 10.965 ;
        RECT 1089.280 10.795 1089.740 10.965 ;
        RECT 1103.540 10.795 1104.000 10.965 ;
        RECT 1117.800 10.795 1118.260 10.965 ;
        RECT 1132.060 10.795 1132.520 10.965 ;
        RECT 1146.320 10.795 1146.780 10.965 ;
        RECT 1160.580 10.795 1161.040 10.965 ;
        RECT 1174.840 10.795 1175.300 10.965 ;
        RECT 1189.100 10.795 1189.560 10.965 ;
        RECT 1203.360 10.795 1203.820 10.965 ;
        RECT 1217.620 10.795 1218.080 10.965 ;
        RECT 1231.880 10.795 1232.340 10.965 ;
        RECT 1246.140 10.795 1246.600 10.965 ;
        RECT 1260.400 10.795 1260.860 10.965 ;
        RECT 1274.660 10.795 1275.120 10.965 ;
        RECT 1288.920 10.795 1289.380 10.965 ;
        RECT 1303.180 10.795 1303.640 10.965 ;
        RECT 1317.440 10.795 1317.900 10.965 ;
        RECT 1331.700 10.795 1332.160 10.965 ;
        RECT 1345.960 10.795 1346.420 10.965 ;
        RECT 1360.220 10.795 1360.680 10.965 ;
        RECT 1374.480 10.795 1374.940 10.965 ;
        RECT 1388.740 10.795 1389.200 10.965 ;
        RECT 1403.000 10.795 1403.460 10.965 ;
        RECT 1417.260 10.795 1417.720 10.965 ;
        RECT 1431.520 10.795 1431.980 10.965 ;
        RECT 1445.780 10.795 1446.240 10.965 ;
        RECT 1460.040 10.795 1460.500 10.965 ;
        RECT 1474.300 10.795 1474.760 10.965 ;
        RECT 1488.560 10.795 1489.020 10.965 ;
        RECT 1502.820 10.795 1503.280 10.965 ;
        RECT 1517.080 10.795 1517.540 10.965 ;
        RECT 1531.340 10.795 1531.800 10.965 ;
        RECT 1545.600 10.795 1546.060 10.965 ;
        RECT 1559.860 10.795 1560.320 10.965 ;
        RECT 1574.120 10.795 1574.580 10.965 ;
        RECT 1588.380 10.795 1588.840 10.965 ;
        RECT 1602.640 10.795 1603.100 10.965 ;
        RECT 1616.900 10.795 1617.360 10.965 ;
        RECT 1631.160 10.795 1631.620 10.965 ;
        RECT 1645.420 10.795 1645.880 10.965 ;
        RECT 1659.680 10.795 1660.140 10.965 ;
        RECT 1673.940 10.795 1674.400 10.965 ;
        RECT 1688.200 10.795 1688.660 10.965 ;
        RECT 1702.460 10.795 1702.920 10.965 ;
        RECT 1716.720 10.795 1717.180 10.965 ;
        RECT 1730.980 10.795 1731.440 10.965 ;
        RECT 1745.240 10.795 1745.700 10.965 ;
        RECT 1759.500 10.795 1759.960 10.965 ;
        RECT 1773.760 10.795 1774.220 10.965 ;
        RECT 1788.020 10.795 1788.480 10.965 ;
        RECT 1802.280 10.795 1802.740 10.965 ;
        RECT 1816.540 10.795 1817.000 10.965 ;
        RECT 1830.800 10.795 1831.260 10.965 ;
        RECT 1845.060 10.795 1845.520 10.965 ;
        RECT 1859.320 10.795 1859.780 10.965 ;
        RECT 1873.580 10.795 1874.040 10.965 ;
        RECT 1887.840 10.795 1888.300 10.965 ;
        RECT 1902.100 10.795 1902.560 10.965 ;
        RECT 1916.360 10.795 1916.820 10.965 ;
        RECT 1930.620 10.795 1931.080 10.965 ;
        RECT 1944.880 10.795 1945.340 10.965 ;
        RECT 1959.140 10.795 1959.600 10.965 ;
        RECT 1973.400 10.795 1973.860 10.965 ;
        RECT 1987.660 10.795 1988.120 10.965 ;
        RECT 2001.920 10.795 2002.380 10.965 ;
        RECT 2016.180 10.795 2016.640 10.965 ;
        RECT 2030.440 10.795 2030.900 10.965 ;
        RECT 2044.700 10.795 2045.160 10.965 ;
        RECT 2058.960 10.795 2059.420 10.965 ;
        RECT 2073.220 10.795 2073.680 10.965 ;
        RECT 2087.480 10.795 2087.940 10.965 ;
        RECT 2101.740 10.795 2102.200 10.965 ;
        RECT 2116.000 10.795 2116.460 10.965 ;
        RECT 2130.260 10.795 2130.720 10.965 ;
        RECT 2144.520 10.795 2144.980 10.965 ;
        RECT 2158.780 10.795 2159.240 10.965 ;
        RECT 2173.040 10.795 2173.500 10.965 ;
        RECT 2187.300 10.795 2187.760 10.965 ;
        RECT 2201.560 10.795 2202.020 10.965 ;
        RECT 2215.820 10.795 2216.280 10.965 ;
        RECT 2230.080 10.795 2230.540 10.965 ;
        RECT 2244.340 10.795 2244.800 10.965 ;
        RECT 2258.600 10.795 2259.060 10.965 ;
        RECT 2272.860 10.795 2273.320 10.965 ;
        RECT 2287.120 10.795 2287.580 10.965 ;
        RECT 2301.380 10.795 2301.840 10.965 ;
        RECT 2315.640 10.795 2316.100 10.965 ;
        RECT 2329.900 10.795 2330.360 10.965 ;
        RECT 2344.160 10.795 2344.620 10.965 ;
        RECT 2358.420 10.795 2358.880 10.965 ;
        RECT 2372.680 10.795 2373.140 10.965 ;
        RECT 2386.940 10.795 2387.400 10.965 ;
        RECT 2401.200 10.795 2401.660 10.965 ;
        RECT 2415.460 10.795 2415.920 10.965 ;
        RECT 2429.720 10.795 2430.180 10.965 ;
        RECT 2443.980 10.795 2444.440 10.965 ;
        RECT 2458.240 10.795 2458.700 10.965 ;
        RECT 2472.500 10.795 2472.960 10.965 ;
        RECT 2486.760 10.795 2487.220 10.965 ;
        RECT 2501.020 10.795 2501.480 10.965 ;
        RECT 2515.280 10.795 2515.740 10.965 ;
        RECT 2529.540 10.795 2530.000 10.965 ;
        RECT 2543.800 10.795 2544.260 10.965 ;
        RECT 2558.060 10.795 2558.520 10.965 ;
        RECT 2572.320 10.795 2572.780 10.965 ;
        RECT 2586.580 10.795 2587.040 10.965 ;
        RECT 2600.840 10.795 2601.300 10.965 ;
        RECT 2615.100 10.795 2615.560 10.965 ;
        RECT 2629.360 10.795 2629.820 10.965 ;
        RECT 2643.620 10.795 2644.080 10.965 ;
        RECT 2657.880 10.795 2658.340 10.965 ;
        RECT 2672.140 10.795 2672.600 10.965 ;
        RECT 2686.400 10.795 2686.860 10.965 ;
        RECT 2700.660 10.795 2701.120 10.965 ;
        RECT 2714.920 10.795 2715.380 10.965 ;
        RECT 2729.180 10.795 2729.640 10.965 ;
        RECT 2743.440 10.795 2743.900 10.965 ;
        RECT 2757.700 10.795 2758.160 10.965 ;
        RECT 2771.960 10.795 2772.420 10.965 ;
        RECT 2786.220 10.795 2786.680 10.965 ;
        RECT 2800.480 10.795 2800.940 10.965 ;
        RECT 2814.740 10.795 2815.200 10.965 ;
        RECT 2829.000 10.795 2829.460 10.965 ;
        RECT 2843.260 10.795 2843.720 10.965 ;
        RECT 2857.520 10.795 2857.980 10.965 ;
        RECT 2871.780 10.795 2872.240 10.965 ;
        RECT 2886.040 10.795 2886.500 10.965 ;
        RECT 2900.300 10.795 2900.760 10.965 ;
        RECT 2909.040 10.795 2910.420 10.965 ;
        RECT 2912.720 10.795 2914.100 10.965 ;
      LAYER mcon ;
        RECT 5.665 3508.715 5.835 3508.885 ;
        RECT 6.125 3508.715 6.295 3508.885 ;
        RECT 6.585 3508.715 6.755 3508.885 ;
        RECT 19.925 3508.715 20.095 3508.885 ;
        RECT 34.185 3508.715 34.355 3508.885 ;
        RECT 48.445 3508.715 48.615 3508.885 ;
        RECT 62.705 3508.715 62.875 3508.885 ;
        RECT 76.965 3508.715 77.135 3508.885 ;
        RECT 91.225 3508.715 91.395 3508.885 ;
        RECT 105.485 3508.715 105.655 3508.885 ;
        RECT 119.745 3508.715 119.915 3508.885 ;
        RECT 134.005 3508.715 134.175 3508.885 ;
        RECT 148.265 3508.715 148.435 3508.885 ;
        RECT 162.525 3508.715 162.695 3508.885 ;
        RECT 176.785 3508.715 176.955 3508.885 ;
        RECT 191.045 3508.715 191.215 3508.885 ;
        RECT 205.305 3508.715 205.475 3508.885 ;
        RECT 219.565 3508.715 219.735 3508.885 ;
        RECT 233.825 3508.715 233.995 3508.885 ;
        RECT 248.085 3508.715 248.255 3508.885 ;
        RECT 262.345 3508.715 262.515 3508.885 ;
        RECT 276.605 3508.715 276.775 3508.885 ;
        RECT 290.865 3508.715 291.035 3508.885 ;
        RECT 305.125 3508.715 305.295 3508.885 ;
        RECT 319.385 3508.715 319.555 3508.885 ;
        RECT 333.645 3508.715 333.815 3508.885 ;
        RECT 347.905 3508.715 348.075 3508.885 ;
        RECT 362.165 3508.715 362.335 3508.885 ;
        RECT 376.425 3508.715 376.595 3508.885 ;
        RECT 390.685 3508.715 390.855 3508.885 ;
        RECT 404.945 3508.715 405.115 3508.885 ;
        RECT 419.205 3508.715 419.375 3508.885 ;
        RECT 433.465 3508.715 433.635 3508.885 ;
        RECT 447.725 3508.715 447.895 3508.885 ;
        RECT 461.985 3508.715 462.155 3508.885 ;
        RECT 476.245 3508.715 476.415 3508.885 ;
        RECT 490.505 3508.715 490.675 3508.885 ;
        RECT 504.765 3508.715 504.935 3508.885 ;
        RECT 519.025 3508.715 519.195 3508.885 ;
        RECT 533.285 3508.715 533.455 3508.885 ;
        RECT 547.545 3508.715 547.715 3508.885 ;
        RECT 561.805 3508.715 561.975 3508.885 ;
        RECT 576.065 3508.715 576.235 3508.885 ;
        RECT 590.325 3508.715 590.495 3508.885 ;
        RECT 604.585 3508.715 604.755 3508.885 ;
        RECT 618.845 3508.715 619.015 3508.885 ;
        RECT 633.105 3508.715 633.275 3508.885 ;
        RECT 647.365 3508.715 647.535 3508.885 ;
        RECT 661.625 3508.715 661.795 3508.885 ;
        RECT 675.885 3508.715 676.055 3508.885 ;
        RECT 690.145 3508.715 690.315 3508.885 ;
        RECT 704.405 3508.715 704.575 3508.885 ;
        RECT 718.665 3508.715 718.835 3508.885 ;
        RECT 732.925 3508.715 733.095 3508.885 ;
        RECT 747.185 3508.715 747.355 3508.885 ;
        RECT 761.445 3508.715 761.615 3508.885 ;
        RECT 775.705 3508.715 775.875 3508.885 ;
        RECT 789.965 3508.715 790.135 3508.885 ;
        RECT 804.225 3508.715 804.395 3508.885 ;
        RECT 818.485 3508.715 818.655 3508.885 ;
        RECT 832.745 3508.715 832.915 3508.885 ;
        RECT 847.005 3508.715 847.175 3508.885 ;
        RECT 861.265 3508.715 861.435 3508.885 ;
        RECT 875.525 3508.715 875.695 3508.885 ;
        RECT 889.785 3508.715 889.955 3508.885 ;
        RECT 904.045 3508.715 904.215 3508.885 ;
        RECT 918.305 3508.715 918.475 3508.885 ;
        RECT 932.565 3508.715 932.735 3508.885 ;
        RECT 946.825 3508.715 946.995 3508.885 ;
        RECT 961.085 3508.715 961.255 3508.885 ;
        RECT 975.345 3508.715 975.515 3508.885 ;
        RECT 989.605 3508.715 989.775 3508.885 ;
        RECT 1003.865 3508.715 1004.035 3508.885 ;
        RECT 1018.125 3508.715 1018.295 3508.885 ;
        RECT 1032.385 3508.715 1032.555 3508.885 ;
        RECT 1046.645 3508.715 1046.815 3508.885 ;
        RECT 1060.905 3508.715 1061.075 3508.885 ;
        RECT 1075.165 3508.715 1075.335 3508.885 ;
        RECT 1089.425 3508.715 1089.595 3508.885 ;
        RECT 1103.685 3508.715 1103.855 3508.885 ;
        RECT 1117.945 3508.715 1118.115 3508.885 ;
        RECT 1132.205 3508.715 1132.375 3508.885 ;
        RECT 1146.465 3508.715 1146.635 3508.885 ;
        RECT 1160.725 3508.715 1160.895 3508.885 ;
        RECT 1174.985 3508.715 1175.155 3508.885 ;
        RECT 1189.245 3508.715 1189.415 3508.885 ;
        RECT 1203.505 3508.715 1203.675 3508.885 ;
        RECT 1217.765 3508.715 1217.935 3508.885 ;
        RECT 1232.025 3508.715 1232.195 3508.885 ;
        RECT 1246.285 3508.715 1246.455 3508.885 ;
        RECT 1260.545 3508.715 1260.715 3508.885 ;
        RECT 1274.805 3508.715 1274.975 3508.885 ;
        RECT 1289.065 3508.715 1289.235 3508.885 ;
        RECT 1303.325 3508.715 1303.495 3508.885 ;
        RECT 1317.585 3508.715 1317.755 3508.885 ;
        RECT 1331.845 3508.715 1332.015 3508.885 ;
        RECT 1346.105 3508.715 1346.275 3508.885 ;
        RECT 1360.365 3508.715 1360.535 3508.885 ;
        RECT 1374.625 3508.715 1374.795 3508.885 ;
        RECT 1388.885 3508.715 1389.055 3508.885 ;
        RECT 1403.145 3508.715 1403.315 3508.885 ;
        RECT 1417.405 3508.715 1417.575 3508.885 ;
        RECT 1431.665 3508.715 1431.835 3508.885 ;
        RECT 1445.925 3508.715 1446.095 3508.885 ;
        RECT 1460.185 3508.715 1460.355 3508.885 ;
        RECT 1474.445 3508.715 1474.615 3508.885 ;
        RECT 1488.705 3508.715 1488.875 3508.885 ;
        RECT 1502.965 3508.715 1503.135 3508.885 ;
        RECT 1517.225 3508.715 1517.395 3508.885 ;
        RECT 1531.485 3508.715 1531.655 3508.885 ;
        RECT 1545.745 3508.715 1545.915 3508.885 ;
        RECT 1560.005 3508.715 1560.175 3508.885 ;
        RECT 1574.265 3508.715 1574.435 3508.885 ;
        RECT 1588.525 3508.715 1588.695 3508.885 ;
        RECT 1602.785 3508.715 1602.955 3508.885 ;
        RECT 1617.045 3508.715 1617.215 3508.885 ;
        RECT 1631.305 3508.715 1631.475 3508.885 ;
        RECT 1645.565 3508.715 1645.735 3508.885 ;
        RECT 1659.825 3508.715 1659.995 3508.885 ;
        RECT 1674.085 3508.715 1674.255 3508.885 ;
        RECT 1688.345 3508.715 1688.515 3508.885 ;
        RECT 1702.605 3508.715 1702.775 3508.885 ;
        RECT 1716.865 3508.715 1717.035 3508.885 ;
        RECT 1731.125 3508.715 1731.295 3508.885 ;
        RECT 1745.385 3508.715 1745.555 3508.885 ;
        RECT 1759.645 3508.715 1759.815 3508.885 ;
        RECT 1773.905 3508.715 1774.075 3508.885 ;
        RECT 1788.165 3508.715 1788.335 3508.885 ;
        RECT 1802.425 3508.715 1802.595 3508.885 ;
        RECT 1816.685 3508.715 1816.855 3508.885 ;
        RECT 1830.945 3508.715 1831.115 3508.885 ;
        RECT 1845.205 3508.715 1845.375 3508.885 ;
        RECT 1859.465 3508.715 1859.635 3508.885 ;
        RECT 1873.725 3508.715 1873.895 3508.885 ;
        RECT 1887.985 3508.715 1888.155 3508.885 ;
        RECT 1902.245 3508.715 1902.415 3508.885 ;
        RECT 1916.505 3508.715 1916.675 3508.885 ;
        RECT 1930.765 3508.715 1930.935 3508.885 ;
        RECT 1945.025 3508.715 1945.195 3508.885 ;
        RECT 1959.285 3508.715 1959.455 3508.885 ;
        RECT 1973.545 3508.715 1973.715 3508.885 ;
        RECT 1987.805 3508.715 1987.975 3508.885 ;
        RECT 2002.065 3508.715 2002.235 3508.885 ;
        RECT 2016.325 3508.715 2016.495 3508.885 ;
        RECT 2030.585 3508.715 2030.755 3508.885 ;
        RECT 2044.845 3508.715 2045.015 3508.885 ;
        RECT 2059.105 3508.715 2059.275 3508.885 ;
        RECT 2073.365 3508.715 2073.535 3508.885 ;
        RECT 2087.625 3508.715 2087.795 3508.885 ;
        RECT 2101.885 3508.715 2102.055 3508.885 ;
        RECT 2116.145 3508.715 2116.315 3508.885 ;
        RECT 2130.405 3508.715 2130.575 3508.885 ;
        RECT 2144.665 3508.715 2144.835 3508.885 ;
        RECT 2158.925 3508.715 2159.095 3508.885 ;
        RECT 2173.185 3508.715 2173.355 3508.885 ;
        RECT 2187.445 3508.715 2187.615 3508.885 ;
        RECT 2201.705 3508.715 2201.875 3508.885 ;
        RECT 2215.965 3508.715 2216.135 3508.885 ;
        RECT 2230.225 3508.715 2230.395 3508.885 ;
        RECT 2244.485 3508.715 2244.655 3508.885 ;
        RECT 2258.745 3508.715 2258.915 3508.885 ;
        RECT 2273.005 3508.715 2273.175 3508.885 ;
        RECT 2287.265 3508.715 2287.435 3508.885 ;
        RECT 2301.525 3508.715 2301.695 3508.885 ;
        RECT 2315.785 3508.715 2315.955 3508.885 ;
        RECT 2330.045 3508.715 2330.215 3508.885 ;
        RECT 2344.305 3508.715 2344.475 3508.885 ;
        RECT 2358.565 3508.715 2358.735 3508.885 ;
        RECT 2372.825 3508.715 2372.995 3508.885 ;
        RECT 2387.085 3508.715 2387.255 3508.885 ;
        RECT 2401.345 3508.715 2401.515 3508.885 ;
        RECT 2415.605 3508.715 2415.775 3508.885 ;
        RECT 2429.865 3508.715 2430.035 3508.885 ;
        RECT 2444.125 3508.715 2444.295 3508.885 ;
        RECT 2458.385 3508.715 2458.555 3508.885 ;
        RECT 2472.645 3508.715 2472.815 3508.885 ;
        RECT 2486.905 3508.715 2487.075 3508.885 ;
        RECT 2501.165 3508.715 2501.335 3508.885 ;
        RECT 2515.425 3508.715 2515.595 3508.885 ;
        RECT 2529.685 3508.715 2529.855 3508.885 ;
        RECT 2543.945 3508.715 2544.115 3508.885 ;
        RECT 2558.205 3508.715 2558.375 3508.885 ;
        RECT 2572.465 3508.715 2572.635 3508.885 ;
        RECT 2586.725 3508.715 2586.895 3508.885 ;
        RECT 2600.985 3508.715 2601.155 3508.885 ;
        RECT 2615.245 3508.715 2615.415 3508.885 ;
        RECT 2629.505 3508.715 2629.675 3508.885 ;
        RECT 2643.765 3508.715 2643.935 3508.885 ;
        RECT 2658.025 3508.715 2658.195 3508.885 ;
        RECT 2672.285 3508.715 2672.455 3508.885 ;
        RECT 2686.545 3508.715 2686.715 3508.885 ;
        RECT 2700.805 3508.715 2700.975 3508.885 ;
        RECT 2715.065 3508.715 2715.235 3508.885 ;
        RECT 2729.325 3508.715 2729.495 3508.885 ;
        RECT 2743.585 3508.715 2743.755 3508.885 ;
        RECT 2757.845 3508.715 2758.015 3508.885 ;
        RECT 2772.105 3508.715 2772.275 3508.885 ;
        RECT 2786.365 3508.715 2786.535 3508.885 ;
        RECT 2800.625 3508.715 2800.795 3508.885 ;
        RECT 2814.885 3508.715 2815.055 3508.885 ;
        RECT 2829.145 3508.715 2829.315 3508.885 ;
        RECT 2843.405 3508.715 2843.575 3508.885 ;
        RECT 2857.665 3508.715 2857.835 3508.885 ;
        RECT 2871.925 3508.715 2872.095 3508.885 ;
        RECT 2886.185 3508.715 2886.355 3508.885 ;
        RECT 2900.445 3508.715 2900.615 3508.885 ;
        RECT 2912.865 3508.715 2913.035 3508.885 ;
        RECT 2913.325 3508.715 2913.495 3508.885 ;
        RECT 2913.785 3508.715 2913.955 3508.885 ;
        RECT 5.665 3503.275 5.835 3503.445 ;
        RECT 6.125 3503.275 6.295 3503.445 ;
        RECT 6.585 3503.275 6.755 3503.445 ;
        RECT 9.805 3503.275 9.975 3503.445 ;
        RECT 10.265 3503.275 10.435 3503.445 ;
        RECT 10.725 3503.275 10.895 3503.445 ;
        RECT 11.185 3503.275 11.355 3503.445 ;
        RECT 11.645 3503.275 11.815 3503.445 ;
        RECT 12.105 3503.275 12.275 3503.445 ;
        RECT 2909.185 3503.275 2909.355 3503.445 ;
        RECT 2909.645 3503.275 2909.815 3503.445 ;
        RECT 2910.105 3503.275 2910.275 3503.445 ;
        RECT 2910.565 3503.275 2910.735 3503.445 ;
        RECT 2911.025 3503.275 2911.195 3503.445 ;
        RECT 2911.485 3503.275 2911.655 3503.445 ;
        RECT 2912.865 3503.275 2913.035 3503.445 ;
        RECT 2913.325 3503.275 2913.495 3503.445 ;
        RECT 2913.785 3503.275 2913.955 3503.445 ;
        RECT 5.665 3497.835 5.835 3498.005 ;
        RECT 6.125 3497.835 6.295 3498.005 ;
        RECT 6.585 3497.835 6.755 3498.005 ;
        RECT 2910.105 3497.835 2910.275 3498.005 ;
        RECT 2912.865 3497.835 2913.035 3498.005 ;
        RECT 2913.325 3497.835 2913.495 3498.005 ;
        RECT 2913.785 3497.835 2913.955 3498.005 ;
        RECT 5.665 3492.395 5.835 3492.565 ;
        RECT 6.125 3492.395 6.295 3492.565 ;
        RECT 6.585 3492.395 6.755 3492.565 ;
        RECT 2910.105 3492.395 2910.275 3492.565 ;
        RECT 2912.865 3492.395 2913.035 3492.565 ;
        RECT 2913.325 3492.395 2913.495 3492.565 ;
        RECT 2913.785 3492.395 2913.955 3492.565 ;
        RECT 5.665 3486.955 5.835 3487.125 ;
        RECT 6.125 3486.955 6.295 3487.125 ;
        RECT 6.585 3486.955 6.755 3487.125 ;
        RECT 2910.105 3486.955 2910.275 3487.125 ;
        RECT 2912.865 3486.955 2913.035 3487.125 ;
        RECT 2913.325 3486.955 2913.495 3487.125 ;
        RECT 2913.785 3486.955 2913.955 3487.125 ;
        RECT 5.665 3481.515 5.835 3481.685 ;
        RECT 6.125 3481.515 6.295 3481.685 ;
        RECT 6.585 3481.515 6.755 3481.685 ;
        RECT 2910.105 3481.515 2910.275 3481.685 ;
        RECT 2912.865 3481.515 2913.035 3481.685 ;
        RECT 2913.325 3481.515 2913.495 3481.685 ;
        RECT 2913.785 3481.515 2913.955 3481.685 ;
        RECT 5.665 3476.075 5.835 3476.245 ;
        RECT 6.125 3476.075 6.295 3476.245 ;
        RECT 6.585 3476.075 6.755 3476.245 ;
        RECT 2910.105 3476.075 2910.275 3476.245 ;
        RECT 2912.865 3476.075 2913.035 3476.245 ;
        RECT 2913.325 3476.075 2913.495 3476.245 ;
        RECT 2913.785 3476.075 2913.955 3476.245 ;
        RECT 5.665 3470.635 5.835 3470.805 ;
        RECT 6.125 3470.635 6.295 3470.805 ;
        RECT 6.585 3470.635 6.755 3470.805 ;
        RECT 2910.105 3470.635 2910.275 3470.805 ;
        RECT 2912.865 3470.635 2913.035 3470.805 ;
        RECT 2913.325 3470.635 2913.495 3470.805 ;
        RECT 2913.785 3470.635 2913.955 3470.805 ;
        RECT 5.665 3465.195 5.835 3465.365 ;
        RECT 6.125 3465.195 6.295 3465.365 ;
        RECT 6.585 3465.195 6.755 3465.365 ;
        RECT 2910.105 3465.195 2910.275 3465.365 ;
        RECT 2912.865 3465.195 2913.035 3465.365 ;
        RECT 2913.325 3465.195 2913.495 3465.365 ;
        RECT 2913.785 3465.195 2913.955 3465.365 ;
        RECT 5.665 3459.755 5.835 3459.925 ;
        RECT 6.125 3459.755 6.295 3459.925 ;
        RECT 6.585 3459.755 6.755 3459.925 ;
        RECT 2910.105 3459.755 2910.275 3459.925 ;
        RECT 2912.865 3459.755 2913.035 3459.925 ;
        RECT 2913.325 3459.755 2913.495 3459.925 ;
        RECT 2913.785 3459.755 2913.955 3459.925 ;
        RECT 5.665 3454.315 5.835 3454.485 ;
        RECT 6.125 3454.315 6.295 3454.485 ;
        RECT 6.585 3454.315 6.755 3454.485 ;
        RECT 2910.105 3454.315 2910.275 3454.485 ;
        RECT 2912.865 3454.315 2913.035 3454.485 ;
        RECT 2913.325 3454.315 2913.495 3454.485 ;
        RECT 2913.785 3454.315 2913.955 3454.485 ;
        RECT 5.665 3448.875 5.835 3449.045 ;
        RECT 6.125 3448.875 6.295 3449.045 ;
        RECT 6.585 3448.875 6.755 3449.045 ;
        RECT 2910.105 3448.875 2910.275 3449.045 ;
        RECT 2912.865 3448.875 2913.035 3449.045 ;
        RECT 2913.325 3448.875 2913.495 3449.045 ;
        RECT 2913.785 3448.875 2913.955 3449.045 ;
        RECT 5.665 3443.435 5.835 3443.605 ;
        RECT 6.125 3443.435 6.295 3443.605 ;
        RECT 6.585 3443.435 6.755 3443.605 ;
        RECT 2910.105 3443.435 2910.275 3443.605 ;
        RECT 2912.865 3443.435 2913.035 3443.605 ;
        RECT 2913.325 3443.435 2913.495 3443.605 ;
        RECT 2913.785 3443.435 2913.955 3443.605 ;
        RECT 5.665 3437.995 5.835 3438.165 ;
        RECT 6.125 3437.995 6.295 3438.165 ;
        RECT 6.585 3437.995 6.755 3438.165 ;
        RECT 2910.105 3437.995 2910.275 3438.165 ;
        RECT 2912.865 3437.995 2913.035 3438.165 ;
        RECT 2913.325 3437.995 2913.495 3438.165 ;
        RECT 2913.785 3437.995 2913.955 3438.165 ;
        RECT 5.665 3432.555 5.835 3432.725 ;
        RECT 6.125 3432.555 6.295 3432.725 ;
        RECT 6.585 3432.555 6.755 3432.725 ;
        RECT 2910.105 3432.555 2910.275 3432.725 ;
        RECT 2912.865 3432.555 2913.035 3432.725 ;
        RECT 2913.325 3432.555 2913.495 3432.725 ;
        RECT 2913.785 3432.555 2913.955 3432.725 ;
        RECT 5.665 3427.115 5.835 3427.285 ;
        RECT 6.125 3427.115 6.295 3427.285 ;
        RECT 6.585 3427.115 6.755 3427.285 ;
        RECT 2910.105 3427.115 2910.275 3427.285 ;
        RECT 2912.865 3427.115 2913.035 3427.285 ;
        RECT 2913.325 3427.115 2913.495 3427.285 ;
        RECT 2913.785 3427.115 2913.955 3427.285 ;
        RECT 5.665 3421.675 5.835 3421.845 ;
        RECT 6.125 3421.675 6.295 3421.845 ;
        RECT 6.585 3421.675 6.755 3421.845 ;
        RECT 2910.105 3421.675 2910.275 3421.845 ;
        RECT 2912.865 3421.675 2913.035 3421.845 ;
        RECT 2913.325 3421.675 2913.495 3421.845 ;
        RECT 2913.785 3421.675 2913.955 3421.845 ;
        RECT 5.665 3416.235 5.835 3416.405 ;
        RECT 6.125 3416.235 6.295 3416.405 ;
        RECT 6.585 3416.235 6.755 3416.405 ;
        RECT 2910.105 3416.235 2910.275 3416.405 ;
        RECT 2912.865 3416.235 2913.035 3416.405 ;
        RECT 2913.325 3416.235 2913.495 3416.405 ;
        RECT 2913.785 3416.235 2913.955 3416.405 ;
        RECT 5.665 3410.795 5.835 3410.965 ;
        RECT 6.125 3410.795 6.295 3410.965 ;
        RECT 6.585 3410.795 6.755 3410.965 ;
        RECT 2910.105 3410.795 2910.275 3410.965 ;
        RECT 2912.865 3410.795 2913.035 3410.965 ;
        RECT 2913.325 3410.795 2913.495 3410.965 ;
        RECT 2913.785 3410.795 2913.955 3410.965 ;
        RECT 5.665 3405.355 5.835 3405.525 ;
        RECT 6.125 3405.355 6.295 3405.525 ;
        RECT 6.585 3405.355 6.755 3405.525 ;
        RECT 2910.105 3405.355 2910.275 3405.525 ;
        RECT 2912.865 3405.355 2913.035 3405.525 ;
        RECT 2913.325 3405.355 2913.495 3405.525 ;
        RECT 2913.785 3405.355 2913.955 3405.525 ;
        RECT 5.665 3399.915 5.835 3400.085 ;
        RECT 6.125 3399.915 6.295 3400.085 ;
        RECT 6.585 3399.915 6.755 3400.085 ;
        RECT 2909.185 3399.915 2909.355 3400.085 ;
        RECT 2909.645 3399.915 2909.815 3400.085 ;
        RECT 2910.105 3399.915 2910.275 3400.085 ;
        RECT 2912.865 3399.915 2913.035 3400.085 ;
        RECT 2913.325 3399.915 2913.495 3400.085 ;
        RECT 2913.785 3399.915 2913.955 3400.085 ;
        RECT 5.665 3394.475 5.835 3394.645 ;
        RECT 6.125 3394.475 6.295 3394.645 ;
        RECT 6.585 3394.475 6.755 3394.645 ;
        RECT 2910.105 3394.475 2910.275 3394.645 ;
        RECT 2912.865 3394.475 2913.035 3394.645 ;
        RECT 2913.325 3394.475 2913.495 3394.645 ;
        RECT 2913.785 3394.475 2913.955 3394.645 ;
        RECT 5.665 3389.035 5.835 3389.205 ;
        RECT 6.125 3389.035 6.295 3389.205 ;
        RECT 6.585 3389.035 6.755 3389.205 ;
        RECT 2910.105 3389.035 2910.275 3389.205 ;
        RECT 2912.865 3389.035 2913.035 3389.205 ;
        RECT 2913.325 3389.035 2913.495 3389.205 ;
        RECT 2913.785 3389.035 2913.955 3389.205 ;
        RECT 5.665 3383.595 5.835 3383.765 ;
        RECT 6.125 3383.595 6.295 3383.765 ;
        RECT 6.585 3383.595 6.755 3383.765 ;
        RECT 2910.105 3383.595 2910.275 3383.765 ;
        RECT 2912.865 3383.595 2913.035 3383.765 ;
        RECT 2913.325 3383.595 2913.495 3383.765 ;
        RECT 2913.785 3383.595 2913.955 3383.765 ;
        RECT 5.665 3378.155 5.835 3378.325 ;
        RECT 6.125 3378.155 6.295 3378.325 ;
        RECT 6.585 3378.155 6.755 3378.325 ;
        RECT 2910.105 3378.155 2910.275 3378.325 ;
        RECT 2912.865 3378.155 2913.035 3378.325 ;
        RECT 2913.325 3378.155 2913.495 3378.325 ;
        RECT 2913.785 3378.155 2913.955 3378.325 ;
        RECT 5.665 3372.715 5.835 3372.885 ;
        RECT 6.125 3372.715 6.295 3372.885 ;
        RECT 6.585 3372.715 6.755 3372.885 ;
        RECT 2910.105 3372.715 2910.275 3372.885 ;
        RECT 2912.865 3372.715 2913.035 3372.885 ;
        RECT 2913.325 3372.715 2913.495 3372.885 ;
        RECT 2913.785 3372.715 2913.955 3372.885 ;
        RECT 5.665 3367.275 5.835 3367.445 ;
        RECT 6.125 3367.275 6.295 3367.445 ;
        RECT 6.585 3367.275 6.755 3367.445 ;
        RECT 2910.105 3367.275 2910.275 3367.445 ;
        RECT 2910.565 3367.275 2910.735 3367.445 ;
        RECT 2911.025 3367.275 2911.195 3367.445 ;
        RECT 2911.485 3367.275 2911.655 3367.445 ;
        RECT 2912.865 3367.275 2913.035 3367.445 ;
        RECT 2913.325 3367.275 2913.495 3367.445 ;
        RECT 2913.785 3367.275 2913.955 3367.445 ;
        RECT 5.665 3361.835 5.835 3362.005 ;
        RECT 6.125 3361.835 6.295 3362.005 ;
        RECT 6.585 3361.835 6.755 3362.005 ;
        RECT 2910.105 3361.835 2910.275 3362.005 ;
        RECT 2912.865 3361.835 2913.035 3362.005 ;
        RECT 2913.325 3361.835 2913.495 3362.005 ;
        RECT 2913.785 3361.835 2913.955 3362.005 ;
        RECT 5.665 3356.395 5.835 3356.565 ;
        RECT 6.125 3356.395 6.295 3356.565 ;
        RECT 6.585 3356.395 6.755 3356.565 ;
        RECT 2910.105 3356.395 2910.275 3356.565 ;
        RECT 2912.865 3356.395 2913.035 3356.565 ;
        RECT 2913.325 3356.395 2913.495 3356.565 ;
        RECT 2913.785 3356.395 2913.955 3356.565 ;
        RECT 5.665 3350.955 5.835 3351.125 ;
        RECT 6.125 3350.955 6.295 3351.125 ;
        RECT 6.585 3350.955 6.755 3351.125 ;
        RECT 2910.105 3350.955 2910.275 3351.125 ;
        RECT 2912.865 3350.955 2913.035 3351.125 ;
        RECT 2913.325 3350.955 2913.495 3351.125 ;
        RECT 2913.785 3350.955 2913.955 3351.125 ;
        RECT 5.665 3345.515 5.835 3345.685 ;
        RECT 6.125 3345.515 6.295 3345.685 ;
        RECT 6.585 3345.515 6.755 3345.685 ;
        RECT 2910.105 3345.515 2910.275 3345.685 ;
        RECT 2912.865 3345.515 2913.035 3345.685 ;
        RECT 2913.325 3345.515 2913.495 3345.685 ;
        RECT 2913.785 3345.515 2913.955 3345.685 ;
        RECT 5.665 3340.075 5.835 3340.245 ;
        RECT 6.125 3340.075 6.295 3340.245 ;
        RECT 6.585 3340.075 6.755 3340.245 ;
        RECT 2910.105 3340.075 2910.275 3340.245 ;
        RECT 2912.865 3340.075 2913.035 3340.245 ;
        RECT 2913.325 3340.075 2913.495 3340.245 ;
        RECT 2913.785 3340.075 2913.955 3340.245 ;
        RECT 5.665 3334.635 5.835 3334.805 ;
        RECT 6.125 3334.635 6.295 3334.805 ;
        RECT 6.585 3334.635 6.755 3334.805 ;
        RECT 2910.105 3334.635 2910.275 3334.805 ;
        RECT 2912.865 3334.635 2913.035 3334.805 ;
        RECT 2913.325 3334.635 2913.495 3334.805 ;
        RECT 2913.785 3334.635 2913.955 3334.805 ;
        RECT 5.665 3329.195 5.835 3329.365 ;
        RECT 6.125 3329.195 6.295 3329.365 ;
        RECT 6.585 3329.195 6.755 3329.365 ;
        RECT 2910.105 3329.195 2910.275 3329.365 ;
        RECT 2912.865 3329.195 2913.035 3329.365 ;
        RECT 2913.325 3329.195 2913.495 3329.365 ;
        RECT 2913.785 3329.195 2913.955 3329.365 ;
        RECT 5.665 3323.755 5.835 3323.925 ;
        RECT 6.125 3323.755 6.295 3323.925 ;
        RECT 6.585 3323.755 6.755 3323.925 ;
        RECT 2910.105 3323.755 2910.275 3323.925 ;
        RECT 2912.865 3323.755 2913.035 3323.925 ;
        RECT 2913.325 3323.755 2913.495 3323.925 ;
        RECT 2913.785 3323.755 2913.955 3323.925 ;
        RECT 5.665 3318.315 5.835 3318.485 ;
        RECT 6.125 3318.315 6.295 3318.485 ;
        RECT 6.585 3318.315 6.755 3318.485 ;
        RECT 2910.105 3318.315 2910.275 3318.485 ;
        RECT 2912.865 3318.315 2913.035 3318.485 ;
        RECT 2913.325 3318.315 2913.495 3318.485 ;
        RECT 2913.785 3318.315 2913.955 3318.485 ;
        RECT 5.665 3312.875 5.835 3313.045 ;
        RECT 6.125 3312.875 6.295 3313.045 ;
        RECT 6.585 3312.875 6.755 3313.045 ;
        RECT 2910.105 3312.875 2910.275 3313.045 ;
        RECT 2912.865 3312.875 2913.035 3313.045 ;
        RECT 2913.325 3312.875 2913.495 3313.045 ;
        RECT 2913.785 3312.875 2913.955 3313.045 ;
        RECT 5.665 3307.435 5.835 3307.605 ;
        RECT 6.125 3307.435 6.295 3307.605 ;
        RECT 6.585 3307.435 6.755 3307.605 ;
        RECT 2910.105 3307.435 2910.275 3307.605 ;
        RECT 2912.865 3307.435 2913.035 3307.605 ;
        RECT 2913.325 3307.435 2913.495 3307.605 ;
        RECT 2913.785 3307.435 2913.955 3307.605 ;
        RECT 5.665 3301.995 5.835 3302.165 ;
        RECT 6.125 3301.995 6.295 3302.165 ;
        RECT 6.585 3301.995 6.755 3302.165 ;
        RECT 2910.105 3301.995 2910.275 3302.165 ;
        RECT 2912.865 3301.995 2913.035 3302.165 ;
        RECT 2913.325 3301.995 2913.495 3302.165 ;
        RECT 2913.785 3301.995 2913.955 3302.165 ;
        RECT 5.665 3296.555 5.835 3296.725 ;
        RECT 6.125 3296.555 6.295 3296.725 ;
        RECT 6.585 3296.555 6.755 3296.725 ;
        RECT 2910.105 3296.555 2910.275 3296.725 ;
        RECT 2912.865 3296.555 2913.035 3296.725 ;
        RECT 2913.325 3296.555 2913.495 3296.725 ;
        RECT 2913.785 3296.555 2913.955 3296.725 ;
        RECT 5.665 3291.115 5.835 3291.285 ;
        RECT 6.125 3291.115 6.295 3291.285 ;
        RECT 6.585 3291.115 6.755 3291.285 ;
        RECT 2910.105 3291.115 2910.275 3291.285 ;
        RECT 2912.865 3291.115 2913.035 3291.285 ;
        RECT 2913.325 3291.115 2913.495 3291.285 ;
        RECT 2913.785 3291.115 2913.955 3291.285 ;
        RECT 5.665 3285.675 5.835 3285.845 ;
        RECT 6.125 3285.675 6.295 3285.845 ;
        RECT 6.585 3285.675 6.755 3285.845 ;
        RECT 2910.105 3285.675 2910.275 3285.845 ;
        RECT 2912.865 3285.675 2913.035 3285.845 ;
        RECT 2913.325 3285.675 2913.495 3285.845 ;
        RECT 2913.785 3285.675 2913.955 3285.845 ;
        RECT 5.665 3280.235 5.835 3280.405 ;
        RECT 6.125 3280.235 6.295 3280.405 ;
        RECT 6.585 3280.235 6.755 3280.405 ;
        RECT 2910.105 3280.235 2910.275 3280.405 ;
        RECT 2912.865 3280.235 2913.035 3280.405 ;
        RECT 2913.325 3280.235 2913.495 3280.405 ;
        RECT 2913.785 3280.235 2913.955 3280.405 ;
        RECT 5.665 3274.795 5.835 3274.965 ;
        RECT 6.125 3274.795 6.295 3274.965 ;
        RECT 6.585 3274.795 6.755 3274.965 ;
        RECT 2910.105 3274.795 2910.275 3274.965 ;
        RECT 2912.865 3274.795 2913.035 3274.965 ;
        RECT 2913.325 3274.795 2913.495 3274.965 ;
        RECT 2913.785 3274.795 2913.955 3274.965 ;
        RECT 5.665 3269.355 5.835 3269.525 ;
        RECT 6.125 3269.355 6.295 3269.525 ;
        RECT 6.585 3269.355 6.755 3269.525 ;
        RECT 2910.105 3269.355 2910.275 3269.525 ;
        RECT 2912.865 3269.355 2913.035 3269.525 ;
        RECT 2913.325 3269.355 2913.495 3269.525 ;
        RECT 2913.785 3269.355 2913.955 3269.525 ;
        RECT 5.665 3263.915 5.835 3264.085 ;
        RECT 6.125 3263.915 6.295 3264.085 ;
        RECT 6.585 3263.915 6.755 3264.085 ;
        RECT 2910.105 3263.915 2910.275 3264.085 ;
        RECT 2912.865 3263.915 2913.035 3264.085 ;
        RECT 2913.325 3263.915 2913.495 3264.085 ;
        RECT 2913.785 3263.915 2913.955 3264.085 ;
        RECT 5.665 3258.475 5.835 3258.645 ;
        RECT 6.125 3258.475 6.295 3258.645 ;
        RECT 6.585 3258.475 6.755 3258.645 ;
        RECT 2910.105 3258.475 2910.275 3258.645 ;
        RECT 2912.865 3258.475 2913.035 3258.645 ;
        RECT 2913.325 3258.475 2913.495 3258.645 ;
        RECT 2913.785 3258.475 2913.955 3258.645 ;
        RECT 5.665 3253.035 5.835 3253.205 ;
        RECT 6.125 3253.035 6.295 3253.205 ;
        RECT 6.585 3253.035 6.755 3253.205 ;
        RECT 2910.105 3253.035 2910.275 3253.205 ;
        RECT 2912.865 3253.035 2913.035 3253.205 ;
        RECT 2913.325 3253.035 2913.495 3253.205 ;
        RECT 2913.785 3253.035 2913.955 3253.205 ;
        RECT 5.665 3247.595 5.835 3247.765 ;
        RECT 6.125 3247.595 6.295 3247.765 ;
        RECT 6.585 3247.595 6.755 3247.765 ;
        RECT 2910.105 3247.595 2910.275 3247.765 ;
        RECT 2912.865 3247.595 2913.035 3247.765 ;
        RECT 2913.325 3247.595 2913.495 3247.765 ;
        RECT 2913.785 3247.595 2913.955 3247.765 ;
        RECT 5.665 3242.155 5.835 3242.325 ;
        RECT 6.125 3242.155 6.295 3242.325 ;
        RECT 6.585 3242.155 6.755 3242.325 ;
        RECT 2910.105 3242.155 2910.275 3242.325 ;
        RECT 2912.865 3242.155 2913.035 3242.325 ;
        RECT 2913.325 3242.155 2913.495 3242.325 ;
        RECT 2913.785 3242.155 2913.955 3242.325 ;
        RECT 5.665 3236.715 5.835 3236.885 ;
        RECT 6.125 3236.715 6.295 3236.885 ;
        RECT 6.585 3236.715 6.755 3236.885 ;
        RECT 2910.105 3236.715 2910.275 3236.885 ;
        RECT 2912.865 3236.715 2913.035 3236.885 ;
        RECT 2913.325 3236.715 2913.495 3236.885 ;
        RECT 2913.785 3236.715 2913.955 3236.885 ;
        RECT 5.665 3231.275 5.835 3231.445 ;
        RECT 6.125 3231.275 6.295 3231.445 ;
        RECT 6.585 3231.275 6.755 3231.445 ;
        RECT 2910.105 3231.275 2910.275 3231.445 ;
        RECT 2912.865 3231.275 2913.035 3231.445 ;
        RECT 2913.325 3231.275 2913.495 3231.445 ;
        RECT 2913.785 3231.275 2913.955 3231.445 ;
        RECT 5.665 3225.835 5.835 3226.005 ;
        RECT 6.125 3225.835 6.295 3226.005 ;
        RECT 6.585 3225.835 6.755 3226.005 ;
        RECT 8.885 3225.835 9.055 3226.005 ;
        RECT 9.345 3225.835 9.515 3226.005 ;
        RECT 9.805 3225.835 9.975 3226.005 ;
        RECT 2910.105 3225.835 2910.275 3226.005 ;
        RECT 2912.865 3225.835 2913.035 3226.005 ;
        RECT 2913.325 3225.835 2913.495 3226.005 ;
        RECT 2913.785 3225.835 2913.955 3226.005 ;
        RECT 5.665 3220.395 5.835 3220.565 ;
        RECT 6.125 3220.395 6.295 3220.565 ;
        RECT 6.585 3220.395 6.755 3220.565 ;
        RECT 2910.105 3220.395 2910.275 3220.565 ;
        RECT 2912.865 3220.395 2913.035 3220.565 ;
        RECT 2913.325 3220.395 2913.495 3220.565 ;
        RECT 2913.785 3220.395 2913.955 3220.565 ;
        RECT 5.665 3214.955 5.835 3215.125 ;
        RECT 6.125 3214.955 6.295 3215.125 ;
        RECT 6.585 3214.955 6.755 3215.125 ;
        RECT 2910.105 3214.955 2910.275 3215.125 ;
        RECT 2912.865 3214.955 2913.035 3215.125 ;
        RECT 2913.325 3214.955 2913.495 3215.125 ;
        RECT 2913.785 3214.955 2913.955 3215.125 ;
        RECT 5.665 3209.515 5.835 3209.685 ;
        RECT 6.125 3209.515 6.295 3209.685 ;
        RECT 6.585 3209.515 6.755 3209.685 ;
        RECT 2910.105 3209.515 2910.275 3209.685 ;
        RECT 2912.865 3209.515 2913.035 3209.685 ;
        RECT 2913.325 3209.515 2913.495 3209.685 ;
        RECT 2913.785 3209.515 2913.955 3209.685 ;
        RECT 5.665 3204.075 5.835 3204.245 ;
        RECT 6.125 3204.075 6.295 3204.245 ;
        RECT 6.585 3204.075 6.755 3204.245 ;
        RECT 2910.105 3204.075 2910.275 3204.245 ;
        RECT 2910.565 3204.075 2910.735 3204.245 ;
        RECT 2911.025 3204.075 2911.195 3204.245 ;
        RECT 2911.485 3204.075 2911.655 3204.245 ;
        RECT 2912.865 3204.075 2913.035 3204.245 ;
        RECT 2913.325 3204.075 2913.495 3204.245 ;
        RECT 2913.785 3204.075 2913.955 3204.245 ;
        RECT 5.665 3198.635 5.835 3198.805 ;
        RECT 6.125 3198.635 6.295 3198.805 ;
        RECT 6.585 3198.635 6.755 3198.805 ;
        RECT 2910.105 3198.635 2910.275 3198.805 ;
        RECT 2912.865 3198.635 2913.035 3198.805 ;
        RECT 2913.325 3198.635 2913.495 3198.805 ;
        RECT 2913.785 3198.635 2913.955 3198.805 ;
        RECT 5.665 3193.195 5.835 3193.365 ;
        RECT 6.125 3193.195 6.295 3193.365 ;
        RECT 6.585 3193.195 6.755 3193.365 ;
        RECT 2910.105 3193.195 2910.275 3193.365 ;
        RECT 2912.865 3193.195 2913.035 3193.365 ;
        RECT 2913.325 3193.195 2913.495 3193.365 ;
        RECT 2913.785 3193.195 2913.955 3193.365 ;
        RECT 5.665 3187.755 5.835 3187.925 ;
        RECT 6.125 3187.755 6.295 3187.925 ;
        RECT 6.585 3187.755 6.755 3187.925 ;
        RECT 2910.105 3187.755 2910.275 3187.925 ;
        RECT 2912.865 3187.755 2913.035 3187.925 ;
        RECT 2913.325 3187.755 2913.495 3187.925 ;
        RECT 2913.785 3187.755 2913.955 3187.925 ;
        RECT 5.665 3182.315 5.835 3182.485 ;
        RECT 6.125 3182.315 6.295 3182.485 ;
        RECT 6.585 3182.315 6.755 3182.485 ;
        RECT 2910.105 3182.315 2910.275 3182.485 ;
        RECT 2912.865 3182.315 2913.035 3182.485 ;
        RECT 2913.325 3182.315 2913.495 3182.485 ;
        RECT 2913.785 3182.315 2913.955 3182.485 ;
        RECT 5.665 3176.875 5.835 3177.045 ;
        RECT 6.125 3176.875 6.295 3177.045 ;
        RECT 6.585 3176.875 6.755 3177.045 ;
        RECT 2910.105 3176.875 2910.275 3177.045 ;
        RECT 2912.865 3176.875 2913.035 3177.045 ;
        RECT 2913.325 3176.875 2913.495 3177.045 ;
        RECT 2913.785 3176.875 2913.955 3177.045 ;
        RECT 5.665 3171.435 5.835 3171.605 ;
        RECT 6.125 3171.435 6.295 3171.605 ;
        RECT 6.585 3171.435 6.755 3171.605 ;
        RECT 2910.105 3171.435 2910.275 3171.605 ;
        RECT 2912.865 3171.435 2913.035 3171.605 ;
        RECT 2913.325 3171.435 2913.495 3171.605 ;
        RECT 2913.785 3171.435 2913.955 3171.605 ;
        RECT 5.665 3165.995 5.835 3166.165 ;
        RECT 6.125 3165.995 6.295 3166.165 ;
        RECT 6.585 3165.995 6.755 3166.165 ;
        RECT 2910.105 3165.995 2910.275 3166.165 ;
        RECT 2912.865 3165.995 2913.035 3166.165 ;
        RECT 2913.325 3165.995 2913.495 3166.165 ;
        RECT 2913.785 3165.995 2913.955 3166.165 ;
        RECT 5.665 3160.555 5.835 3160.725 ;
        RECT 6.125 3160.555 6.295 3160.725 ;
        RECT 6.585 3160.555 6.755 3160.725 ;
        RECT 2910.105 3160.555 2910.275 3160.725 ;
        RECT 2912.865 3160.555 2913.035 3160.725 ;
        RECT 2913.325 3160.555 2913.495 3160.725 ;
        RECT 2913.785 3160.555 2913.955 3160.725 ;
        RECT 5.665 3155.115 5.835 3155.285 ;
        RECT 6.125 3155.115 6.295 3155.285 ;
        RECT 6.585 3155.115 6.755 3155.285 ;
        RECT 2910.105 3155.115 2910.275 3155.285 ;
        RECT 2912.865 3155.115 2913.035 3155.285 ;
        RECT 2913.325 3155.115 2913.495 3155.285 ;
        RECT 2913.785 3155.115 2913.955 3155.285 ;
        RECT 5.665 3149.675 5.835 3149.845 ;
        RECT 6.125 3149.675 6.295 3149.845 ;
        RECT 6.585 3149.675 6.755 3149.845 ;
        RECT 2910.105 3149.675 2910.275 3149.845 ;
        RECT 2912.865 3149.675 2913.035 3149.845 ;
        RECT 2913.325 3149.675 2913.495 3149.845 ;
        RECT 2913.785 3149.675 2913.955 3149.845 ;
        RECT 5.665 3144.235 5.835 3144.405 ;
        RECT 6.125 3144.235 6.295 3144.405 ;
        RECT 6.585 3144.235 6.755 3144.405 ;
        RECT 2910.105 3144.235 2910.275 3144.405 ;
        RECT 2912.865 3144.235 2913.035 3144.405 ;
        RECT 2913.325 3144.235 2913.495 3144.405 ;
        RECT 2913.785 3144.235 2913.955 3144.405 ;
        RECT 5.665 3138.795 5.835 3138.965 ;
        RECT 6.125 3138.795 6.295 3138.965 ;
        RECT 6.585 3138.795 6.755 3138.965 ;
        RECT 2910.105 3138.795 2910.275 3138.965 ;
        RECT 2912.865 3138.795 2913.035 3138.965 ;
        RECT 2913.325 3138.795 2913.495 3138.965 ;
        RECT 2913.785 3138.795 2913.955 3138.965 ;
        RECT 5.665 3133.355 5.835 3133.525 ;
        RECT 6.125 3133.355 6.295 3133.525 ;
        RECT 6.585 3133.355 6.755 3133.525 ;
        RECT 2910.105 3133.355 2910.275 3133.525 ;
        RECT 2912.865 3133.355 2913.035 3133.525 ;
        RECT 2913.325 3133.355 2913.495 3133.525 ;
        RECT 2913.785 3133.355 2913.955 3133.525 ;
        RECT 5.665 3127.915 5.835 3128.085 ;
        RECT 6.125 3127.915 6.295 3128.085 ;
        RECT 6.585 3127.915 6.755 3128.085 ;
        RECT 2910.105 3127.915 2910.275 3128.085 ;
        RECT 2912.865 3127.915 2913.035 3128.085 ;
        RECT 2913.325 3127.915 2913.495 3128.085 ;
        RECT 2913.785 3127.915 2913.955 3128.085 ;
        RECT 5.665 3122.475 5.835 3122.645 ;
        RECT 6.125 3122.475 6.295 3122.645 ;
        RECT 6.585 3122.475 6.755 3122.645 ;
        RECT 2910.105 3122.475 2910.275 3122.645 ;
        RECT 2912.865 3122.475 2913.035 3122.645 ;
        RECT 2913.325 3122.475 2913.495 3122.645 ;
        RECT 2913.785 3122.475 2913.955 3122.645 ;
        RECT 5.665 3117.035 5.835 3117.205 ;
        RECT 6.125 3117.035 6.295 3117.205 ;
        RECT 6.585 3117.035 6.755 3117.205 ;
        RECT 2910.105 3117.035 2910.275 3117.205 ;
        RECT 2912.865 3117.035 2913.035 3117.205 ;
        RECT 2913.325 3117.035 2913.495 3117.205 ;
        RECT 2913.785 3117.035 2913.955 3117.205 ;
        RECT 5.665 3111.595 5.835 3111.765 ;
        RECT 6.125 3111.595 6.295 3111.765 ;
        RECT 6.585 3111.595 6.755 3111.765 ;
        RECT 2910.105 3111.595 2910.275 3111.765 ;
        RECT 2912.865 3111.595 2913.035 3111.765 ;
        RECT 2913.325 3111.595 2913.495 3111.765 ;
        RECT 2913.785 3111.595 2913.955 3111.765 ;
        RECT 5.665 3106.155 5.835 3106.325 ;
        RECT 6.125 3106.155 6.295 3106.325 ;
        RECT 6.585 3106.155 6.755 3106.325 ;
        RECT 2910.105 3106.155 2910.275 3106.325 ;
        RECT 2912.865 3106.155 2913.035 3106.325 ;
        RECT 2913.325 3106.155 2913.495 3106.325 ;
        RECT 2913.785 3106.155 2913.955 3106.325 ;
        RECT 5.665 3100.715 5.835 3100.885 ;
        RECT 6.125 3100.715 6.295 3100.885 ;
        RECT 6.585 3100.715 6.755 3100.885 ;
        RECT 2910.105 3100.715 2910.275 3100.885 ;
        RECT 2912.865 3100.715 2913.035 3100.885 ;
        RECT 2913.325 3100.715 2913.495 3100.885 ;
        RECT 2913.785 3100.715 2913.955 3100.885 ;
        RECT 5.665 3095.275 5.835 3095.445 ;
        RECT 6.125 3095.275 6.295 3095.445 ;
        RECT 6.585 3095.275 6.755 3095.445 ;
        RECT 2909.185 3095.275 2909.355 3095.445 ;
        RECT 2909.645 3095.275 2909.815 3095.445 ;
        RECT 2910.105 3095.275 2910.275 3095.445 ;
        RECT 2912.865 3095.275 2913.035 3095.445 ;
        RECT 2913.325 3095.275 2913.495 3095.445 ;
        RECT 2913.785 3095.275 2913.955 3095.445 ;
        RECT 5.665 3089.835 5.835 3090.005 ;
        RECT 6.125 3089.835 6.295 3090.005 ;
        RECT 6.585 3089.835 6.755 3090.005 ;
        RECT 2910.105 3089.835 2910.275 3090.005 ;
        RECT 2912.865 3089.835 2913.035 3090.005 ;
        RECT 2913.325 3089.835 2913.495 3090.005 ;
        RECT 2913.785 3089.835 2913.955 3090.005 ;
        RECT 5.665 3084.395 5.835 3084.565 ;
        RECT 6.125 3084.395 6.295 3084.565 ;
        RECT 6.585 3084.395 6.755 3084.565 ;
        RECT 2910.105 3084.395 2910.275 3084.565 ;
        RECT 2912.865 3084.395 2913.035 3084.565 ;
        RECT 2913.325 3084.395 2913.495 3084.565 ;
        RECT 2913.785 3084.395 2913.955 3084.565 ;
        RECT 5.665 3078.955 5.835 3079.125 ;
        RECT 6.125 3078.955 6.295 3079.125 ;
        RECT 6.585 3078.955 6.755 3079.125 ;
        RECT 2910.105 3078.955 2910.275 3079.125 ;
        RECT 2912.865 3078.955 2913.035 3079.125 ;
        RECT 2913.325 3078.955 2913.495 3079.125 ;
        RECT 2913.785 3078.955 2913.955 3079.125 ;
        RECT 5.665 3073.515 5.835 3073.685 ;
        RECT 6.125 3073.515 6.295 3073.685 ;
        RECT 6.585 3073.515 6.755 3073.685 ;
        RECT 2910.105 3073.515 2910.275 3073.685 ;
        RECT 2912.865 3073.515 2913.035 3073.685 ;
        RECT 2913.325 3073.515 2913.495 3073.685 ;
        RECT 2913.785 3073.515 2913.955 3073.685 ;
        RECT 5.665 3068.075 5.835 3068.245 ;
        RECT 6.125 3068.075 6.295 3068.245 ;
        RECT 6.585 3068.075 6.755 3068.245 ;
        RECT 2910.105 3068.075 2910.275 3068.245 ;
        RECT 2912.865 3068.075 2913.035 3068.245 ;
        RECT 2913.325 3068.075 2913.495 3068.245 ;
        RECT 2913.785 3068.075 2913.955 3068.245 ;
        RECT 5.665 3062.635 5.835 3062.805 ;
        RECT 6.125 3062.635 6.295 3062.805 ;
        RECT 6.585 3062.635 6.755 3062.805 ;
        RECT 2910.105 3062.635 2910.275 3062.805 ;
        RECT 2912.865 3062.635 2913.035 3062.805 ;
        RECT 2913.325 3062.635 2913.495 3062.805 ;
        RECT 2913.785 3062.635 2913.955 3062.805 ;
        RECT 5.665 3057.195 5.835 3057.365 ;
        RECT 6.125 3057.195 6.295 3057.365 ;
        RECT 6.585 3057.195 6.755 3057.365 ;
        RECT 2910.105 3057.195 2910.275 3057.365 ;
        RECT 2912.865 3057.195 2913.035 3057.365 ;
        RECT 2913.325 3057.195 2913.495 3057.365 ;
        RECT 2913.785 3057.195 2913.955 3057.365 ;
        RECT 5.665 3051.755 5.835 3051.925 ;
        RECT 6.125 3051.755 6.295 3051.925 ;
        RECT 6.585 3051.755 6.755 3051.925 ;
        RECT 2910.105 3051.755 2910.275 3051.925 ;
        RECT 2912.865 3051.755 2913.035 3051.925 ;
        RECT 2913.325 3051.755 2913.495 3051.925 ;
        RECT 2913.785 3051.755 2913.955 3051.925 ;
        RECT 5.665 3046.315 5.835 3046.485 ;
        RECT 6.125 3046.315 6.295 3046.485 ;
        RECT 6.585 3046.315 6.755 3046.485 ;
        RECT 2910.105 3046.315 2910.275 3046.485 ;
        RECT 2912.865 3046.315 2913.035 3046.485 ;
        RECT 2913.325 3046.315 2913.495 3046.485 ;
        RECT 2913.785 3046.315 2913.955 3046.485 ;
        RECT 5.665 3040.875 5.835 3041.045 ;
        RECT 6.125 3040.875 6.295 3041.045 ;
        RECT 6.585 3040.875 6.755 3041.045 ;
        RECT 2910.105 3040.875 2910.275 3041.045 ;
        RECT 2912.865 3040.875 2913.035 3041.045 ;
        RECT 2913.325 3040.875 2913.495 3041.045 ;
        RECT 2913.785 3040.875 2913.955 3041.045 ;
        RECT 5.665 3035.435 5.835 3035.605 ;
        RECT 6.125 3035.435 6.295 3035.605 ;
        RECT 6.585 3035.435 6.755 3035.605 ;
        RECT 2910.105 3035.435 2910.275 3035.605 ;
        RECT 2912.865 3035.435 2913.035 3035.605 ;
        RECT 2913.325 3035.435 2913.495 3035.605 ;
        RECT 2913.785 3035.435 2913.955 3035.605 ;
        RECT 5.665 3029.995 5.835 3030.165 ;
        RECT 6.125 3029.995 6.295 3030.165 ;
        RECT 6.585 3029.995 6.755 3030.165 ;
        RECT 2910.105 3029.995 2910.275 3030.165 ;
        RECT 2912.865 3029.995 2913.035 3030.165 ;
        RECT 2913.325 3029.995 2913.495 3030.165 ;
        RECT 2913.785 3029.995 2913.955 3030.165 ;
        RECT 5.665 3024.555 5.835 3024.725 ;
        RECT 6.125 3024.555 6.295 3024.725 ;
        RECT 6.585 3024.555 6.755 3024.725 ;
        RECT 2910.105 3024.555 2910.275 3024.725 ;
        RECT 2912.865 3024.555 2913.035 3024.725 ;
        RECT 2913.325 3024.555 2913.495 3024.725 ;
        RECT 2913.785 3024.555 2913.955 3024.725 ;
        RECT 5.665 3019.115 5.835 3019.285 ;
        RECT 6.125 3019.115 6.295 3019.285 ;
        RECT 6.585 3019.115 6.755 3019.285 ;
        RECT 2910.105 3019.115 2910.275 3019.285 ;
        RECT 2912.865 3019.115 2913.035 3019.285 ;
        RECT 2913.325 3019.115 2913.495 3019.285 ;
        RECT 2913.785 3019.115 2913.955 3019.285 ;
        RECT 5.665 3013.675 5.835 3013.845 ;
        RECT 6.125 3013.675 6.295 3013.845 ;
        RECT 6.585 3013.675 6.755 3013.845 ;
        RECT 8.885 3013.675 9.055 3013.845 ;
        RECT 9.345 3013.675 9.515 3013.845 ;
        RECT 9.805 3013.675 9.975 3013.845 ;
        RECT 2910.105 3013.675 2910.275 3013.845 ;
        RECT 2912.865 3013.675 2913.035 3013.845 ;
        RECT 2913.325 3013.675 2913.495 3013.845 ;
        RECT 2913.785 3013.675 2913.955 3013.845 ;
        RECT 5.665 3008.235 5.835 3008.405 ;
        RECT 6.125 3008.235 6.295 3008.405 ;
        RECT 6.585 3008.235 6.755 3008.405 ;
        RECT 2910.105 3008.235 2910.275 3008.405 ;
        RECT 2912.865 3008.235 2913.035 3008.405 ;
        RECT 2913.325 3008.235 2913.495 3008.405 ;
        RECT 2913.785 3008.235 2913.955 3008.405 ;
        RECT 5.665 3002.795 5.835 3002.965 ;
        RECT 6.125 3002.795 6.295 3002.965 ;
        RECT 6.585 3002.795 6.755 3002.965 ;
        RECT 2910.105 3002.795 2910.275 3002.965 ;
        RECT 2912.865 3002.795 2913.035 3002.965 ;
        RECT 2913.325 3002.795 2913.495 3002.965 ;
        RECT 2913.785 3002.795 2913.955 3002.965 ;
        RECT 5.665 2997.355 5.835 2997.525 ;
        RECT 6.125 2997.355 6.295 2997.525 ;
        RECT 6.585 2997.355 6.755 2997.525 ;
        RECT 2910.105 2997.355 2910.275 2997.525 ;
        RECT 2912.865 2997.355 2913.035 2997.525 ;
        RECT 2913.325 2997.355 2913.495 2997.525 ;
        RECT 2913.785 2997.355 2913.955 2997.525 ;
        RECT 5.665 2991.915 5.835 2992.085 ;
        RECT 6.125 2991.915 6.295 2992.085 ;
        RECT 6.585 2991.915 6.755 2992.085 ;
        RECT 2910.105 2991.915 2910.275 2992.085 ;
        RECT 2912.865 2991.915 2913.035 2992.085 ;
        RECT 2913.325 2991.915 2913.495 2992.085 ;
        RECT 2913.785 2991.915 2913.955 2992.085 ;
        RECT 5.665 2986.475 5.835 2986.645 ;
        RECT 6.125 2986.475 6.295 2986.645 ;
        RECT 6.585 2986.475 6.755 2986.645 ;
        RECT 2910.105 2986.475 2910.275 2986.645 ;
        RECT 2912.865 2986.475 2913.035 2986.645 ;
        RECT 2913.325 2986.475 2913.495 2986.645 ;
        RECT 2913.785 2986.475 2913.955 2986.645 ;
        RECT 5.665 2981.035 5.835 2981.205 ;
        RECT 6.125 2981.035 6.295 2981.205 ;
        RECT 6.585 2981.035 6.755 2981.205 ;
        RECT 2910.105 2981.035 2910.275 2981.205 ;
        RECT 2912.865 2981.035 2913.035 2981.205 ;
        RECT 2913.325 2981.035 2913.495 2981.205 ;
        RECT 2913.785 2981.035 2913.955 2981.205 ;
        RECT 5.665 2975.595 5.835 2975.765 ;
        RECT 6.125 2975.595 6.295 2975.765 ;
        RECT 6.585 2975.595 6.755 2975.765 ;
        RECT 2910.105 2975.595 2910.275 2975.765 ;
        RECT 2912.865 2975.595 2913.035 2975.765 ;
        RECT 2913.325 2975.595 2913.495 2975.765 ;
        RECT 2913.785 2975.595 2913.955 2975.765 ;
        RECT 5.665 2970.155 5.835 2970.325 ;
        RECT 6.125 2970.155 6.295 2970.325 ;
        RECT 6.585 2970.155 6.755 2970.325 ;
        RECT 8.885 2970.155 9.055 2970.325 ;
        RECT 9.345 2970.155 9.515 2970.325 ;
        RECT 9.805 2970.155 9.975 2970.325 ;
        RECT 2910.105 2970.155 2910.275 2970.325 ;
        RECT 2912.865 2970.155 2913.035 2970.325 ;
        RECT 2913.325 2970.155 2913.495 2970.325 ;
        RECT 2913.785 2970.155 2913.955 2970.325 ;
        RECT 5.665 2964.715 5.835 2964.885 ;
        RECT 6.125 2964.715 6.295 2964.885 ;
        RECT 6.585 2964.715 6.755 2964.885 ;
        RECT 2910.105 2964.715 2910.275 2964.885 ;
        RECT 2912.865 2964.715 2913.035 2964.885 ;
        RECT 2913.325 2964.715 2913.495 2964.885 ;
        RECT 2913.785 2964.715 2913.955 2964.885 ;
        RECT 5.665 2959.275 5.835 2959.445 ;
        RECT 6.125 2959.275 6.295 2959.445 ;
        RECT 6.585 2959.275 6.755 2959.445 ;
        RECT 2910.105 2959.275 2910.275 2959.445 ;
        RECT 2912.865 2959.275 2913.035 2959.445 ;
        RECT 2913.325 2959.275 2913.495 2959.445 ;
        RECT 2913.785 2959.275 2913.955 2959.445 ;
        RECT 5.665 2953.835 5.835 2954.005 ;
        RECT 6.125 2953.835 6.295 2954.005 ;
        RECT 6.585 2953.835 6.755 2954.005 ;
        RECT 8.885 2953.835 9.055 2954.005 ;
        RECT 9.345 2953.835 9.515 2954.005 ;
        RECT 9.805 2953.835 9.975 2954.005 ;
        RECT 2910.105 2953.835 2910.275 2954.005 ;
        RECT 2912.865 2953.835 2913.035 2954.005 ;
        RECT 2913.325 2953.835 2913.495 2954.005 ;
        RECT 2913.785 2953.835 2913.955 2954.005 ;
        RECT 5.665 2948.395 5.835 2948.565 ;
        RECT 6.125 2948.395 6.295 2948.565 ;
        RECT 6.585 2948.395 6.755 2948.565 ;
        RECT 2910.105 2948.395 2910.275 2948.565 ;
        RECT 2912.865 2948.395 2913.035 2948.565 ;
        RECT 2913.325 2948.395 2913.495 2948.565 ;
        RECT 2913.785 2948.395 2913.955 2948.565 ;
        RECT 5.665 2942.955 5.835 2943.125 ;
        RECT 6.125 2942.955 6.295 2943.125 ;
        RECT 6.585 2942.955 6.755 2943.125 ;
        RECT 2910.105 2942.955 2910.275 2943.125 ;
        RECT 2912.865 2942.955 2913.035 2943.125 ;
        RECT 2913.325 2942.955 2913.495 2943.125 ;
        RECT 2913.785 2942.955 2913.955 2943.125 ;
        RECT 5.665 2937.515 5.835 2937.685 ;
        RECT 6.125 2937.515 6.295 2937.685 ;
        RECT 6.585 2937.515 6.755 2937.685 ;
        RECT 2910.105 2937.515 2910.275 2937.685 ;
        RECT 2912.865 2937.515 2913.035 2937.685 ;
        RECT 2913.325 2937.515 2913.495 2937.685 ;
        RECT 2913.785 2937.515 2913.955 2937.685 ;
        RECT 5.665 2932.075 5.835 2932.245 ;
        RECT 6.125 2932.075 6.295 2932.245 ;
        RECT 6.585 2932.075 6.755 2932.245 ;
        RECT 2910.105 2932.075 2910.275 2932.245 ;
        RECT 2912.865 2932.075 2913.035 2932.245 ;
        RECT 2913.325 2932.075 2913.495 2932.245 ;
        RECT 2913.785 2932.075 2913.955 2932.245 ;
        RECT 5.665 2926.635 5.835 2926.805 ;
        RECT 6.125 2926.635 6.295 2926.805 ;
        RECT 6.585 2926.635 6.755 2926.805 ;
        RECT 2910.105 2926.635 2910.275 2926.805 ;
        RECT 2912.865 2926.635 2913.035 2926.805 ;
        RECT 2913.325 2926.635 2913.495 2926.805 ;
        RECT 2913.785 2926.635 2913.955 2926.805 ;
        RECT 5.665 2921.195 5.835 2921.365 ;
        RECT 6.125 2921.195 6.295 2921.365 ;
        RECT 6.585 2921.195 6.755 2921.365 ;
        RECT 2910.105 2921.195 2910.275 2921.365 ;
        RECT 2912.865 2921.195 2913.035 2921.365 ;
        RECT 2913.325 2921.195 2913.495 2921.365 ;
        RECT 2913.785 2921.195 2913.955 2921.365 ;
        RECT 5.665 2915.755 5.835 2915.925 ;
        RECT 6.125 2915.755 6.295 2915.925 ;
        RECT 6.585 2915.755 6.755 2915.925 ;
        RECT 2910.105 2915.755 2910.275 2915.925 ;
        RECT 2910.565 2915.755 2910.735 2915.925 ;
        RECT 2911.025 2915.755 2911.195 2915.925 ;
        RECT 2911.485 2915.755 2911.655 2915.925 ;
        RECT 2912.865 2915.755 2913.035 2915.925 ;
        RECT 2913.325 2915.755 2913.495 2915.925 ;
        RECT 2913.785 2915.755 2913.955 2915.925 ;
        RECT 5.665 2910.315 5.835 2910.485 ;
        RECT 6.125 2910.315 6.295 2910.485 ;
        RECT 6.585 2910.315 6.755 2910.485 ;
        RECT 2910.105 2910.315 2910.275 2910.485 ;
        RECT 2912.865 2910.315 2913.035 2910.485 ;
        RECT 2913.325 2910.315 2913.495 2910.485 ;
        RECT 2913.785 2910.315 2913.955 2910.485 ;
        RECT 5.665 2904.875 5.835 2905.045 ;
        RECT 6.125 2904.875 6.295 2905.045 ;
        RECT 6.585 2904.875 6.755 2905.045 ;
        RECT 2910.105 2904.875 2910.275 2905.045 ;
        RECT 2912.865 2904.875 2913.035 2905.045 ;
        RECT 2913.325 2904.875 2913.495 2905.045 ;
        RECT 2913.785 2904.875 2913.955 2905.045 ;
        RECT 5.665 2899.435 5.835 2899.605 ;
        RECT 6.125 2899.435 6.295 2899.605 ;
        RECT 6.585 2899.435 6.755 2899.605 ;
        RECT 2910.105 2899.435 2910.275 2899.605 ;
        RECT 2912.865 2899.435 2913.035 2899.605 ;
        RECT 2913.325 2899.435 2913.495 2899.605 ;
        RECT 2913.785 2899.435 2913.955 2899.605 ;
        RECT 5.665 2893.995 5.835 2894.165 ;
        RECT 6.125 2893.995 6.295 2894.165 ;
        RECT 6.585 2893.995 6.755 2894.165 ;
        RECT 2910.105 2893.995 2910.275 2894.165 ;
        RECT 2912.865 2893.995 2913.035 2894.165 ;
        RECT 2913.325 2893.995 2913.495 2894.165 ;
        RECT 2913.785 2893.995 2913.955 2894.165 ;
        RECT 5.665 2888.555 5.835 2888.725 ;
        RECT 6.125 2888.555 6.295 2888.725 ;
        RECT 6.585 2888.555 6.755 2888.725 ;
        RECT 2910.105 2888.555 2910.275 2888.725 ;
        RECT 2912.865 2888.555 2913.035 2888.725 ;
        RECT 2913.325 2888.555 2913.495 2888.725 ;
        RECT 2913.785 2888.555 2913.955 2888.725 ;
        RECT 5.665 2883.115 5.835 2883.285 ;
        RECT 6.125 2883.115 6.295 2883.285 ;
        RECT 6.585 2883.115 6.755 2883.285 ;
        RECT 8.885 2883.115 9.055 2883.285 ;
        RECT 9.345 2883.115 9.515 2883.285 ;
        RECT 9.805 2883.115 9.975 2883.285 ;
        RECT 2910.105 2883.115 2910.275 2883.285 ;
        RECT 2912.865 2883.115 2913.035 2883.285 ;
        RECT 2913.325 2883.115 2913.495 2883.285 ;
        RECT 2913.785 2883.115 2913.955 2883.285 ;
        RECT 5.665 2877.675 5.835 2877.845 ;
        RECT 6.125 2877.675 6.295 2877.845 ;
        RECT 6.585 2877.675 6.755 2877.845 ;
        RECT 2910.105 2877.675 2910.275 2877.845 ;
        RECT 2912.865 2877.675 2913.035 2877.845 ;
        RECT 2913.325 2877.675 2913.495 2877.845 ;
        RECT 2913.785 2877.675 2913.955 2877.845 ;
        RECT 5.665 2872.235 5.835 2872.405 ;
        RECT 6.125 2872.235 6.295 2872.405 ;
        RECT 6.585 2872.235 6.755 2872.405 ;
        RECT 8.885 2872.235 9.055 2872.405 ;
        RECT 9.345 2872.235 9.515 2872.405 ;
        RECT 9.805 2872.235 9.975 2872.405 ;
        RECT 2910.105 2872.235 2910.275 2872.405 ;
        RECT 2912.865 2872.235 2913.035 2872.405 ;
        RECT 2913.325 2872.235 2913.495 2872.405 ;
        RECT 2913.785 2872.235 2913.955 2872.405 ;
        RECT 5.665 2866.795 5.835 2866.965 ;
        RECT 6.125 2866.795 6.295 2866.965 ;
        RECT 6.585 2866.795 6.755 2866.965 ;
        RECT 2910.105 2866.795 2910.275 2866.965 ;
        RECT 2912.865 2866.795 2913.035 2866.965 ;
        RECT 2913.325 2866.795 2913.495 2866.965 ;
        RECT 2913.785 2866.795 2913.955 2866.965 ;
        RECT 5.665 2861.355 5.835 2861.525 ;
        RECT 6.125 2861.355 6.295 2861.525 ;
        RECT 6.585 2861.355 6.755 2861.525 ;
        RECT 2910.105 2861.355 2910.275 2861.525 ;
        RECT 2912.865 2861.355 2913.035 2861.525 ;
        RECT 2913.325 2861.355 2913.495 2861.525 ;
        RECT 2913.785 2861.355 2913.955 2861.525 ;
        RECT 5.665 2855.915 5.835 2856.085 ;
        RECT 6.125 2855.915 6.295 2856.085 ;
        RECT 6.585 2855.915 6.755 2856.085 ;
        RECT 2910.105 2855.915 2910.275 2856.085 ;
        RECT 2912.865 2855.915 2913.035 2856.085 ;
        RECT 2913.325 2855.915 2913.495 2856.085 ;
        RECT 2913.785 2855.915 2913.955 2856.085 ;
        RECT 5.665 2850.475 5.835 2850.645 ;
        RECT 6.125 2850.475 6.295 2850.645 ;
        RECT 6.585 2850.475 6.755 2850.645 ;
        RECT 2910.105 2850.475 2910.275 2850.645 ;
        RECT 2912.865 2850.475 2913.035 2850.645 ;
        RECT 2913.325 2850.475 2913.495 2850.645 ;
        RECT 2913.785 2850.475 2913.955 2850.645 ;
        RECT 5.665 2845.035 5.835 2845.205 ;
        RECT 6.125 2845.035 6.295 2845.205 ;
        RECT 6.585 2845.035 6.755 2845.205 ;
        RECT 2910.105 2845.035 2910.275 2845.205 ;
        RECT 2912.865 2845.035 2913.035 2845.205 ;
        RECT 2913.325 2845.035 2913.495 2845.205 ;
        RECT 2913.785 2845.035 2913.955 2845.205 ;
        RECT 5.665 2839.595 5.835 2839.765 ;
        RECT 6.125 2839.595 6.295 2839.765 ;
        RECT 6.585 2839.595 6.755 2839.765 ;
        RECT 2910.105 2839.595 2910.275 2839.765 ;
        RECT 2912.865 2839.595 2913.035 2839.765 ;
        RECT 2913.325 2839.595 2913.495 2839.765 ;
        RECT 2913.785 2839.595 2913.955 2839.765 ;
        RECT 5.665 2834.155 5.835 2834.325 ;
        RECT 6.125 2834.155 6.295 2834.325 ;
        RECT 6.585 2834.155 6.755 2834.325 ;
        RECT 2910.105 2834.155 2910.275 2834.325 ;
        RECT 2912.865 2834.155 2913.035 2834.325 ;
        RECT 2913.325 2834.155 2913.495 2834.325 ;
        RECT 2913.785 2834.155 2913.955 2834.325 ;
        RECT 5.665 2828.715 5.835 2828.885 ;
        RECT 6.125 2828.715 6.295 2828.885 ;
        RECT 6.585 2828.715 6.755 2828.885 ;
        RECT 2910.105 2828.715 2910.275 2828.885 ;
        RECT 2912.865 2828.715 2913.035 2828.885 ;
        RECT 2913.325 2828.715 2913.495 2828.885 ;
        RECT 2913.785 2828.715 2913.955 2828.885 ;
        RECT 5.665 2823.275 5.835 2823.445 ;
        RECT 6.125 2823.275 6.295 2823.445 ;
        RECT 6.585 2823.275 6.755 2823.445 ;
        RECT 2910.105 2823.275 2910.275 2823.445 ;
        RECT 2912.865 2823.275 2913.035 2823.445 ;
        RECT 2913.325 2823.275 2913.495 2823.445 ;
        RECT 2913.785 2823.275 2913.955 2823.445 ;
        RECT 5.665 2817.835 5.835 2818.005 ;
        RECT 6.125 2817.835 6.295 2818.005 ;
        RECT 6.585 2817.835 6.755 2818.005 ;
        RECT 2910.105 2817.835 2910.275 2818.005 ;
        RECT 2912.865 2817.835 2913.035 2818.005 ;
        RECT 2913.325 2817.835 2913.495 2818.005 ;
        RECT 2913.785 2817.835 2913.955 2818.005 ;
        RECT 5.665 2812.395 5.835 2812.565 ;
        RECT 6.125 2812.395 6.295 2812.565 ;
        RECT 6.585 2812.395 6.755 2812.565 ;
        RECT 2910.105 2812.395 2910.275 2812.565 ;
        RECT 2912.865 2812.395 2913.035 2812.565 ;
        RECT 2913.325 2812.395 2913.495 2812.565 ;
        RECT 2913.785 2812.395 2913.955 2812.565 ;
        RECT 5.665 2806.955 5.835 2807.125 ;
        RECT 6.125 2806.955 6.295 2807.125 ;
        RECT 6.585 2806.955 6.755 2807.125 ;
        RECT 2910.105 2806.955 2910.275 2807.125 ;
        RECT 2912.865 2806.955 2913.035 2807.125 ;
        RECT 2913.325 2806.955 2913.495 2807.125 ;
        RECT 2913.785 2806.955 2913.955 2807.125 ;
        RECT 5.665 2801.515 5.835 2801.685 ;
        RECT 6.125 2801.515 6.295 2801.685 ;
        RECT 6.585 2801.515 6.755 2801.685 ;
        RECT 2910.105 2801.515 2910.275 2801.685 ;
        RECT 2912.865 2801.515 2913.035 2801.685 ;
        RECT 2913.325 2801.515 2913.495 2801.685 ;
        RECT 2913.785 2801.515 2913.955 2801.685 ;
        RECT 5.665 2796.075 5.835 2796.245 ;
        RECT 6.125 2796.075 6.295 2796.245 ;
        RECT 6.585 2796.075 6.755 2796.245 ;
        RECT 2910.105 2796.075 2910.275 2796.245 ;
        RECT 2912.865 2796.075 2913.035 2796.245 ;
        RECT 2913.325 2796.075 2913.495 2796.245 ;
        RECT 2913.785 2796.075 2913.955 2796.245 ;
        RECT 5.665 2790.635 5.835 2790.805 ;
        RECT 6.125 2790.635 6.295 2790.805 ;
        RECT 6.585 2790.635 6.755 2790.805 ;
        RECT 2910.105 2790.635 2910.275 2790.805 ;
        RECT 2912.865 2790.635 2913.035 2790.805 ;
        RECT 2913.325 2790.635 2913.495 2790.805 ;
        RECT 2913.785 2790.635 2913.955 2790.805 ;
        RECT 5.665 2785.195 5.835 2785.365 ;
        RECT 6.125 2785.195 6.295 2785.365 ;
        RECT 6.585 2785.195 6.755 2785.365 ;
        RECT 2910.105 2785.195 2910.275 2785.365 ;
        RECT 2912.865 2785.195 2913.035 2785.365 ;
        RECT 2913.325 2785.195 2913.495 2785.365 ;
        RECT 2913.785 2785.195 2913.955 2785.365 ;
        RECT 5.665 2779.755 5.835 2779.925 ;
        RECT 6.125 2779.755 6.295 2779.925 ;
        RECT 6.585 2779.755 6.755 2779.925 ;
        RECT 2910.105 2779.755 2910.275 2779.925 ;
        RECT 2912.865 2779.755 2913.035 2779.925 ;
        RECT 2913.325 2779.755 2913.495 2779.925 ;
        RECT 2913.785 2779.755 2913.955 2779.925 ;
        RECT 5.665 2774.315 5.835 2774.485 ;
        RECT 6.125 2774.315 6.295 2774.485 ;
        RECT 6.585 2774.315 6.755 2774.485 ;
        RECT 2909.185 2774.315 2909.355 2774.485 ;
        RECT 2909.645 2774.315 2909.815 2774.485 ;
        RECT 2910.105 2774.315 2910.275 2774.485 ;
        RECT 2912.865 2774.315 2913.035 2774.485 ;
        RECT 2913.325 2774.315 2913.495 2774.485 ;
        RECT 2913.785 2774.315 2913.955 2774.485 ;
        RECT 5.665 2768.875 5.835 2769.045 ;
        RECT 6.125 2768.875 6.295 2769.045 ;
        RECT 6.585 2768.875 6.755 2769.045 ;
        RECT 2910.105 2768.875 2910.275 2769.045 ;
        RECT 2912.865 2768.875 2913.035 2769.045 ;
        RECT 2913.325 2768.875 2913.495 2769.045 ;
        RECT 2913.785 2768.875 2913.955 2769.045 ;
        RECT 5.665 2763.435 5.835 2763.605 ;
        RECT 6.125 2763.435 6.295 2763.605 ;
        RECT 6.585 2763.435 6.755 2763.605 ;
        RECT 2910.105 2763.435 2910.275 2763.605 ;
        RECT 2912.865 2763.435 2913.035 2763.605 ;
        RECT 2913.325 2763.435 2913.495 2763.605 ;
        RECT 2913.785 2763.435 2913.955 2763.605 ;
        RECT 5.665 2757.995 5.835 2758.165 ;
        RECT 6.125 2757.995 6.295 2758.165 ;
        RECT 6.585 2757.995 6.755 2758.165 ;
        RECT 2910.105 2757.995 2910.275 2758.165 ;
        RECT 2912.865 2757.995 2913.035 2758.165 ;
        RECT 2913.325 2757.995 2913.495 2758.165 ;
        RECT 2913.785 2757.995 2913.955 2758.165 ;
        RECT 5.665 2752.555 5.835 2752.725 ;
        RECT 6.125 2752.555 6.295 2752.725 ;
        RECT 6.585 2752.555 6.755 2752.725 ;
        RECT 2910.105 2752.555 2910.275 2752.725 ;
        RECT 2912.865 2752.555 2913.035 2752.725 ;
        RECT 2913.325 2752.555 2913.495 2752.725 ;
        RECT 2913.785 2752.555 2913.955 2752.725 ;
        RECT 5.665 2747.115 5.835 2747.285 ;
        RECT 6.125 2747.115 6.295 2747.285 ;
        RECT 6.585 2747.115 6.755 2747.285 ;
        RECT 2910.105 2747.115 2910.275 2747.285 ;
        RECT 2912.865 2747.115 2913.035 2747.285 ;
        RECT 2913.325 2747.115 2913.495 2747.285 ;
        RECT 2913.785 2747.115 2913.955 2747.285 ;
        RECT 5.665 2741.675 5.835 2741.845 ;
        RECT 6.125 2741.675 6.295 2741.845 ;
        RECT 6.585 2741.675 6.755 2741.845 ;
        RECT 2910.105 2741.675 2910.275 2741.845 ;
        RECT 2912.865 2741.675 2913.035 2741.845 ;
        RECT 2913.325 2741.675 2913.495 2741.845 ;
        RECT 2913.785 2741.675 2913.955 2741.845 ;
        RECT 5.665 2736.235 5.835 2736.405 ;
        RECT 6.125 2736.235 6.295 2736.405 ;
        RECT 6.585 2736.235 6.755 2736.405 ;
        RECT 2910.105 2736.235 2910.275 2736.405 ;
        RECT 2912.865 2736.235 2913.035 2736.405 ;
        RECT 2913.325 2736.235 2913.495 2736.405 ;
        RECT 2913.785 2736.235 2913.955 2736.405 ;
        RECT 5.665 2730.795 5.835 2730.965 ;
        RECT 6.125 2730.795 6.295 2730.965 ;
        RECT 6.585 2730.795 6.755 2730.965 ;
        RECT 2910.105 2730.795 2910.275 2730.965 ;
        RECT 2912.865 2730.795 2913.035 2730.965 ;
        RECT 2913.325 2730.795 2913.495 2730.965 ;
        RECT 2913.785 2730.795 2913.955 2730.965 ;
        RECT 5.665 2725.355 5.835 2725.525 ;
        RECT 6.125 2725.355 6.295 2725.525 ;
        RECT 6.585 2725.355 6.755 2725.525 ;
        RECT 2910.105 2725.355 2910.275 2725.525 ;
        RECT 2912.865 2725.355 2913.035 2725.525 ;
        RECT 2913.325 2725.355 2913.495 2725.525 ;
        RECT 2913.785 2725.355 2913.955 2725.525 ;
        RECT 5.665 2719.915 5.835 2720.085 ;
        RECT 6.125 2719.915 6.295 2720.085 ;
        RECT 6.585 2719.915 6.755 2720.085 ;
        RECT 2910.105 2719.915 2910.275 2720.085 ;
        RECT 2912.865 2719.915 2913.035 2720.085 ;
        RECT 2913.325 2719.915 2913.495 2720.085 ;
        RECT 2913.785 2719.915 2913.955 2720.085 ;
        RECT 5.665 2714.475 5.835 2714.645 ;
        RECT 6.125 2714.475 6.295 2714.645 ;
        RECT 6.585 2714.475 6.755 2714.645 ;
        RECT 2910.105 2714.475 2910.275 2714.645 ;
        RECT 2912.865 2714.475 2913.035 2714.645 ;
        RECT 2913.325 2714.475 2913.495 2714.645 ;
        RECT 2913.785 2714.475 2913.955 2714.645 ;
        RECT 5.665 2709.035 5.835 2709.205 ;
        RECT 6.125 2709.035 6.295 2709.205 ;
        RECT 6.585 2709.035 6.755 2709.205 ;
        RECT 2910.105 2709.035 2910.275 2709.205 ;
        RECT 2912.865 2709.035 2913.035 2709.205 ;
        RECT 2913.325 2709.035 2913.495 2709.205 ;
        RECT 2913.785 2709.035 2913.955 2709.205 ;
        RECT 5.665 2703.595 5.835 2703.765 ;
        RECT 6.125 2703.595 6.295 2703.765 ;
        RECT 6.585 2703.595 6.755 2703.765 ;
        RECT 2910.105 2703.595 2910.275 2703.765 ;
        RECT 2912.865 2703.595 2913.035 2703.765 ;
        RECT 2913.325 2703.595 2913.495 2703.765 ;
        RECT 2913.785 2703.595 2913.955 2703.765 ;
        RECT 5.665 2698.155 5.835 2698.325 ;
        RECT 6.125 2698.155 6.295 2698.325 ;
        RECT 6.585 2698.155 6.755 2698.325 ;
        RECT 2910.105 2698.155 2910.275 2698.325 ;
        RECT 2912.865 2698.155 2913.035 2698.325 ;
        RECT 2913.325 2698.155 2913.495 2698.325 ;
        RECT 2913.785 2698.155 2913.955 2698.325 ;
        RECT 5.665 2692.715 5.835 2692.885 ;
        RECT 6.125 2692.715 6.295 2692.885 ;
        RECT 6.585 2692.715 6.755 2692.885 ;
        RECT 2912.865 2692.715 2913.035 2692.885 ;
        RECT 2913.325 2692.715 2913.495 2692.885 ;
        RECT 2913.785 2692.715 2913.955 2692.885 ;
        RECT 5.665 2687.275 5.835 2687.445 ;
        RECT 6.125 2687.275 6.295 2687.445 ;
        RECT 6.585 2687.275 6.755 2687.445 ;
        RECT 2906.425 2687.275 2906.595 2687.445 ;
        RECT 2912.865 2687.275 2913.035 2687.445 ;
        RECT 2913.325 2687.275 2913.495 2687.445 ;
        RECT 2913.785 2687.275 2913.955 2687.445 ;
        RECT 5.665 2681.835 5.835 2682.005 ;
        RECT 6.125 2681.835 6.295 2682.005 ;
        RECT 6.585 2681.835 6.755 2682.005 ;
        RECT 2906.425 2681.835 2906.595 2682.005 ;
        RECT 2912.865 2681.835 2913.035 2682.005 ;
        RECT 2913.325 2681.835 2913.495 2682.005 ;
        RECT 2913.785 2681.835 2913.955 2682.005 ;
        RECT 5.665 2676.395 5.835 2676.565 ;
        RECT 6.125 2676.395 6.295 2676.565 ;
        RECT 6.585 2676.395 6.755 2676.565 ;
        RECT 2906.425 2676.395 2906.595 2676.565 ;
        RECT 2912.865 2676.395 2913.035 2676.565 ;
        RECT 2913.325 2676.395 2913.495 2676.565 ;
        RECT 2913.785 2676.395 2913.955 2676.565 ;
        RECT 5.665 2670.955 5.835 2671.125 ;
        RECT 6.125 2670.955 6.295 2671.125 ;
        RECT 6.585 2670.955 6.755 2671.125 ;
        RECT 2906.425 2670.955 2906.595 2671.125 ;
        RECT 2912.865 2670.955 2913.035 2671.125 ;
        RECT 2913.325 2670.955 2913.495 2671.125 ;
        RECT 2913.785 2670.955 2913.955 2671.125 ;
        RECT 5.665 2665.515 5.835 2665.685 ;
        RECT 6.125 2665.515 6.295 2665.685 ;
        RECT 6.585 2665.515 6.755 2665.685 ;
        RECT 2906.425 2665.515 2906.595 2665.685 ;
        RECT 2912.865 2665.515 2913.035 2665.685 ;
        RECT 2913.325 2665.515 2913.495 2665.685 ;
        RECT 2913.785 2665.515 2913.955 2665.685 ;
        RECT 5.665 2660.075 5.835 2660.245 ;
        RECT 6.125 2660.075 6.295 2660.245 ;
        RECT 6.585 2660.075 6.755 2660.245 ;
        RECT 2906.425 2660.075 2906.595 2660.245 ;
        RECT 2912.865 2660.075 2913.035 2660.245 ;
        RECT 2913.325 2660.075 2913.495 2660.245 ;
        RECT 2913.785 2660.075 2913.955 2660.245 ;
        RECT 5.665 2654.635 5.835 2654.805 ;
        RECT 6.125 2654.635 6.295 2654.805 ;
        RECT 6.585 2654.635 6.755 2654.805 ;
        RECT 2906.425 2654.635 2906.595 2654.805 ;
        RECT 2912.865 2654.635 2913.035 2654.805 ;
        RECT 2913.325 2654.635 2913.495 2654.805 ;
        RECT 2913.785 2654.635 2913.955 2654.805 ;
        RECT 5.665 2649.195 5.835 2649.365 ;
        RECT 6.125 2649.195 6.295 2649.365 ;
        RECT 6.585 2649.195 6.755 2649.365 ;
        RECT 2906.425 2649.195 2906.595 2649.365 ;
        RECT 2912.865 2649.195 2913.035 2649.365 ;
        RECT 2913.325 2649.195 2913.495 2649.365 ;
        RECT 2913.785 2649.195 2913.955 2649.365 ;
        RECT 5.665 2643.755 5.835 2643.925 ;
        RECT 6.125 2643.755 6.295 2643.925 ;
        RECT 6.585 2643.755 6.755 2643.925 ;
        RECT 2906.425 2643.755 2906.595 2643.925 ;
        RECT 2912.865 2643.755 2913.035 2643.925 ;
        RECT 2913.325 2643.755 2913.495 2643.925 ;
        RECT 2913.785 2643.755 2913.955 2643.925 ;
        RECT 5.665 2638.315 5.835 2638.485 ;
        RECT 6.125 2638.315 6.295 2638.485 ;
        RECT 6.585 2638.315 6.755 2638.485 ;
        RECT 2906.425 2638.315 2906.595 2638.485 ;
        RECT 2912.865 2638.315 2913.035 2638.485 ;
        RECT 2913.325 2638.315 2913.495 2638.485 ;
        RECT 2913.785 2638.315 2913.955 2638.485 ;
        RECT 5.665 2632.875 5.835 2633.045 ;
        RECT 6.125 2632.875 6.295 2633.045 ;
        RECT 6.585 2632.875 6.755 2633.045 ;
        RECT 2906.425 2632.875 2906.595 2633.045 ;
        RECT 2912.865 2632.875 2913.035 2633.045 ;
        RECT 2913.325 2632.875 2913.495 2633.045 ;
        RECT 2913.785 2632.875 2913.955 2633.045 ;
        RECT 5.665 2627.435 5.835 2627.605 ;
        RECT 6.125 2627.435 6.295 2627.605 ;
        RECT 6.585 2627.435 6.755 2627.605 ;
        RECT 2906.425 2627.435 2906.595 2627.605 ;
        RECT 2909.185 2627.435 2909.355 2627.605 ;
        RECT 2909.645 2627.435 2909.815 2627.605 ;
        RECT 2910.105 2627.435 2910.275 2627.605 ;
        RECT 2912.865 2627.435 2913.035 2627.605 ;
        RECT 2913.325 2627.435 2913.495 2627.605 ;
        RECT 2913.785 2627.435 2913.955 2627.605 ;
        RECT 5.665 2621.995 5.835 2622.165 ;
        RECT 6.125 2621.995 6.295 2622.165 ;
        RECT 6.585 2621.995 6.755 2622.165 ;
        RECT 2906.425 2621.995 2906.595 2622.165 ;
        RECT 2912.865 2621.995 2913.035 2622.165 ;
        RECT 2913.325 2621.995 2913.495 2622.165 ;
        RECT 2913.785 2621.995 2913.955 2622.165 ;
        RECT 5.665 2616.555 5.835 2616.725 ;
        RECT 6.125 2616.555 6.295 2616.725 ;
        RECT 6.585 2616.555 6.755 2616.725 ;
        RECT 2906.425 2616.555 2906.595 2616.725 ;
        RECT 2912.865 2616.555 2913.035 2616.725 ;
        RECT 2913.325 2616.555 2913.495 2616.725 ;
        RECT 2913.785 2616.555 2913.955 2616.725 ;
        RECT 5.665 2611.115 5.835 2611.285 ;
        RECT 6.125 2611.115 6.295 2611.285 ;
        RECT 6.585 2611.115 6.755 2611.285 ;
        RECT 2906.425 2611.115 2906.595 2611.285 ;
        RECT 2912.865 2611.115 2913.035 2611.285 ;
        RECT 2913.325 2611.115 2913.495 2611.285 ;
        RECT 2913.785 2611.115 2913.955 2611.285 ;
        RECT 5.665 2605.675 5.835 2605.845 ;
        RECT 6.125 2605.675 6.295 2605.845 ;
        RECT 6.585 2605.675 6.755 2605.845 ;
        RECT 2906.425 2605.675 2906.595 2605.845 ;
        RECT 2912.865 2605.675 2913.035 2605.845 ;
        RECT 2913.325 2605.675 2913.495 2605.845 ;
        RECT 2913.785 2605.675 2913.955 2605.845 ;
        RECT 5.665 2600.235 5.835 2600.405 ;
        RECT 6.125 2600.235 6.295 2600.405 ;
        RECT 6.585 2600.235 6.755 2600.405 ;
        RECT 2906.425 2600.235 2906.595 2600.405 ;
        RECT 2909.185 2600.235 2909.355 2600.405 ;
        RECT 2909.645 2600.235 2909.815 2600.405 ;
        RECT 2910.105 2600.235 2910.275 2600.405 ;
        RECT 2912.865 2600.235 2913.035 2600.405 ;
        RECT 2913.325 2600.235 2913.495 2600.405 ;
        RECT 2913.785 2600.235 2913.955 2600.405 ;
        RECT 5.665 2594.795 5.835 2594.965 ;
        RECT 6.125 2594.795 6.295 2594.965 ;
        RECT 6.585 2594.795 6.755 2594.965 ;
        RECT 2906.425 2594.795 2906.595 2594.965 ;
        RECT 2912.865 2594.795 2913.035 2594.965 ;
        RECT 2913.325 2594.795 2913.495 2594.965 ;
        RECT 2913.785 2594.795 2913.955 2594.965 ;
        RECT 5.665 2589.355 5.835 2589.525 ;
        RECT 6.125 2589.355 6.295 2589.525 ;
        RECT 6.585 2589.355 6.755 2589.525 ;
        RECT 2906.425 2589.355 2906.595 2589.525 ;
        RECT 2912.865 2589.355 2913.035 2589.525 ;
        RECT 2913.325 2589.355 2913.495 2589.525 ;
        RECT 2913.785 2589.355 2913.955 2589.525 ;
        RECT 5.665 2583.915 5.835 2584.085 ;
        RECT 6.125 2583.915 6.295 2584.085 ;
        RECT 6.585 2583.915 6.755 2584.085 ;
        RECT 2906.425 2583.915 2906.595 2584.085 ;
        RECT 2912.865 2583.915 2913.035 2584.085 ;
        RECT 2913.325 2583.915 2913.495 2584.085 ;
        RECT 2913.785 2583.915 2913.955 2584.085 ;
        RECT 5.665 2578.475 5.835 2578.645 ;
        RECT 6.125 2578.475 6.295 2578.645 ;
        RECT 6.585 2578.475 6.755 2578.645 ;
        RECT 2906.425 2578.475 2906.595 2578.645 ;
        RECT 2912.865 2578.475 2913.035 2578.645 ;
        RECT 2913.325 2578.475 2913.495 2578.645 ;
        RECT 2913.785 2578.475 2913.955 2578.645 ;
        RECT 5.665 2573.035 5.835 2573.205 ;
        RECT 6.125 2573.035 6.295 2573.205 ;
        RECT 6.585 2573.035 6.755 2573.205 ;
        RECT 2906.425 2573.035 2906.595 2573.205 ;
        RECT 2912.865 2573.035 2913.035 2573.205 ;
        RECT 2913.325 2573.035 2913.495 2573.205 ;
        RECT 2913.785 2573.035 2913.955 2573.205 ;
        RECT 5.665 2567.595 5.835 2567.765 ;
        RECT 6.125 2567.595 6.295 2567.765 ;
        RECT 6.585 2567.595 6.755 2567.765 ;
        RECT 2906.425 2567.595 2906.595 2567.765 ;
        RECT 2912.865 2567.595 2913.035 2567.765 ;
        RECT 2913.325 2567.595 2913.495 2567.765 ;
        RECT 2913.785 2567.595 2913.955 2567.765 ;
        RECT 5.665 2562.155 5.835 2562.325 ;
        RECT 6.125 2562.155 6.295 2562.325 ;
        RECT 6.585 2562.155 6.755 2562.325 ;
        RECT 2906.425 2562.155 2906.595 2562.325 ;
        RECT 2912.865 2562.155 2913.035 2562.325 ;
        RECT 2913.325 2562.155 2913.495 2562.325 ;
        RECT 2913.785 2562.155 2913.955 2562.325 ;
        RECT 5.665 2556.715 5.835 2556.885 ;
        RECT 6.125 2556.715 6.295 2556.885 ;
        RECT 6.585 2556.715 6.755 2556.885 ;
        RECT 2906.425 2556.715 2906.595 2556.885 ;
        RECT 2912.865 2556.715 2913.035 2556.885 ;
        RECT 2913.325 2556.715 2913.495 2556.885 ;
        RECT 2913.785 2556.715 2913.955 2556.885 ;
        RECT 5.665 2551.275 5.835 2551.445 ;
        RECT 6.125 2551.275 6.295 2551.445 ;
        RECT 6.585 2551.275 6.755 2551.445 ;
        RECT 2906.425 2551.275 2906.595 2551.445 ;
        RECT 2912.865 2551.275 2913.035 2551.445 ;
        RECT 2913.325 2551.275 2913.495 2551.445 ;
        RECT 2913.785 2551.275 2913.955 2551.445 ;
        RECT 5.665 2545.835 5.835 2546.005 ;
        RECT 6.125 2545.835 6.295 2546.005 ;
        RECT 6.585 2545.835 6.755 2546.005 ;
        RECT 2906.425 2545.835 2906.595 2546.005 ;
        RECT 2912.865 2545.835 2913.035 2546.005 ;
        RECT 2913.325 2545.835 2913.495 2546.005 ;
        RECT 2913.785 2545.835 2913.955 2546.005 ;
        RECT 5.665 2540.395 5.835 2540.565 ;
        RECT 6.125 2540.395 6.295 2540.565 ;
        RECT 6.585 2540.395 6.755 2540.565 ;
        RECT 2906.425 2540.395 2906.595 2540.565 ;
        RECT 2912.865 2540.395 2913.035 2540.565 ;
        RECT 2913.325 2540.395 2913.495 2540.565 ;
        RECT 2913.785 2540.395 2913.955 2540.565 ;
        RECT 5.665 2534.955 5.835 2535.125 ;
        RECT 6.125 2534.955 6.295 2535.125 ;
        RECT 6.585 2534.955 6.755 2535.125 ;
        RECT 2906.425 2534.955 2906.595 2535.125 ;
        RECT 2912.865 2534.955 2913.035 2535.125 ;
        RECT 2913.325 2534.955 2913.495 2535.125 ;
        RECT 2913.785 2534.955 2913.955 2535.125 ;
        RECT 5.665 2529.515 5.835 2529.685 ;
        RECT 6.125 2529.515 6.295 2529.685 ;
        RECT 6.585 2529.515 6.755 2529.685 ;
        RECT 2906.425 2529.515 2906.595 2529.685 ;
        RECT 2912.865 2529.515 2913.035 2529.685 ;
        RECT 2913.325 2529.515 2913.495 2529.685 ;
        RECT 2913.785 2529.515 2913.955 2529.685 ;
        RECT 5.665 2524.075 5.835 2524.245 ;
        RECT 6.125 2524.075 6.295 2524.245 ;
        RECT 6.585 2524.075 6.755 2524.245 ;
        RECT 2906.425 2524.075 2906.595 2524.245 ;
        RECT 2912.865 2524.075 2913.035 2524.245 ;
        RECT 2913.325 2524.075 2913.495 2524.245 ;
        RECT 2913.785 2524.075 2913.955 2524.245 ;
        RECT 5.665 2518.635 5.835 2518.805 ;
        RECT 6.125 2518.635 6.295 2518.805 ;
        RECT 6.585 2518.635 6.755 2518.805 ;
        RECT 2906.425 2518.635 2906.595 2518.805 ;
        RECT 2912.865 2518.635 2913.035 2518.805 ;
        RECT 2913.325 2518.635 2913.495 2518.805 ;
        RECT 2913.785 2518.635 2913.955 2518.805 ;
        RECT 5.665 2513.195 5.835 2513.365 ;
        RECT 6.125 2513.195 6.295 2513.365 ;
        RECT 6.585 2513.195 6.755 2513.365 ;
        RECT 2906.425 2513.195 2906.595 2513.365 ;
        RECT 2912.865 2513.195 2913.035 2513.365 ;
        RECT 2913.325 2513.195 2913.495 2513.365 ;
        RECT 2913.785 2513.195 2913.955 2513.365 ;
        RECT 5.665 2507.755 5.835 2507.925 ;
        RECT 6.125 2507.755 6.295 2507.925 ;
        RECT 6.585 2507.755 6.755 2507.925 ;
        RECT 2906.425 2507.755 2906.595 2507.925 ;
        RECT 2912.865 2507.755 2913.035 2507.925 ;
        RECT 2913.325 2507.755 2913.495 2507.925 ;
        RECT 2913.785 2507.755 2913.955 2507.925 ;
        RECT 5.665 2502.315 5.835 2502.485 ;
        RECT 6.125 2502.315 6.295 2502.485 ;
        RECT 6.585 2502.315 6.755 2502.485 ;
        RECT 8.885 2502.315 9.055 2502.485 ;
        RECT 9.345 2502.315 9.515 2502.485 ;
        RECT 9.805 2502.315 9.975 2502.485 ;
        RECT 2906.425 2502.315 2906.595 2502.485 ;
        RECT 2912.865 2502.315 2913.035 2502.485 ;
        RECT 2913.325 2502.315 2913.495 2502.485 ;
        RECT 2913.785 2502.315 2913.955 2502.485 ;
        RECT 5.665 2496.875 5.835 2497.045 ;
        RECT 6.125 2496.875 6.295 2497.045 ;
        RECT 6.585 2496.875 6.755 2497.045 ;
        RECT 2906.425 2496.875 2906.595 2497.045 ;
        RECT 2912.865 2496.875 2913.035 2497.045 ;
        RECT 2913.325 2496.875 2913.495 2497.045 ;
        RECT 2913.785 2496.875 2913.955 2497.045 ;
        RECT 5.665 2491.435 5.835 2491.605 ;
        RECT 6.125 2491.435 6.295 2491.605 ;
        RECT 6.585 2491.435 6.755 2491.605 ;
        RECT 2906.425 2491.435 2906.595 2491.605 ;
        RECT 2912.865 2491.435 2913.035 2491.605 ;
        RECT 2913.325 2491.435 2913.495 2491.605 ;
        RECT 2913.785 2491.435 2913.955 2491.605 ;
        RECT 5.665 2485.995 5.835 2486.165 ;
        RECT 6.125 2485.995 6.295 2486.165 ;
        RECT 6.585 2485.995 6.755 2486.165 ;
        RECT 2906.425 2485.995 2906.595 2486.165 ;
        RECT 2912.865 2485.995 2913.035 2486.165 ;
        RECT 2913.325 2485.995 2913.495 2486.165 ;
        RECT 2913.785 2485.995 2913.955 2486.165 ;
        RECT 5.665 2480.555 5.835 2480.725 ;
        RECT 6.125 2480.555 6.295 2480.725 ;
        RECT 6.585 2480.555 6.755 2480.725 ;
        RECT 2906.425 2480.555 2906.595 2480.725 ;
        RECT 2912.865 2480.555 2913.035 2480.725 ;
        RECT 2913.325 2480.555 2913.495 2480.725 ;
        RECT 2913.785 2480.555 2913.955 2480.725 ;
        RECT 5.665 2475.115 5.835 2475.285 ;
        RECT 6.125 2475.115 6.295 2475.285 ;
        RECT 6.585 2475.115 6.755 2475.285 ;
        RECT 2906.425 2475.115 2906.595 2475.285 ;
        RECT 2912.865 2475.115 2913.035 2475.285 ;
        RECT 2913.325 2475.115 2913.495 2475.285 ;
        RECT 2913.785 2475.115 2913.955 2475.285 ;
        RECT 5.665 2469.675 5.835 2469.845 ;
        RECT 6.125 2469.675 6.295 2469.845 ;
        RECT 6.585 2469.675 6.755 2469.845 ;
        RECT 2906.425 2469.675 2906.595 2469.845 ;
        RECT 2912.865 2469.675 2913.035 2469.845 ;
        RECT 2913.325 2469.675 2913.495 2469.845 ;
        RECT 2913.785 2469.675 2913.955 2469.845 ;
        RECT 5.665 2464.235 5.835 2464.405 ;
        RECT 6.125 2464.235 6.295 2464.405 ;
        RECT 6.585 2464.235 6.755 2464.405 ;
        RECT 2906.425 2464.235 2906.595 2464.405 ;
        RECT 2909.185 2464.235 2909.355 2464.405 ;
        RECT 2909.645 2464.235 2909.815 2464.405 ;
        RECT 2910.105 2464.235 2910.275 2464.405 ;
        RECT 2912.865 2464.235 2913.035 2464.405 ;
        RECT 2913.325 2464.235 2913.495 2464.405 ;
        RECT 2913.785 2464.235 2913.955 2464.405 ;
        RECT 5.665 2458.795 5.835 2458.965 ;
        RECT 6.125 2458.795 6.295 2458.965 ;
        RECT 6.585 2458.795 6.755 2458.965 ;
        RECT 2906.425 2458.795 2906.595 2458.965 ;
        RECT 2912.865 2458.795 2913.035 2458.965 ;
        RECT 2913.325 2458.795 2913.495 2458.965 ;
        RECT 2913.785 2458.795 2913.955 2458.965 ;
        RECT 5.665 2453.355 5.835 2453.525 ;
        RECT 6.125 2453.355 6.295 2453.525 ;
        RECT 6.585 2453.355 6.755 2453.525 ;
        RECT 2906.425 2453.355 2906.595 2453.525 ;
        RECT 2912.865 2453.355 2913.035 2453.525 ;
        RECT 2913.325 2453.355 2913.495 2453.525 ;
        RECT 2913.785 2453.355 2913.955 2453.525 ;
        RECT 5.665 2447.915 5.835 2448.085 ;
        RECT 6.125 2447.915 6.295 2448.085 ;
        RECT 6.585 2447.915 6.755 2448.085 ;
        RECT 2906.425 2447.915 2906.595 2448.085 ;
        RECT 2912.865 2447.915 2913.035 2448.085 ;
        RECT 2913.325 2447.915 2913.495 2448.085 ;
        RECT 2913.785 2447.915 2913.955 2448.085 ;
        RECT 5.665 2442.475 5.835 2442.645 ;
        RECT 6.125 2442.475 6.295 2442.645 ;
        RECT 6.585 2442.475 6.755 2442.645 ;
        RECT 2906.425 2442.475 2906.595 2442.645 ;
        RECT 2912.865 2442.475 2913.035 2442.645 ;
        RECT 2913.325 2442.475 2913.495 2442.645 ;
        RECT 2913.785 2442.475 2913.955 2442.645 ;
        RECT 5.665 2437.035 5.835 2437.205 ;
        RECT 6.125 2437.035 6.295 2437.205 ;
        RECT 6.585 2437.035 6.755 2437.205 ;
        RECT 2906.425 2437.035 2906.595 2437.205 ;
        RECT 2912.865 2437.035 2913.035 2437.205 ;
        RECT 2913.325 2437.035 2913.495 2437.205 ;
        RECT 2913.785 2437.035 2913.955 2437.205 ;
        RECT 5.665 2431.595 5.835 2431.765 ;
        RECT 6.125 2431.595 6.295 2431.765 ;
        RECT 6.585 2431.595 6.755 2431.765 ;
        RECT 2906.425 2431.595 2906.595 2431.765 ;
        RECT 2909.185 2431.595 2909.355 2431.765 ;
        RECT 2909.645 2431.595 2909.815 2431.765 ;
        RECT 2910.105 2431.595 2910.275 2431.765 ;
        RECT 2912.865 2431.595 2913.035 2431.765 ;
        RECT 2913.325 2431.595 2913.495 2431.765 ;
        RECT 2913.785 2431.595 2913.955 2431.765 ;
        RECT 5.665 2426.155 5.835 2426.325 ;
        RECT 6.125 2426.155 6.295 2426.325 ;
        RECT 6.585 2426.155 6.755 2426.325 ;
        RECT 2906.425 2426.155 2906.595 2426.325 ;
        RECT 2912.865 2426.155 2913.035 2426.325 ;
        RECT 2913.325 2426.155 2913.495 2426.325 ;
        RECT 2913.785 2426.155 2913.955 2426.325 ;
        RECT 5.665 2420.715 5.835 2420.885 ;
        RECT 6.125 2420.715 6.295 2420.885 ;
        RECT 6.585 2420.715 6.755 2420.885 ;
        RECT 2906.425 2420.715 2906.595 2420.885 ;
        RECT 2912.865 2420.715 2913.035 2420.885 ;
        RECT 2913.325 2420.715 2913.495 2420.885 ;
        RECT 2913.785 2420.715 2913.955 2420.885 ;
        RECT 5.665 2415.275 5.835 2415.445 ;
        RECT 6.125 2415.275 6.295 2415.445 ;
        RECT 6.585 2415.275 6.755 2415.445 ;
        RECT 2906.425 2415.275 2906.595 2415.445 ;
        RECT 2912.865 2415.275 2913.035 2415.445 ;
        RECT 2913.325 2415.275 2913.495 2415.445 ;
        RECT 2913.785 2415.275 2913.955 2415.445 ;
        RECT 5.665 2409.835 5.835 2410.005 ;
        RECT 6.125 2409.835 6.295 2410.005 ;
        RECT 6.585 2409.835 6.755 2410.005 ;
        RECT 2906.425 2409.835 2906.595 2410.005 ;
        RECT 2912.865 2409.835 2913.035 2410.005 ;
        RECT 2913.325 2409.835 2913.495 2410.005 ;
        RECT 2913.785 2409.835 2913.955 2410.005 ;
        RECT 5.665 2404.395 5.835 2404.565 ;
        RECT 6.125 2404.395 6.295 2404.565 ;
        RECT 6.585 2404.395 6.755 2404.565 ;
        RECT 2906.425 2404.395 2906.595 2404.565 ;
        RECT 2912.865 2404.395 2913.035 2404.565 ;
        RECT 2913.325 2404.395 2913.495 2404.565 ;
        RECT 2913.785 2404.395 2913.955 2404.565 ;
        RECT 5.665 2398.955 5.835 2399.125 ;
        RECT 6.125 2398.955 6.295 2399.125 ;
        RECT 6.585 2398.955 6.755 2399.125 ;
        RECT 2906.425 2398.955 2906.595 2399.125 ;
        RECT 2912.865 2398.955 2913.035 2399.125 ;
        RECT 2913.325 2398.955 2913.495 2399.125 ;
        RECT 2913.785 2398.955 2913.955 2399.125 ;
        RECT 5.665 2393.515 5.835 2393.685 ;
        RECT 6.125 2393.515 6.295 2393.685 ;
        RECT 6.585 2393.515 6.755 2393.685 ;
        RECT 2906.425 2393.515 2906.595 2393.685 ;
        RECT 2912.865 2393.515 2913.035 2393.685 ;
        RECT 2913.325 2393.515 2913.495 2393.685 ;
        RECT 2913.785 2393.515 2913.955 2393.685 ;
        RECT 5.665 2388.075 5.835 2388.245 ;
        RECT 6.125 2388.075 6.295 2388.245 ;
        RECT 6.585 2388.075 6.755 2388.245 ;
        RECT 2906.425 2388.075 2906.595 2388.245 ;
        RECT 2909.185 2388.075 2909.355 2388.245 ;
        RECT 2909.645 2388.075 2909.815 2388.245 ;
        RECT 2910.105 2388.075 2910.275 2388.245 ;
        RECT 2912.865 2388.075 2913.035 2388.245 ;
        RECT 2913.325 2388.075 2913.495 2388.245 ;
        RECT 2913.785 2388.075 2913.955 2388.245 ;
        RECT 5.665 2382.635 5.835 2382.805 ;
        RECT 6.125 2382.635 6.295 2382.805 ;
        RECT 6.585 2382.635 6.755 2382.805 ;
        RECT 8.885 2382.635 9.055 2382.805 ;
        RECT 9.345 2382.635 9.515 2382.805 ;
        RECT 9.805 2382.635 9.975 2382.805 ;
        RECT 2906.425 2382.635 2906.595 2382.805 ;
        RECT 2912.865 2382.635 2913.035 2382.805 ;
        RECT 2913.325 2382.635 2913.495 2382.805 ;
        RECT 2913.785 2382.635 2913.955 2382.805 ;
        RECT 5.665 2377.195 5.835 2377.365 ;
        RECT 6.125 2377.195 6.295 2377.365 ;
        RECT 6.585 2377.195 6.755 2377.365 ;
        RECT 2906.425 2377.195 2906.595 2377.365 ;
        RECT 2912.865 2377.195 2913.035 2377.365 ;
        RECT 2913.325 2377.195 2913.495 2377.365 ;
        RECT 2913.785 2377.195 2913.955 2377.365 ;
        RECT 5.665 2371.755 5.835 2371.925 ;
        RECT 6.125 2371.755 6.295 2371.925 ;
        RECT 6.585 2371.755 6.755 2371.925 ;
        RECT 2906.425 2371.755 2906.595 2371.925 ;
        RECT 2912.865 2371.755 2913.035 2371.925 ;
        RECT 2913.325 2371.755 2913.495 2371.925 ;
        RECT 2913.785 2371.755 2913.955 2371.925 ;
        RECT 5.665 2366.315 5.835 2366.485 ;
        RECT 6.125 2366.315 6.295 2366.485 ;
        RECT 6.585 2366.315 6.755 2366.485 ;
        RECT 2906.425 2366.315 2906.595 2366.485 ;
        RECT 2912.865 2366.315 2913.035 2366.485 ;
        RECT 2913.325 2366.315 2913.495 2366.485 ;
        RECT 2913.785 2366.315 2913.955 2366.485 ;
        RECT 5.665 2360.875 5.835 2361.045 ;
        RECT 6.125 2360.875 6.295 2361.045 ;
        RECT 6.585 2360.875 6.755 2361.045 ;
        RECT 2906.425 2360.875 2906.595 2361.045 ;
        RECT 2912.865 2360.875 2913.035 2361.045 ;
        RECT 2913.325 2360.875 2913.495 2361.045 ;
        RECT 2913.785 2360.875 2913.955 2361.045 ;
        RECT 5.665 2355.435 5.835 2355.605 ;
        RECT 6.125 2355.435 6.295 2355.605 ;
        RECT 6.585 2355.435 6.755 2355.605 ;
        RECT 2906.425 2355.435 2906.595 2355.605 ;
        RECT 2912.865 2355.435 2913.035 2355.605 ;
        RECT 2913.325 2355.435 2913.495 2355.605 ;
        RECT 2913.785 2355.435 2913.955 2355.605 ;
        RECT 5.665 2349.995 5.835 2350.165 ;
        RECT 6.125 2349.995 6.295 2350.165 ;
        RECT 6.585 2349.995 6.755 2350.165 ;
        RECT 2906.425 2349.995 2906.595 2350.165 ;
        RECT 2912.865 2349.995 2913.035 2350.165 ;
        RECT 2913.325 2349.995 2913.495 2350.165 ;
        RECT 2913.785 2349.995 2913.955 2350.165 ;
        RECT 5.665 2344.555 5.835 2344.725 ;
        RECT 6.125 2344.555 6.295 2344.725 ;
        RECT 6.585 2344.555 6.755 2344.725 ;
        RECT 2906.425 2344.555 2906.595 2344.725 ;
        RECT 2912.865 2344.555 2913.035 2344.725 ;
        RECT 2913.325 2344.555 2913.495 2344.725 ;
        RECT 2913.785 2344.555 2913.955 2344.725 ;
        RECT 5.665 2339.115 5.835 2339.285 ;
        RECT 6.125 2339.115 6.295 2339.285 ;
        RECT 6.585 2339.115 6.755 2339.285 ;
        RECT 2906.425 2339.115 2906.595 2339.285 ;
        RECT 2912.865 2339.115 2913.035 2339.285 ;
        RECT 2913.325 2339.115 2913.495 2339.285 ;
        RECT 2913.785 2339.115 2913.955 2339.285 ;
        RECT 5.665 2333.675 5.835 2333.845 ;
        RECT 6.125 2333.675 6.295 2333.845 ;
        RECT 6.585 2333.675 6.755 2333.845 ;
        RECT 2906.425 2333.675 2906.595 2333.845 ;
        RECT 2912.865 2333.675 2913.035 2333.845 ;
        RECT 2913.325 2333.675 2913.495 2333.845 ;
        RECT 2913.785 2333.675 2913.955 2333.845 ;
        RECT 5.665 2328.235 5.835 2328.405 ;
        RECT 6.125 2328.235 6.295 2328.405 ;
        RECT 6.585 2328.235 6.755 2328.405 ;
        RECT 2906.425 2328.235 2906.595 2328.405 ;
        RECT 2912.865 2328.235 2913.035 2328.405 ;
        RECT 2913.325 2328.235 2913.495 2328.405 ;
        RECT 2913.785 2328.235 2913.955 2328.405 ;
        RECT 5.665 2322.795 5.835 2322.965 ;
        RECT 6.125 2322.795 6.295 2322.965 ;
        RECT 6.585 2322.795 6.755 2322.965 ;
        RECT 2906.425 2322.795 2906.595 2322.965 ;
        RECT 2912.865 2322.795 2913.035 2322.965 ;
        RECT 2913.325 2322.795 2913.495 2322.965 ;
        RECT 2913.785 2322.795 2913.955 2322.965 ;
        RECT 5.665 2317.355 5.835 2317.525 ;
        RECT 6.125 2317.355 6.295 2317.525 ;
        RECT 6.585 2317.355 6.755 2317.525 ;
        RECT 2906.425 2317.355 2906.595 2317.525 ;
        RECT 2912.865 2317.355 2913.035 2317.525 ;
        RECT 2913.325 2317.355 2913.495 2317.525 ;
        RECT 2913.785 2317.355 2913.955 2317.525 ;
        RECT 5.665 2311.915 5.835 2312.085 ;
        RECT 6.125 2311.915 6.295 2312.085 ;
        RECT 6.585 2311.915 6.755 2312.085 ;
        RECT 2906.425 2311.915 2906.595 2312.085 ;
        RECT 2912.865 2311.915 2913.035 2312.085 ;
        RECT 2913.325 2311.915 2913.495 2312.085 ;
        RECT 2913.785 2311.915 2913.955 2312.085 ;
        RECT 5.665 2306.475 5.835 2306.645 ;
        RECT 6.125 2306.475 6.295 2306.645 ;
        RECT 6.585 2306.475 6.755 2306.645 ;
        RECT 2906.425 2306.475 2906.595 2306.645 ;
        RECT 2912.865 2306.475 2913.035 2306.645 ;
        RECT 2913.325 2306.475 2913.495 2306.645 ;
        RECT 2913.785 2306.475 2913.955 2306.645 ;
        RECT 5.665 2301.035 5.835 2301.205 ;
        RECT 6.125 2301.035 6.295 2301.205 ;
        RECT 6.585 2301.035 6.755 2301.205 ;
        RECT 2906.425 2301.035 2906.595 2301.205 ;
        RECT 2912.865 2301.035 2913.035 2301.205 ;
        RECT 2913.325 2301.035 2913.495 2301.205 ;
        RECT 2913.785 2301.035 2913.955 2301.205 ;
        RECT 5.665 2295.595 5.835 2295.765 ;
        RECT 6.125 2295.595 6.295 2295.765 ;
        RECT 6.585 2295.595 6.755 2295.765 ;
        RECT 2906.425 2295.595 2906.595 2295.765 ;
        RECT 2912.865 2295.595 2913.035 2295.765 ;
        RECT 2913.325 2295.595 2913.495 2295.765 ;
        RECT 2913.785 2295.595 2913.955 2295.765 ;
        RECT 5.665 2290.155 5.835 2290.325 ;
        RECT 6.125 2290.155 6.295 2290.325 ;
        RECT 6.585 2290.155 6.755 2290.325 ;
        RECT 2906.425 2290.155 2906.595 2290.325 ;
        RECT 2912.865 2290.155 2913.035 2290.325 ;
        RECT 2913.325 2290.155 2913.495 2290.325 ;
        RECT 2913.785 2290.155 2913.955 2290.325 ;
        RECT 5.665 2284.715 5.835 2284.885 ;
        RECT 6.125 2284.715 6.295 2284.885 ;
        RECT 6.585 2284.715 6.755 2284.885 ;
        RECT 2906.425 2284.715 2906.595 2284.885 ;
        RECT 2912.865 2284.715 2913.035 2284.885 ;
        RECT 2913.325 2284.715 2913.495 2284.885 ;
        RECT 2913.785 2284.715 2913.955 2284.885 ;
        RECT 5.665 2279.275 5.835 2279.445 ;
        RECT 6.125 2279.275 6.295 2279.445 ;
        RECT 6.585 2279.275 6.755 2279.445 ;
        RECT 2906.425 2279.275 2906.595 2279.445 ;
        RECT 2912.865 2279.275 2913.035 2279.445 ;
        RECT 2913.325 2279.275 2913.495 2279.445 ;
        RECT 2913.785 2279.275 2913.955 2279.445 ;
        RECT 5.665 2273.835 5.835 2274.005 ;
        RECT 6.125 2273.835 6.295 2274.005 ;
        RECT 6.585 2273.835 6.755 2274.005 ;
        RECT 2906.425 2273.835 2906.595 2274.005 ;
        RECT 2912.865 2273.835 2913.035 2274.005 ;
        RECT 2913.325 2273.835 2913.495 2274.005 ;
        RECT 2913.785 2273.835 2913.955 2274.005 ;
        RECT 5.665 2268.395 5.835 2268.565 ;
        RECT 6.125 2268.395 6.295 2268.565 ;
        RECT 6.585 2268.395 6.755 2268.565 ;
        RECT 2906.425 2268.395 2906.595 2268.565 ;
        RECT 2912.865 2268.395 2913.035 2268.565 ;
        RECT 2913.325 2268.395 2913.495 2268.565 ;
        RECT 2913.785 2268.395 2913.955 2268.565 ;
        RECT 5.665 2262.955 5.835 2263.125 ;
        RECT 6.125 2262.955 6.295 2263.125 ;
        RECT 6.585 2262.955 6.755 2263.125 ;
        RECT 2906.425 2262.955 2906.595 2263.125 ;
        RECT 2909.185 2262.955 2909.355 2263.125 ;
        RECT 2909.645 2262.955 2909.815 2263.125 ;
        RECT 2910.105 2262.955 2910.275 2263.125 ;
        RECT 2912.865 2262.955 2913.035 2263.125 ;
        RECT 2913.325 2262.955 2913.495 2263.125 ;
        RECT 2913.785 2262.955 2913.955 2263.125 ;
        RECT 5.665 2257.515 5.835 2257.685 ;
        RECT 6.125 2257.515 6.295 2257.685 ;
        RECT 6.585 2257.515 6.755 2257.685 ;
        RECT 2906.425 2257.515 2906.595 2257.685 ;
        RECT 2912.865 2257.515 2913.035 2257.685 ;
        RECT 2913.325 2257.515 2913.495 2257.685 ;
        RECT 2913.785 2257.515 2913.955 2257.685 ;
        RECT 5.665 2252.075 5.835 2252.245 ;
        RECT 6.125 2252.075 6.295 2252.245 ;
        RECT 6.585 2252.075 6.755 2252.245 ;
        RECT 2906.425 2252.075 2906.595 2252.245 ;
        RECT 2912.865 2252.075 2913.035 2252.245 ;
        RECT 2913.325 2252.075 2913.495 2252.245 ;
        RECT 2913.785 2252.075 2913.955 2252.245 ;
        RECT 5.665 2246.635 5.835 2246.805 ;
        RECT 6.125 2246.635 6.295 2246.805 ;
        RECT 6.585 2246.635 6.755 2246.805 ;
        RECT 2906.425 2246.635 2906.595 2246.805 ;
        RECT 2912.865 2246.635 2913.035 2246.805 ;
        RECT 2913.325 2246.635 2913.495 2246.805 ;
        RECT 2913.785 2246.635 2913.955 2246.805 ;
        RECT 5.665 2241.195 5.835 2241.365 ;
        RECT 6.125 2241.195 6.295 2241.365 ;
        RECT 6.585 2241.195 6.755 2241.365 ;
        RECT 2906.425 2241.195 2906.595 2241.365 ;
        RECT 2912.865 2241.195 2913.035 2241.365 ;
        RECT 2913.325 2241.195 2913.495 2241.365 ;
        RECT 2913.785 2241.195 2913.955 2241.365 ;
        RECT 5.665 2235.755 5.835 2235.925 ;
        RECT 6.125 2235.755 6.295 2235.925 ;
        RECT 6.585 2235.755 6.755 2235.925 ;
        RECT 2906.425 2235.755 2906.595 2235.925 ;
        RECT 2912.865 2235.755 2913.035 2235.925 ;
        RECT 2913.325 2235.755 2913.495 2235.925 ;
        RECT 2913.785 2235.755 2913.955 2235.925 ;
        RECT 5.665 2230.315 5.835 2230.485 ;
        RECT 6.125 2230.315 6.295 2230.485 ;
        RECT 6.585 2230.315 6.755 2230.485 ;
        RECT 2906.425 2230.315 2906.595 2230.485 ;
        RECT 2912.865 2230.315 2913.035 2230.485 ;
        RECT 2913.325 2230.315 2913.495 2230.485 ;
        RECT 2913.785 2230.315 2913.955 2230.485 ;
        RECT 5.665 2224.875 5.835 2225.045 ;
        RECT 6.125 2224.875 6.295 2225.045 ;
        RECT 6.585 2224.875 6.755 2225.045 ;
        RECT 2906.425 2224.875 2906.595 2225.045 ;
        RECT 2912.865 2224.875 2913.035 2225.045 ;
        RECT 2913.325 2224.875 2913.495 2225.045 ;
        RECT 2913.785 2224.875 2913.955 2225.045 ;
        RECT 5.665 2219.435 5.835 2219.605 ;
        RECT 6.125 2219.435 6.295 2219.605 ;
        RECT 6.585 2219.435 6.755 2219.605 ;
        RECT 2906.425 2219.435 2906.595 2219.605 ;
        RECT 2912.865 2219.435 2913.035 2219.605 ;
        RECT 2913.325 2219.435 2913.495 2219.605 ;
        RECT 2913.785 2219.435 2913.955 2219.605 ;
        RECT 5.665 2213.995 5.835 2214.165 ;
        RECT 6.125 2213.995 6.295 2214.165 ;
        RECT 6.585 2213.995 6.755 2214.165 ;
        RECT 2906.425 2213.995 2906.595 2214.165 ;
        RECT 2912.865 2213.995 2913.035 2214.165 ;
        RECT 2913.325 2213.995 2913.495 2214.165 ;
        RECT 2913.785 2213.995 2913.955 2214.165 ;
        RECT 5.665 2208.555 5.835 2208.725 ;
        RECT 6.125 2208.555 6.295 2208.725 ;
        RECT 6.585 2208.555 6.755 2208.725 ;
        RECT 2906.425 2208.555 2906.595 2208.725 ;
        RECT 2912.865 2208.555 2913.035 2208.725 ;
        RECT 2913.325 2208.555 2913.495 2208.725 ;
        RECT 2913.785 2208.555 2913.955 2208.725 ;
        RECT 5.665 2203.115 5.835 2203.285 ;
        RECT 6.125 2203.115 6.295 2203.285 ;
        RECT 6.585 2203.115 6.755 2203.285 ;
        RECT 2906.425 2203.115 2906.595 2203.285 ;
        RECT 2912.865 2203.115 2913.035 2203.285 ;
        RECT 2913.325 2203.115 2913.495 2203.285 ;
        RECT 2913.785 2203.115 2913.955 2203.285 ;
        RECT 5.665 2197.675 5.835 2197.845 ;
        RECT 6.125 2197.675 6.295 2197.845 ;
        RECT 6.585 2197.675 6.755 2197.845 ;
        RECT 2906.425 2197.675 2906.595 2197.845 ;
        RECT 2912.865 2197.675 2913.035 2197.845 ;
        RECT 2913.325 2197.675 2913.495 2197.845 ;
        RECT 2913.785 2197.675 2913.955 2197.845 ;
        RECT 5.665 2192.235 5.835 2192.405 ;
        RECT 6.125 2192.235 6.295 2192.405 ;
        RECT 6.585 2192.235 6.755 2192.405 ;
        RECT 2906.425 2192.235 2906.595 2192.405 ;
        RECT 2912.865 2192.235 2913.035 2192.405 ;
        RECT 2913.325 2192.235 2913.495 2192.405 ;
        RECT 2913.785 2192.235 2913.955 2192.405 ;
        RECT 5.665 2186.795 5.835 2186.965 ;
        RECT 6.125 2186.795 6.295 2186.965 ;
        RECT 6.585 2186.795 6.755 2186.965 ;
        RECT 2906.425 2186.795 2906.595 2186.965 ;
        RECT 2912.865 2186.795 2913.035 2186.965 ;
        RECT 2913.325 2186.795 2913.495 2186.965 ;
        RECT 2913.785 2186.795 2913.955 2186.965 ;
        RECT 5.665 2181.355 5.835 2181.525 ;
        RECT 6.125 2181.355 6.295 2181.525 ;
        RECT 6.585 2181.355 6.755 2181.525 ;
        RECT 2906.425 2181.355 2906.595 2181.525 ;
        RECT 2912.865 2181.355 2913.035 2181.525 ;
        RECT 2913.325 2181.355 2913.495 2181.525 ;
        RECT 2913.785 2181.355 2913.955 2181.525 ;
        RECT 5.665 2175.915 5.835 2176.085 ;
        RECT 6.125 2175.915 6.295 2176.085 ;
        RECT 6.585 2175.915 6.755 2176.085 ;
        RECT 2906.425 2175.915 2906.595 2176.085 ;
        RECT 2912.865 2175.915 2913.035 2176.085 ;
        RECT 2913.325 2175.915 2913.495 2176.085 ;
        RECT 2913.785 2175.915 2913.955 2176.085 ;
        RECT 5.665 2170.475 5.835 2170.645 ;
        RECT 6.125 2170.475 6.295 2170.645 ;
        RECT 6.585 2170.475 6.755 2170.645 ;
        RECT 2906.425 2170.475 2906.595 2170.645 ;
        RECT 2912.865 2170.475 2913.035 2170.645 ;
        RECT 2913.325 2170.475 2913.495 2170.645 ;
        RECT 2913.785 2170.475 2913.955 2170.645 ;
        RECT 5.665 2165.035 5.835 2165.205 ;
        RECT 6.125 2165.035 6.295 2165.205 ;
        RECT 6.585 2165.035 6.755 2165.205 ;
        RECT 2906.425 2165.035 2906.595 2165.205 ;
        RECT 2912.865 2165.035 2913.035 2165.205 ;
        RECT 2913.325 2165.035 2913.495 2165.205 ;
        RECT 2913.785 2165.035 2913.955 2165.205 ;
        RECT 5.665 2159.595 5.835 2159.765 ;
        RECT 6.125 2159.595 6.295 2159.765 ;
        RECT 6.585 2159.595 6.755 2159.765 ;
        RECT 2906.425 2159.595 2906.595 2159.765 ;
        RECT 2912.865 2159.595 2913.035 2159.765 ;
        RECT 2913.325 2159.595 2913.495 2159.765 ;
        RECT 2913.785 2159.595 2913.955 2159.765 ;
        RECT 5.665 2154.155 5.835 2154.325 ;
        RECT 6.125 2154.155 6.295 2154.325 ;
        RECT 6.585 2154.155 6.755 2154.325 ;
        RECT 2906.425 2154.155 2906.595 2154.325 ;
        RECT 2912.865 2154.155 2913.035 2154.325 ;
        RECT 2913.325 2154.155 2913.495 2154.325 ;
        RECT 2913.785 2154.155 2913.955 2154.325 ;
        RECT 5.665 2148.715 5.835 2148.885 ;
        RECT 6.125 2148.715 6.295 2148.885 ;
        RECT 6.585 2148.715 6.755 2148.885 ;
        RECT 2906.425 2148.715 2906.595 2148.885 ;
        RECT 2912.865 2148.715 2913.035 2148.885 ;
        RECT 2913.325 2148.715 2913.495 2148.885 ;
        RECT 2913.785 2148.715 2913.955 2148.885 ;
        RECT 5.665 2143.275 5.835 2143.445 ;
        RECT 6.125 2143.275 6.295 2143.445 ;
        RECT 6.585 2143.275 6.755 2143.445 ;
        RECT 2906.425 2143.275 2906.595 2143.445 ;
        RECT 2912.865 2143.275 2913.035 2143.445 ;
        RECT 2913.325 2143.275 2913.495 2143.445 ;
        RECT 2913.785 2143.275 2913.955 2143.445 ;
        RECT 5.665 2137.835 5.835 2138.005 ;
        RECT 6.125 2137.835 6.295 2138.005 ;
        RECT 6.585 2137.835 6.755 2138.005 ;
        RECT 2906.425 2137.835 2906.595 2138.005 ;
        RECT 2912.865 2137.835 2913.035 2138.005 ;
        RECT 2913.325 2137.835 2913.495 2138.005 ;
        RECT 2913.785 2137.835 2913.955 2138.005 ;
        RECT 5.665 2132.395 5.835 2132.565 ;
        RECT 6.125 2132.395 6.295 2132.565 ;
        RECT 6.585 2132.395 6.755 2132.565 ;
        RECT 2906.425 2132.395 2906.595 2132.565 ;
        RECT 2912.865 2132.395 2913.035 2132.565 ;
        RECT 2913.325 2132.395 2913.495 2132.565 ;
        RECT 2913.785 2132.395 2913.955 2132.565 ;
        RECT 5.665 2126.955 5.835 2127.125 ;
        RECT 6.125 2126.955 6.295 2127.125 ;
        RECT 6.585 2126.955 6.755 2127.125 ;
        RECT 2906.425 2126.955 2906.595 2127.125 ;
        RECT 2912.865 2126.955 2913.035 2127.125 ;
        RECT 2913.325 2126.955 2913.495 2127.125 ;
        RECT 2913.785 2126.955 2913.955 2127.125 ;
        RECT 5.665 2121.515 5.835 2121.685 ;
        RECT 6.125 2121.515 6.295 2121.685 ;
        RECT 6.585 2121.515 6.755 2121.685 ;
        RECT 2906.425 2121.515 2906.595 2121.685 ;
        RECT 2912.865 2121.515 2913.035 2121.685 ;
        RECT 2913.325 2121.515 2913.495 2121.685 ;
        RECT 2913.785 2121.515 2913.955 2121.685 ;
        RECT 5.665 2116.075 5.835 2116.245 ;
        RECT 6.125 2116.075 6.295 2116.245 ;
        RECT 6.585 2116.075 6.755 2116.245 ;
        RECT 2906.425 2116.075 2906.595 2116.245 ;
        RECT 2909.185 2116.075 2909.355 2116.245 ;
        RECT 2909.645 2116.075 2909.815 2116.245 ;
        RECT 2910.105 2116.075 2910.275 2116.245 ;
        RECT 2912.865 2116.075 2913.035 2116.245 ;
        RECT 2913.325 2116.075 2913.495 2116.245 ;
        RECT 2913.785 2116.075 2913.955 2116.245 ;
        RECT 5.665 2110.635 5.835 2110.805 ;
        RECT 6.125 2110.635 6.295 2110.805 ;
        RECT 6.585 2110.635 6.755 2110.805 ;
        RECT 2906.425 2110.635 2906.595 2110.805 ;
        RECT 2912.865 2110.635 2913.035 2110.805 ;
        RECT 2913.325 2110.635 2913.495 2110.805 ;
        RECT 2913.785 2110.635 2913.955 2110.805 ;
        RECT 5.665 2105.195 5.835 2105.365 ;
        RECT 6.125 2105.195 6.295 2105.365 ;
        RECT 6.585 2105.195 6.755 2105.365 ;
        RECT 2906.425 2105.195 2906.595 2105.365 ;
        RECT 2912.865 2105.195 2913.035 2105.365 ;
        RECT 2913.325 2105.195 2913.495 2105.365 ;
        RECT 2913.785 2105.195 2913.955 2105.365 ;
        RECT 5.665 2099.755 5.835 2099.925 ;
        RECT 6.125 2099.755 6.295 2099.925 ;
        RECT 6.585 2099.755 6.755 2099.925 ;
        RECT 2906.425 2099.755 2906.595 2099.925 ;
        RECT 2912.865 2099.755 2913.035 2099.925 ;
        RECT 2913.325 2099.755 2913.495 2099.925 ;
        RECT 2913.785 2099.755 2913.955 2099.925 ;
        RECT 5.665 2094.315 5.835 2094.485 ;
        RECT 6.125 2094.315 6.295 2094.485 ;
        RECT 6.585 2094.315 6.755 2094.485 ;
        RECT 2906.425 2094.315 2906.595 2094.485 ;
        RECT 2912.865 2094.315 2913.035 2094.485 ;
        RECT 2913.325 2094.315 2913.495 2094.485 ;
        RECT 2913.785 2094.315 2913.955 2094.485 ;
        RECT 5.665 2088.875 5.835 2089.045 ;
        RECT 6.125 2088.875 6.295 2089.045 ;
        RECT 6.585 2088.875 6.755 2089.045 ;
        RECT 2906.425 2088.875 2906.595 2089.045 ;
        RECT 2912.865 2088.875 2913.035 2089.045 ;
        RECT 2913.325 2088.875 2913.495 2089.045 ;
        RECT 2913.785 2088.875 2913.955 2089.045 ;
        RECT 5.665 2083.435 5.835 2083.605 ;
        RECT 6.125 2083.435 6.295 2083.605 ;
        RECT 6.585 2083.435 6.755 2083.605 ;
        RECT 2906.425 2083.435 2906.595 2083.605 ;
        RECT 2912.865 2083.435 2913.035 2083.605 ;
        RECT 2913.325 2083.435 2913.495 2083.605 ;
        RECT 2913.785 2083.435 2913.955 2083.605 ;
        RECT 5.665 2077.995 5.835 2078.165 ;
        RECT 6.125 2077.995 6.295 2078.165 ;
        RECT 6.585 2077.995 6.755 2078.165 ;
        RECT 2906.425 2077.995 2906.595 2078.165 ;
        RECT 2912.865 2077.995 2913.035 2078.165 ;
        RECT 2913.325 2077.995 2913.495 2078.165 ;
        RECT 2913.785 2077.995 2913.955 2078.165 ;
        RECT 5.665 2072.555 5.835 2072.725 ;
        RECT 6.125 2072.555 6.295 2072.725 ;
        RECT 6.585 2072.555 6.755 2072.725 ;
        RECT 2906.425 2072.555 2906.595 2072.725 ;
        RECT 2912.865 2072.555 2913.035 2072.725 ;
        RECT 2913.325 2072.555 2913.495 2072.725 ;
        RECT 2913.785 2072.555 2913.955 2072.725 ;
        RECT 5.665 2067.115 5.835 2067.285 ;
        RECT 6.125 2067.115 6.295 2067.285 ;
        RECT 6.585 2067.115 6.755 2067.285 ;
        RECT 2906.425 2067.115 2906.595 2067.285 ;
        RECT 2912.865 2067.115 2913.035 2067.285 ;
        RECT 2913.325 2067.115 2913.495 2067.285 ;
        RECT 2913.785 2067.115 2913.955 2067.285 ;
        RECT 5.665 2061.675 5.835 2061.845 ;
        RECT 6.125 2061.675 6.295 2061.845 ;
        RECT 6.585 2061.675 6.755 2061.845 ;
        RECT 2906.425 2061.675 2906.595 2061.845 ;
        RECT 2912.865 2061.675 2913.035 2061.845 ;
        RECT 2913.325 2061.675 2913.495 2061.845 ;
        RECT 2913.785 2061.675 2913.955 2061.845 ;
        RECT 5.665 2056.235 5.835 2056.405 ;
        RECT 6.125 2056.235 6.295 2056.405 ;
        RECT 6.585 2056.235 6.755 2056.405 ;
        RECT 2906.425 2056.235 2906.595 2056.405 ;
        RECT 2912.865 2056.235 2913.035 2056.405 ;
        RECT 2913.325 2056.235 2913.495 2056.405 ;
        RECT 2913.785 2056.235 2913.955 2056.405 ;
        RECT 5.665 2050.795 5.835 2050.965 ;
        RECT 6.125 2050.795 6.295 2050.965 ;
        RECT 6.585 2050.795 6.755 2050.965 ;
        RECT 2906.425 2050.795 2906.595 2050.965 ;
        RECT 2912.865 2050.795 2913.035 2050.965 ;
        RECT 2913.325 2050.795 2913.495 2050.965 ;
        RECT 2913.785 2050.795 2913.955 2050.965 ;
        RECT 5.665 2045.355 5.835 2045.525 ;
        RECT 6.125 2045.355 6.295 2045.525 ;
        RECT 6.585 2045.355 6.755 2045.525 ;
        RECT 2906.425 2045.355 2906.595 2045.525 ;
        RECT 2912.865 2045.355 2913.035 2045.525 ;
        RECT 2913.325 2045.355 2913.495 2045.525 ;
        RECT 2913.785 2045.355 2913.955 2045.525 ;
        RECT 5.665 2039.915 5.835 2040.085 ;
        RECT 6.125 2039.915 6.295 2040.085 ;
        RECT 6.585 2039.915 6.755 2040.085 ;
        RECT 2906.425 2039.915 2906.595 2040.085 ;
        RECT 2912.865 2039.915 2913.035 2040.085 ;
        RECT 2913.325 2039.915 2913.495 2040.085 ;
        RECT 2913.785 2039.915 2913.955 2040.085 ;
        RECT 5.665 2034.475 5.835 2034.645 ;
        RECT 6.125 2034.475 6.295 2034.645 ;
        RECT 6.585 2034.475 6.755 2034.645 ;
        RECT 2906.425 2034.475 2906.595 2034.645 ;
        RECT 2912.865 2034.475 2913.035 2034.645 ;
        RECT 2913.325 2034.475 2913.495 2034.645 ;
        RECT 2913.785 2034.475 2913.955 2034.645 ;
        RECT 5.665 2029.035 5.835 2029.205 ;
        RECT 6.125 2029.035 6.295 2029.205 ;
        RECT 6.585 2029.035 6.755 2029.205 ;
        RECT 2906.425 2029.035 2906.595 2029.205 ;
        RECT 2912.865 2029.035 2913.035 2029.205 ;
        RECT 2913.325 2029.035 2913.495 2029.205 ;
        RECT 2913.785 2029.035 2913.955 2029.205 ;
        RECT 5.665 2023.595 5.835 2023.765 ;
        RECT 6.125 2023.595 6.295 2023.765 ;
        RECT 6.585 2023.595 6.755 2023.765 ;
        RECT 2906.425 2023.595 2906.595 2023.765 ;
        RECT 2912.865 2023.595 2913.035 2023.765 ;
        RECT 2913.325 2023.595 2913.495 2023.765 ;
        RECT 2913.785 2023.595 2913.955 2023.765 ;
        RECT 5.665 2018.155 5.835 2018.325 ;
        RECT 6.125 2018.155 6.295 2018.325 ;
        RECT 6.585 2018.155 6.755 2018.325 ;
        RECT 2906.425 2018.155 2906.595 2018.325 ;
        RECT 2912.865 2018.155 2913.035 2018.325 ;
        RECT 2913.325 2018.155 2913.495 2018.325 ;
        RECT 2913.785 2018.155 2913.955 2018.325 ;
        RECT 5.665 2012.715 5.835 2012.885 ;
        RECT 6.125 2012.715 6.295 2012.885 ;
        RECT 6.585 2012.715 6.755 2012.885 ;
        RECT 2906.425 2012.715 2906.595 2012.885 ;
        RECT 2912.865 2012.715 2913.035 2012.885 ;
        RECT 2913.325 2012.715 2913.495 2012.885 ;
        RECT 2913.785 2012.715 2913.955 2012.885 ;
        RECT 5.665 2007.275 5.835 2007.445 ;
        RECT 6.125 2007.275 6.295 2007.445 ;
        RECT 6.585 2007.275 6.755 2007.445 ;
        RECT 2906.425 2007.275 2906.595 2007.445 ;
        RECT 2912.865 2007.275 2913.035 2007.445 ;
        RECT 2913.325 2007.275 2913.495 2007.445 ;
        RECT 2913.785 2007.275 2913.955 2007.445 ;
        RECT 5.665 2001.835 5.835 2002.005 ;
        RECT 6.125 2001.835 6.295 2002.005 ;
        RECT 6.585 2001.835 6.755 2002.005 ;
        RECT 2906.425 2001.835 2906.595 2002.005 ;
        RECT 2912.865 2001.835 2913.035 2002.005 ;
        RECT 2913.325 2001.835 2913.495 2002.005 ;
        RECT 2913.785 2001.835 2913.955 2002.005 ;
        RECT 5.665 1996.395 5.835 1996.565 ;
        RECT 6.125 1996.395 6.295 1996.565 ;
        RECT 6.585 1996.395 6.755 1996.565 ;
        RECT 2906.425 1996.395 2906.595 1996.565 ;
        RECT 2912.865 1996.395 2913.035 1996.565 ;
        RECT 2913.325 1996.395 2913.495 1996.565 ;
        RECT 2913.785 1996.395 2913.955 1996.565 ;
        RECT 5.665 1990.955 5.835 1991.125 ;
        RECT 6.125 1990.955 6.295 1991.125 ;
        RECT 6.585 1990.955 6.755 1991.125 ;
        RECT 2906.425 1990.955 2906.595 1991.125 ;
        RECT 2912.865 1990.955 2913.035 1991.125 ;
        RECT 2913.325 1990.955 2913.495 1991.125 ;
        RECT 2913.785 1990.955 2913.955 1991.125 ;
        RECT 5.665 1985.515 5.835 1985.685 ;
        RECT 6.125 1985.515 6.295 1985.685 ;
        RECT 6.585 1985.515 6.755 1985.685 ;
        RECT 8.885 1985.515 9.055 1985.685 ;
        RECT 9.345 1985.515 9.515 1985.685 ;
        RECT 9.805 1985.515 9.975 1985.685 ;
        RECT 2906.425 1985.515 2906.595 1985.685 ;
        RECT 2912.865 1985.515 2913.035 1985.685 ;
        RECT 2913.325 1985.515 2913.495 1985.685 ;
        RECT 2913.785 1985.515 2913.955 1985.685 ;
        RECT 5.665 1980.075 5.835 1980.245 ;
        RECT 6.125 1980.075 6.295 1980.245 ;
        RECT 6.585 1980.075 6.755 1980.245 ;
        RECT 2906.425 1980.075 2906.595 1980.245 ;
        RECT 2912.865 1980.075 2913.035 1980.245 ;
        RECT 2913.325 1980.075 2913.495 1980.245 ;
        RECT 2913.785 1980.075 2913.955 1980.245 ;
        RECT 5.665 1974.635 5.835 1974.805 ;
        RECT 6.125 1974.635 6.295 1974.805 ;
        RECT 6.585 1974.635 6.755 1974.805 ;
        RECT 2906.425 1974.635 2906.595 1974.805 ;
        RECT 2912.865 1974.635 2913.035 1974.805 ;
        RECT 2913.325 1974.635 2913.495 1974.805 ;
        RECT 2913.785 1974.635 2913.955 1974.805 ;
        RECT 5.665 1969.195 5.835 1969.365 ;
        RECT 6.125 1969.195 6.295 1969.365 ;
        RECT 6.585 1969.195 6.755 1969.365 ;
        RECT 2906.425 1969.195 2906.595 1969.365 ;
        RECT 2912.865 1969.195 2913.035 1969.365 ;
        RECT 2913.325 1969.195 2913.495 1969.365 ;
        RECT 2913.785 1969.195 2913.955 1969.365 ;
        RECT 5.665 1963.755 5.835 1963.925 ;
        RECT 6.125 1963.755 6.295 1963.925 ;
        RECT 6.585 1963.755 6.755 1963.925 ;
        RECT 2906.425 1963.755 2906.595 1963.925 ;
        RECT 2912.865 1963.755 2913.035 1963.925 ;
        RECT 2913.325 1963.755 2913.495 1963.925 ;
        RECT 2913.785 1963.755 2913.955 1963.925 ;
        RECT 5.665 1958.315 5.835 1958.485 ;
        RECT 6.125 1958.315 6.295 1958.485 ;
        RECT 6.585 1958.315 6.755 1958.485 ;
        RECT 2906.425 1958.315 2906.595 1958.485 ;
        RECT 2912.865 1958.315 2913.035 1958.485 ;
        RECT 2913.325 1958.315 2913.495 1958.485 ;
        RECT 2913.785 1958.315 2913.955 1958.485 ;
        RECT 5.665 1952.875 5.835 1953.045 ;
        RECT 6.125 1952.875 6.295 1953.045 ;
        RECT 6.585 1952.875 6.755 1953.045 ;
        RECT 8.885 1952.875 9.055 1953.045 ;
        RECT 9.345 1952.875 9.515 1953.045 ;
        RECT 9.805 1952.875 9.975 1953.045 ;
        RECT 2906.425 1952.875 2906.595 1953.045 ;
        RECT 2912.865 1952.875 2913.035 1953.045 ;
        RECT 2913.325 1952.875 2913.495 1953.045 ;
        RECT 2913.785 1952.875 2913.955 1953.045 ;
        RECT 5.665 1947.435 5.835 1947.605 ;
        RECT 6.125 1947.435 6.295 1947.605 ;
        RECT 6.585 1947.435 6.755 1947.605 ;
        RECT 2906.425 1947.435 2906.595 1947.605 ;
        RECT 2912.865 1947.435 2913.035 1947.605 ;
        RECT 2913.325 1947.435 2913.495 1947.605 ;
        RECT 2913.785 1947.435 2913.955 1947.605 ;
        RECT 5.665 1941.995 5.835 1942.165 ;
        RECT 6.125 1941.995 6.295 1942.165 ;
        RECT 6.585 1941.995 6.755 1942.165 ;
        RECT 2906.425 1941.995 2906.595 1942.165 ;
        RECT 2912.865 1941.995 2913.035 1942.165 ;
        RECT 2913.325 1941.995 2913.495 1942.165 ;
        RECT 2913.785 1941.995 2913.955 1942.165 ;
        RECT 5.665 1936.555 5.835 1936.725 ;
        RECT 6.125 1936.555 6.295 1936.725 ;
        RECT 6.585 1936.555 6.755 1936.725 ;
        RECT 2906.425 1936.555 2906.595 1936.725 ;
        RECT 2909.185 1936.555 2909.355 1936.725 ;
        RECT 2909.645 1936.555 2909.815 1936.725 ;
        RECT 2910.105 1936.555 2910.275 1936.725 ;
        RECT 2912.865 1936.555 2913.035 1936.725 ;
        RECT 2913.325 1936.555 2913.495 1936.725 ;
        RECT 2913.785 1936.555 2913.955 1936.725 ;
        RECT 5.665 1931.115 5.835 1931.285 ;
        RECT 6.125 1931.115 6.295 1931.285 ;
        RECT 6.585 1931.115 6.755 1931.285 ;
        RECT 2906.425 1931.115 2906.595 1931.285 ;
        RECT 2912.865 1931.115 2913.035 1931.285 ;
        RECT 2913.325 1931.115 2913.495 1931.285 ;
        RECT 2913.785 1931.115 2913.955 1931.285 ;
        RECT 5.665 1925.675 5.835 1925.845 ;
        RECT 6.125 1925.675 6.295 1925.845 ;
        RECT 6.585 1925.675 6.755 1925.845 ;
        RECT 2906.425 1925.675 2906.595 1925.845 ;
        RECT 2912.865 1925.675 2913.035 1925.845 ;
        RECT 2913.325 1925.675 2913.495 1925.845 ;
        RECT 2913.785 1925.675 2913.955 1925.845 ;
        RECT 5.665 1920.235 5.835 1920.405 ;
        RECT 6.125 1920.235 6.295 1920.405 ;
        RECT 6.585 1920.235 6.755 1920.405 ;
        RECT 2906.425 1920.235 2906.595 1920.405 ;
        RECT 2912.865 1920.235 2913.035 1920.405 ;
        RECT 2913.325 1920.235 2913.495 1920.405 ;
        RECT 2913.785 1920.235 2913.955 1920.405 ;
        RECT 5.665 1914.795 5.835 1914.965 ;
        RECT 6.125 1914.795 6.295 1914.965 ;
        RECT 6.585 1914.795 6.755 1914.965 ;
        RECT 2906.425 1914.795 2906.595 1914.965 ;
        RECT 2912.865 1914.795 2913.035 1914.965 ;
        RECT 2913.325 1914.795 2913.495 1914.965 ;
        RECT 2913.785 1914.795 2913.955 1914.965 ;
        RECT 5.665 1909.355 5.835 1909.525 ;
        RECT 6.125 1909.355 6.295 1909.525 ;
        RECT 6.585 1909.355 6.755 1909.525 ;
        RECT 2906.425 1909.355 2906.595 1909.525 ;
        RECT 2912.865 1909.355 2913.035 1909.525 ;
        RECT 2913.325 1909.355 2913.495 1909.525 ;
        RECT 2913.785 1909.355 2913.955 1909.525 ;
        RECT 5.665 1903.915 5.835 1904.085 ;
        RECT 6.125 1903.915 6.295 1904.085 ;
        RECT 6.585 1903.915 6.755 1904.085 ;
        RECT 2906.425 1903.915 2906.595 1904.085 ;
        RECT 2912.865 1903.915 2913.035 1904.085 ;
        RECT 2913.325 1903.915 2913.495 1904.085 ;
        RECT 2913.785 1903.915 2913.955 1904.085 ;
        RECT 5.665 1898.475 5.835 1898.645 ;
        RECT 6.125 1898.475 6.295 1898.645 ;
        RECT 6.585 1898.475 6.755 1898.645 ;
        RECT 2906.425 1898.475 2906.595 1898.645 ;
        RECT 2912.865 1898.475 2913.035 1898.645 ;
        RECT 2913.325 1898.475 2913.495 1898.645 ;
        RECT 2913.785 1898.475 2913.955 1898.645 ;
        RECT 5.665 1893.035 5.835 1893.205 ;
        RECT 6.125 1893.035 6.295 1893.205 ;
        RECT 6.585 1893.035 6.755 1893.205 ;
        RECT 2906.425 1893.035 2906.595 1893.205 ;
        RECT 2912.865 1893.035 2913.035 1893.205 ;
        RECT 2913.325 1893.035 2913.495 1893.205 ;
        RECT 2913.785 1893.035 2913.955 1893.205 ;
        RECT 5.665 1887.595 5.835 1887.765 ;
        RECT 6.125 1887.595 6.295 1887.765 ;
        RECT 6.585 1887.595 6.755 1887.765 ;
        RECT 2906.425 1887.595 2906.595 1887.765 ;
        RECT 2912.865 1887.595 2913.035 1887.765 ;
        RECT 2913.325 1887.595 2913.495 1887.765 ;
        RECT 2913.785 1887.595 2913.955 1887.765 ;
        RECT 5.665 1882.155 5.835 1882.325 ;
        RECT 6.125 1882.155 6.295 1882.325 ;
        RECT 6.585 1882.155 6.755 1882.325 ;
        RECT 2906.425 1882.155 2906.595 1882.325 ;
        RECT 2912.865 1882.155 2913.035 1882.325 ;
        RECT 2913.325 1882.155 2913.495 1882.325 ;
        RECT 2913.785 1882.155 2913.955 1882.325 ;
        RECT 5.665 1876.715 5.835 1876.885 ;
        RECT 6.125 1876.715 6.295 1876.885 ;
        RECT 6.585 1876.715 6.755 1876.885 ;
        RECT 2906.425 1876.715 2906.595 1876.885 ;
        RECT 2912.865 1876.715 2913.035 1876.885 ;
        RECT 2913.325 1876.715 2913.495 1876.885 ;
        RECT 2913.785 1876.715 2913.955 1876.885 ;
        RECT 5.665 1871.275 5.835 1871.445 ;
        RECT 6.125 1871.275 6.295 1871.445 ;
        RECT 6.585 1871.275 6.755 1871.445 ;
        RECT 2906.425 1871.275 2906.595 1871.445 ;
        RECT 2912.865 1871.275 2913.035 1871.445 ;
        RECT 2913.325 1871.275 2913.495 1871.445 ;
        RECT 2913.785 1871.275 2913.955 1871.445 ;
        RECT 5.665 1865.835 5.835 1866.005 ;
        RECT 6.125 1865.835 6.295 1866.005 ;
        RECT 6.585 1865.835 6.755 1866.005 ;
        RECT 2906.425 1865.835 2906.595 1866.005 ;
        RECT 2912.865 1865.835 2913.035 1866.005 ;
        RECT 2913.325 1865.835 2913.495 1866.005 ;
        RECT 2913.785 1865.835 2913.955 1866.005 ;
        RECT 5.665 1860.395 5.835 1860.565 ;
        RECT 6.125 1860.395 6.295 1860.565 ;
        RECT 6.585 1860.395 6.755 1860.565 ;
        RECT 2906.425 1860.395 2906.595 1860.565 ;
        RECT 2912.865 1860.395 2913.035 1860.565 ;
        RECT 2913.325 1860.395 2913.495 1860.565 ;
        RECT 2913.785 1860.395 2913.955 1860.565 ;
        RECT 5.665 1854.955 5.835 1855.125 ;
        RECT 6.125 1854.955 6.295 1855.125 ;
        RECT 6.585 1854.955 6.755 1855.125 ;
        RECT 2906.425 1854.955 2906.595 1855.125 ;
        RECT 2912.865 1854.955 2913.035 1855.125 ;
        RECT 2913.325 1854.955 2913.495 1855.125 ;
        RECT 2913.785 1854.955 2913.955 1855.125 ;
        RECT 5.665 1849.515 5.835 1849.685 ;
        RECT 6.125 1849.515 6.295 1849.685 ;
        RECT 6.585 1849.515 6.755 1849.685 ;
        RECT 2906.425 1849.515 2906.595 1849.685 ;
        RECT 2912.865 1849.515 2913.035 1849.685 ;
        RECT 2913.325 1849.515 2913.495 1849.685 ;
        RECT 2913.785 1849.515 2913.955 1849.685 ;
        RECT 5.665 1844.075 5.835 1844.245 ;
        RECT 6.125 1844.075 6.295 1844.245 ;
        RECT 6.585 1844.075 6.755 1844.245 ;
        RECT 2906.425 1844.075 2906.595 1844.245 ;
        RECT 2912.865 1844.075 2913.035 1844.245 ;
        RECT 2913.325 1844.075 2913.495 1844.245 ;
        RECT 2913.785 1844.075 2913.955 1844.245 ;
        RECT 5.665 1838.635 5.835 1838.805 ;
        RECT 6.125 1838.635 6.295 1838.805 ;
        RECT 6.585 1838.635 6.755 1838.805 ;
        RECT 2906.425 1838.635 2906.595 1838.805 ;
        RECT 2912.865 1838.635 2913.035 1838.805 ;
        RECT 2913.325 1838.635 2913.495 1838.805 ;
        RECT 2913.785 1838.635 2913.955 1838.805 ;
        RECT 5.665 1833.195 5.835 1833.365 ;
        RECT 6.125 1833.195 6.295 1833.365 ;
        RECT 6.585 1833.195 6.755 1833.365 ;
        RECT 2906.425 1833.195 2906.595 1833.365 ;
        RECT 2912.865 1833.195 2913.035 1833.365 ;
        RECT 2913.325 1833.195 2913.495 1833.365 ;
        RECT 2913.785 1833.195 2913.955 1833.365 ;
        RECT 5.665 1827.755 5.835 1827.925 ;
        RECT 6.125 1827.755 6.295 1827.925 ;
        RECT 6.585 1827.755 6.755 1827.925 ;
        RECT 2906.425 1827.755 2906.595 1827.925 ;
        RECT 2912.865 1827.755 2913.035 1827.925 ;
        RECT 2913.325 1827.755 2913.495 1827.925 ;
        RECT 2913.785 1827.755 2913.955 1827.925 ;
        RECT 5.665 1822.315 5.835 1822.485 ;
        RECT 6.125 1822.315 6.295 1822.485 ;
        RECT 6.585 1822.315 6.755 1822.485 ;
        RECT 2906.425 1822.315 2906.595 1822.485 ;
        RECT 2912.865 1822.315 2913.035 1822.485 ;
        RECT 2913.325 1822.315 2913.495 1822.485 ;
        RECT 2913.785 1822.315 2913.955 1822.485 ;
        RECT 5.665 1816.875 5.835 1817.045 ;
        RECT 6.125 1816.875 6.295 1817.045 ;
        RECT 6.585 1816.875 6.755 1817.045 ;
        RECT 2906.425 1816.875 2906.595 1817.045 ;
        RECT 2912.865 1816.875 2913.035 1817.045 ;
        RECT 2913.325 1816.875 2913.495 1817.045 ;
        RECT 2913.785 1816.875 2913.955 1817.045 ;
        RECT 5.665 1811.435 5.835 1811.605 ;
        RECT 6.125 1811.435 6.295 1811.605 ;
        RECT 6.585 1811.435 6.755 1811.605 ;
        RECT 2906.425 1811.435 2906.595 1811.605 ;
        RECT 2912.865 1811.435 2913.035 1811.605 ;
        RECT 2913.325 1811.435 2913.495 1811.605 ;
        RECT 2913.785 1811.435 2913.955 1811.605 ;
        RECT 5.665 1805.995 5.835 1806.165 ;
        RECT 6.125 1805.995 6.295 1806.165 ;
        RECT 6.585 1805.995 6.755 1806.165 ;
        RECT 2906.425 1805.995 2906.595 1806.165 ;
        RECT 2912.865 1805.995 2913.035 1806.165 ;
        RECT 2913.325 1805.995 2913.495 1806.165 ;
        RECT 2913.785 1805.995 2913.955 1806.165 ;
        RECT 5.665 1800.555 5.835 1800.725 ;
        RECT 6.125 1800.555 6.295 1800.725 ;
        RECT 6.585 1800.555 6.755 1800.725 ;
        RECT 2906.425 1800.555 2906.595 1800.725 ;
        RECT 2912.865 1800.555 2913.035 1800.725 ;
        RECT 2913.325 1800.555 2913.495 1800.725 ;
        RECT 2913.785 1800.555 2913.955 1800.725 ;
        RECT 5.665 1795.115 5.835 1795.285 ;
        RECT 6.125 1795.115 6.295 1795.285 ;
        RECT 6.585 1795.115 6.755 1795.285 ;
        RECT 2906.425 1795.115 2906.595 1795.285 ;
        RECT 2912.865 1795.115 2913.035 1795.285 ;
        RECT 2913.325 1795.115 2913.495 1795.285 ;
        RECT 2913.785 1795.115 2913.955 1795.285 ;
        RECT 5.665 1789.675 5.835 1789.845 ;
        RECT 6.125 1789.675 6.295 1789.845 ;
        RECT 6.585 1789.675 6.755 1789.845 ;
        RECT 2906.425 1789.675 2906.595 1789.845 ;
        RECT 2912.865 1789.675 2913.035 1789.845 ;
        RECT 2913.325 1789.675 2913.495 1789.845 ;
        RECT 2913.785 1789.675 2913.955 1789.845 ;
        RECT 5.665 1784.235 5.835 1784.405 ;
        RECT 6.125 1784.235 6.295 1784.405 ;
        RECT 6.585 1784.235 6.755 1784.405 ;
        RECT 2906.425 1784.235 2906.595 1784.405 ;
        RECT 2912.865 1784.235 2913.035 1784.405 ;
        RECT 2913.325 1784.235 2913.495 1784.405 ;
        RECT 2913.785 1784.235 2913.955 1784.405 ;
        RECT 5.665 1778.795 5.835 1778.965 ;
        RECT 6.125 1778.795 6.295 1778.965 ;
        RECT 6.585 1778.795 6.755 1778.965 ;
        RECT 8.885 1778.795 9.055 1778.965 ;
        RECT 9.345 1778.795 9.515 1778.965 ;
        RECT 9.805 1778.795 9.975 1778.965 ;
        RECT 2906.425 1778.795 2906.595 1778.965 ;
        RECT 2912.865 1778.795 2913.035 1778.965 ;
        RECT 2913.325 1778.795 2913.495 1778.965 ;
        RECT 2913.785 1778.795 2913.955 1778.965 ;
        RECT 5.665 1773.355 5.835 1773.525 ;
        RECT 6.125 1773.355 6.295 1773.525 ;
        RECT 6.585 1773.355 6.755 1773.525 ;
        RECT 2906.425 1773.355 2906.595 1773.525 ;
        RECT 2912.865 1773.355 2913.035 1773.525 ;
        RECT 2913.325 1773.355 2913.495 1773.525 ;
        RECT 2913.785 1773.355 2913.955 1773.525 ;
        RECT 5.665 1767.915 5.835 1768.085 ;
        RECT 6.125 1767.915 6.295 1768.085 ;
        RECT 6.585 1767.915 6.755 1768.085 ;
        RECT 2906.425 1767.915 2906.595 1768.085 ;
        RECT 2912.865 1767.915 2913.035 1768.085 ;
        RECT 2913.325 1767.915 2913.495 1768.085 ;
        RECT 2913.785 1767.915 2913.955 1768.085 ;
        RECT 5.665 1762.475 5.835 1762.645 ;
        RECT 6.125 1762.475 6.295 1762.645 ;
        RECT 6.585 1762.475 6.755 1762.645 ;
        RECT 2906.425 1762.475 2906.595 1762.645 ;
        RECT 2912.865 1762.475 2913.035 1762.645 ;
        RECT 2913.325 1762.475 2913.495 1762.645 ;
        RECT 2913.785 1762.475 2913.955 1762.645 ;
        RECT 5.665 1757.035 5.835 1757.205 ;
        RECT 6.125 1757.035 6.295 1757.205 ;
        RECT 6.585 1757.035 6.755 1757.205 ;
        RECT 2906.425 1757.035 2906.595 1757.205 ;
        RECT 2912.865 1757.035 2913.035 1757.205 ;
        RECT 2913.325 1757.035 2913.495 1757.205 ;
        RECT 2913.785 1757.035 2913.955 1757.205 ;
        RECT 5.665 1751.595 5.835 1751.765 ;
        RECT 6.125 1751.595 6.295 1751.765 ;
        RECT 6.585 1751.595 6.755 1751.765 ;
        RECT 2906.425 1751.595 2906.595 1751.765 ;
        RECT 2912.865 1751.595 2913.035 1751.765 ;
        RECT 2913.325 1751.595 2913.495 1751.765 ;
        RECT 2913.785 1751.595 2913.955 1751.765 ;
        RECT 5.665 1746.155 5.835 1746.325 ;
        RECT 6.125 1746.155 6.295 1746.325 ;
        RECT 6.585 1746.155 6.755 1746.325 ;
        RECT 2906.425 1746.155 2906.595 1746.325 ;
        RECT 2912.865 1746.155 2913.035 1746.325 ;
        RECT 2913.325 1746.155 2913.495 1746.325 ;
        RECT 2913.785 1746.155 2913.955 1746.325 ;
        RECT 5.665 1740.715 5.835 1740.885 ;
        RECT 6.125 1740.715 6.295 1740.885 ;
        RECT 6.585 1740.715 6.755 1740.885 ;
        RECT 2906.425 1740.715 2906.595 1740.885 ;
        RECT 2912.865 1740.715 2913.035 1740.885 ;
        RECT 2913.325 1740.715 2913.495 1740.885 ;
        RECT 2913.785 1740.715 2913.955 1740.885 ;
        RECT 5.665 1735.275 5.835 1735.445 ;
        RECT 6.125 1735.275 6.295 1735.445 ;
        RECT 6.585 1735.275 6.755 1735.445 ;
        RECT 2906.425 1735.275 2906.595 1735.445 ;
        RECT 2912.865 1735.275 2913.035 1735.445 ;
        RECT 2913.325 1735.275 2913.495 1735.445 ;
        RECT 2913.785 1735.275 2913.955 1735.445 ;
        RECT 5.665 1729.835 5.835 1730.005 ;
        RECT 6.125 1729.835 6.295 1730.005 ;
        RECT 6.585 1729.835 6.755 1730.005 ;
        RECT 2906.425 1729.835 2906.595 1730.005 ;
        RECT 2912.865 1729.835 2913.035 1730.005 ;
        RECT 2913.325 1729.835 2913.495 1730.005 ;
        RECT 2913.785 1729.835 2913.955 1730.005 ;
        RECT 5.665 1724.395 5.835 1724.565 ;
        RECT 6.125 1724.395 6.295 1724.565 ;
        RECT 6.585 1724.395 6.755 1724.565 ;
        RECT 2906.425 1724.395 2906.595 1724.565 ;
        RECT 2912.865 1724.395 2913.035 1724.565 ;
        RECT 2913.325 1724.395 2913.495 1724.565 ;
        RECT 2913.785 1724.395 2913.955 1724.565 ;
        RECT 5.665 1718.955 5.835 1719.125 ;
        RECT 6.125 1718.955 6.295 1719.125 ;
        RECT 6.585 1718.955 6.755 1719.125 ;
        RECT 2906.425 1718.955 2906.595 1719.125 ;
        RECT 2912.865 1718.955 2913.035 1719.125 ;
        RECT 2913.325 1718.955 2913.495 1719.125 ;
        RECT 2913.785 1718.955 2913.955 1719.125 ;
        RECT 5.665 1713.515 5.835 1713.685 ;
        RECT 6.125 1713.515 6.295 1713.685 ;
        RECT 6.585 1713.515 6.755 1713.685 ;
        RECT 2906.425 1713.515 2906.595 1713.685 ;
        RECT 2912.865 1713.515 2913.035 1713.685 ;
        RECT 2913.325 1713.515 2913.495 1713.685 ;
        RECT 2913.785 1713.515 2913.955 1713.685 ;
        RECT 5.665 1708.075 5.835 1708.245 ;
        RECT 6.125 1708.075 6.295 1708.245 ;
        RECT 6.585 1708.075 6.755 1708.245 ;
        RECT 8.885 1708.075 9.055 1708.245 ;
        RECT 9.345 1708.075 9.515 1708.245 ;
        RECT 9.805 1708.075 9.975 1708.245 ;
        RECT 2906.425 1708.075 2906.595 1708.245 ;
        RECT 2912.865 1708.075 2913.035 1708.245 ;
        RECT 2913.325 1708.075 2913.495 1708.245 ;
        RECT 2913.785 1708.075 2913.955 1708.245 ;
        RECT 5.665 1702.635 5.835 1702.805 ;
        RECT 6.125 1702.635 6.295 1702.805 ;
        RECT 6.585 1702.635 6.755 1702.805 ;
        RECT 2906.425 1702.635 2906.595 1702.805 ;
        RECT 2912.865 1702.635 2913.035 1702.805 ;
        RECT 2913.325 1702.635 2913.495 1702.805 ;
        RECT 2913.785 1702.635 2913.955 1702.805 ;
        RECT 5.665 1697.195 5.835 1697.365 ;
        RECT 6.125 1697.195 6.295 1697.365 ;
        RECT 6.585 1697.195 6.755 1697.365 ;
        RECT 2906.425 1697.195 2906.595 1697.365 ;
        RECT 2912.865 1697.195 2913.035 1697.365 ;
        RECT 2913.325 1697.195 2913.495 1697.365 ;
        RECT 2913.785 1697.195 2913.955 1697.365 ;
        RECT 5.665 1691.755 5.835 1691.925 ;
        RECT 6.125 1691.755 6.295 1691.925 ;
        RECT 6.585 1691.755 6.755 1691.925 ;
        RECT 2906.425 1691.755 2906.595 1691.925 ;
        RECT 2912.865 1691.755 2913.035 1691.925 ;
        RECT 2913.325 1691.755 2913.495 1691.925 ;
        RECT 2913.785 1691.755 2913.955 1691.925 ;
        RECT 5.665 1686.315 5.835 1686.485 ;
        RECT 6.125 1686.315 6.295 1686.485 ;
        RECT 6.585 1686.315 6.755 1686.485 ;
        RECT 2906.425 1686.315 2906.595 1686.485 ;
        RECT 2912.865 1686.315 2913.035 1686.485 ;
        RECT 2913.325 1686.315 2913.495 1686.485 ;
        RECT 2913.785 1686.315 2913.955 1686.485 ;
        RECT 5.665 1680.875 5.835 1681.045 ;
        RECT 6.125 1680.875 6.295 1681.045 ;
        RECT 6.585 1680.875 6.755 1681.045 ;
        RECT 2906.425 1680.875 2906.595 1681.045 ;
        RECT 2912.865 1680.875 2913.035 1681.045 ;
        RECT 2913.325 1680.875 2913.495 1681.045 ;
        RECT 2913.785 1680.875 2913.955 1681.045 ;
        RECT 5.665 1675.435 5.835 1675.605 ;
        RECT 6.125 1675.435 6.295 1675.605 ;
        RECT 6.585 1675.435 6.755 1675.605 ;
        RECT 2906.425 1675.435 2906.595 1675.605 ;
        RECT 2912.865 1675.435 2913.035 1675.605 ;
        RECT 2913.325 1675.435 2913.495 1675.605 ;
        RECT 2913.785 1675.435 2913.955 1675.605 ;
        RECT 5.665 1669.995 5.835 1670.165 ;
        RECT 6.125 1669.995 6.295 1670.165 ;
        RECT 6.585 1669.995 6.755 1670.165 ;
        RECT 2906.425 1669.995 2906.595 1670.165 ;
        RECT 2909.185 1669.995 2909.355 1670.165 ;
        RECT 2909.645 1669.995 2909.815 1670.165 ;
        RECT 2910.105 1669.995 2910.275 1670.165 ;
        RECT 2912.865 1669.995 2913.035 1670.165 ;
        RECT 2913.325 1669.995 2913.495 1670.165 ;
        RECT 2913.785 1669.995 2913.955 1670.165 ;
        RECT 5.665 1664.555 5.835 1664.725 ;
        RECT 6.125 1664.555 6.295 1664.725 ;
        RECT 6.585 1664.555 6.755 1664.725 ;
        RECT 2906.425 1664.555 2906.595 1664.725 ;
        RECT 2912.865 1664.555 2913.035 1664.725 ;
        RECT 2913.325 1664.555 2913.495 1664.725 ;
        RECT 2913.785 1664.555 2913.955 1664.725 ;
        RECT 5.665 1659.115 5.835 1659.285 ;
        RECT 6.125 1659.115 6.295 1659.285 ;
        RECT 6.585 1659.115 6.755 1659.285 ;
        RECT 2906.425 1659.115 2906.595 1659.285 ;
        RECT 2912.865 1659.115 2913.035 1659.285 ;
        RECT 2913.325 1659.115 2913.495 1659.285 ;
        RECT 2913.785 1659.115 2913.955 1659.285 ;
        RECT 5.665 1653.675 5.835 1653.845 ;
        RECT 6.125 1653.675 6.295 1653.845 ;
        RECT 6.585 1653.675 6.755 1653.845 ;
        RECT 2906.425 1653.675 2906.595 1653.845 ;
        RECT 2912.865 1653.675 2913.035 1653.845 ;
        RECT 2913.325 1653.675 2913.495 1653.845 ;
        RECT 2913.785 1653.675 2913.955 1653.845 ;
        RECT 5.665 1648.235 5.835 1648.405 ;
        RECT 6.125 1648.235 6.295 1648.405 ;
        RECT 6.585 1648.235 6.755 1648.405 ;
        RECT 2906.425 1648.235 2906.595 1648.405 ;
        RECT 2912.865 1648.235 2913.035 1648.405 ;
        RECT 2913.325 1648.235 2913.495 1648.405 ;
        RECT 2913.785 1648.235 2913.955 1648.405 ;
        RECT 5.665 1642.795 5.835 1642.965 ;
        RECT 6.125 1642.795 6.295 1642.965 ;
        RECT 6.585 1642.795 6.755 1642.965 ;
        RECT 2906.425 1642.795 2906.595 1642.965 ;
        RECT 2912.865 1642.795 2913.035 1642.965 ;
        RECT 2913.325 1642.795 2913.495 1642.965 ;
        RECT 2913.785 1642.795 2913.955 1642.965 ;
        RECT 5.665 1637.355 5.835 1637.525 ;
        RECT 6.125 1637.355 6.295 1637.525 ;
        RECT 6.585 1637.355 6.755 1637.525 ;
        RECT 2906.425 1637.355 2906.595 1637.525 ;
        RECT 2912.865 1637.355 2913.035 1637.525 ;
        RECT 2913.325 1637.355 2913.495 1637.525 ;
        RECT 2913.785 1637.355 2913.955 1637.525 ;
        RECT 5.665 1631.915 5.835 1632.085 ;
        RECT 6.125 1631.915 6.295 1632.085 ;
        RECT 6.585 1631.915 6.755 1632.085 ;
        RECT 2906.425 1631.915 2906.595 1632.085 ;
        RECT 2912.865 1631.915 2913.035 1632.085 ;
        RECT 2913.325 1631.915 2913.495 1632.085 ;
        RECT 2913.785 1631.915 2913.955 1632.085 ;
        RECT 5.665 1626.475 5.835 1626.645 ;
        RECT 6.125 1626.475 6.295 1626.645 ;
        RECT 6.585 1626.475 6.755 1626.645 ;
        RECT 2906.425 1626.475 2906.595 1626.645 ;
        RECT 2912.865 1626.475 2913.035 1626.645 ;
        RECT 2913.325 1626.475 2913.495 1626.645 ;
        RECT 2913.785 1626.475 2913.955 1626.645 ;
        RECT 5.665 1621.035 5.835 1621.205 ;
        RECT 6.125 1621.035 6.295 1621.205 ;
        RECT 6.585 1621.035 6.755 1621.205 ;
        RECT 2906.425 1621.035 2906.595 1621.205 ;
        RECT 2912.865 1621.035 2913.035 1621.205 ;
        RECT 2913.325 1621.035 2913.495 1621.205 ;
        RECT 2913.785 1621.035 2913.955 1621.205 ;
        RECT 5.665 1615.595 5.835 1615.765 ;
        RECT 6.125 1615.595 6.295 1615.765 ;
        RECT 6.585 1615.595 6.755 1615.765 ;
        RECT 2906.425 1615.595 2906.595 1615.765 ;
        RECT 2912.865 1615.595 2913.035 1615.765 ;
        RECT 2913.325 1615.595 2913.495 1615.765 ;
        RECT 2913.785 1615.595 2913.955 1615.765 ;
        RECT 5.665 1610.155 5.835 1610.325 ;
        RECT 6.125 1610.155 6.295 1610.325 ;
        RECT 6.585 1610.155 6.755 1610.325 ;
        RECT 2906.425 1610.155 2906.595 1610.325 ;
        RECT 2912.865 1610.155 2913.035 1610.325 ;
        RECT 2913.325 1610.155 2913.495 1610.325 ;
        RECT 2913.785 1610.155 2913.955 1610.325 ;
        RECT 5.665 1604.715 5.835 1604.885 ;
        RECT 6.125 1604.715 6.295 1604.885 ;
        RECT 6.585 1604.715 6.755 1604.885 ;
        RECT 2906.425 1604.715 2906.595 1604.885 ;
        RECT 2912.865 1604.715 2913.035 1604.885 ;
        RECT 2913.325 1604.715 2913.495 1604.885 ;
        RECT 2913.785 1604.715 2913.955 1604.885 ;
        RECT 5.665 1599.275 5.835 1599.445 ;
        RECT 6.125 1599.275 6.295 1599.445 ;
        RECT 6.585 1599.275 6.755 1599.445 ;
        RECT 2906.425 1599.275 2906.595 1599.445 ;
        RECT 2912.865 1599.275 2913.035 1599.445 ;
        RECT 2913.325 1599.275 2913.495 1599.445 ;
        RECT 2913.785 1599.275 2913.955 1599.445 ;
        RECT 5.665 1593.835 5.835 1594.005 ;
        RECT 6.125 1593.835 6.295 1594.005 ;
        RECT 6.585 1593.835 6.755 1594.005 ;
        RECT 2906.425 1593.835 2906.595 1594.005 ;
        RECT 2912.865 1593.835 2913.035 1594.005 ;
        RECT 2913.325 1593.835 2913.495 1594.005 ;
        RECT 2913.785 1593.835 2913.955 1594.005 ;
        RECT 5.665 1588.395 5.835 1588.565 ;
        RECT 6.125 1588.395 6.295 1588.565 ;
        RECT 6.585 1588.395 6.755 1588.565 ;
        RECT 2906.425 1588.395 2906.595 1588.565 ;
        RECT 2912.865 1588.395 2913.035 1588.565 ;
        RECT 2913.325 1588.395 2913.495 1588.565 ;
        RECT 2913.785 1588.395 2913.955 1588.565 ;
        RECT 5.665 1582.955 5.835 1583.125 ;
        RECT 6.125 1582.955 6.295 1583.125 ;
        RECT 6.585 1582.955 6.755 1583.125 ;
        RECT 8.885 1582.955 9.055 1583.125 ;
        RECT 9.345 1582.955 9.515 1583.125 ;
        RECT 9.805 1582.955 9.975 1583.125 ;
        RECT 2906.425 1582.955 2906.595 1583.125 ;
        RECT 2912.865 1582.955 2913.035 1583.125 ;
        RECT 2913.325 1582.955 2913.495 1583.125 ;
        RECT 2913.785 1582.955 2913.955 1583.125 ;
        RECT 5.665 1577.515 5.835 1577.685 ;
        RECT 6.125 1577.515 6.295 1577.685 ;
        RECT 6.585 1577.515 6.755 1577.685 ;
        RECT 2906.425 1577.515 2906.595 1577.685 ;
        RECT 2912.865 1577.515 2913.035 1577.685 ;
        RECT 2913.325 1577.515 2913.495 1577.685 ;
        RECT 2913.785 1577.515 2913.955 1577.685 ;
        RECT 5.665 1572.075 5.835 1572.245 ;
        RECT 6.125 1572.075 6.295 1572.245 ;
        RECT 6.585 1572.075 6.755 1572.245 ;
        RECT 2906.425 1572.075 2906.595 1572.245 ;
        RECT 2912.865 1572.075 2913.035 1572.245 ;
        RECT 2913.325 1572.075 2913.495 1572.245 ;
        RECT 2913.785 1572.075 2913.955 1572.245 ;
        RECT 5.665 1566.635 5.835 1566.805 ;
        RECT 6.125 1566.635 6.295 1566.805 ;
        RECT 6.585 1566.635 6.755 1566.805 ;
        RECT 2906.425 1566.635 2906.595 1566.805 ;
        RECT 2912.865 1566.635 2913.035 1566.805 ;
        RECT 2913.325 1566.635 2913.495 1566.805 ;
        RECT 2913.785 1566.635 2913.955 1566.805 ;
        RECT 5.665 1561.195 5.835 1561.365 ;
        RECT 6.125 1561.195 6.295 1561.365 ;
        RECT 6.585 1561.195 6.755 1561.365 ;
        RECT 2906.425 1561.195 2906.595 1561.365 ;
        RECT 2912.865 1561.195 2913.035 1561.365 ;
        RECT 2913.325 1561.195 2913.495 1561.365 ;
        RECT 2913.785 1561.195 2913.955 1561.365 ;
        RECT 5.665 1555.755 5.835 1555.925 ;
        RECT 6.125 1555.755 6.295 1555.925 ;
        RECT 6.585 1555.755 6.755 1555.925 ;
        RECT 2906.425 1555.755 2906.595 1555.925 ;
        RECT 2912.865 1555.755 2913.035 1555.925 ;
        RECT 2913.325 1555.755 2913.495 1555.925 ;
        RECT 2913.785 1555.755 2913.955 1555.925 ;
        RECT 5.665 1550.315 5.835 1550.485 ;
        RECT 6.125 1550.315 6.295 1550.485 ;
        RECT 6.585 1550.315 6.755 1550.485 ;
        RECT 2906.425 1550.315 2906.595 1550.485 ;
        RECT 2912.865 1550.315 2913.035 1550.485 ;
        RECT 2913.325 1550.315 2913.495 1550.485 ;
        RECT 2913.785 1550.315 2913.955 1550.485 ;
        RECT 5.665 1544.875 5.835 1545.045 ;
        RECT 6.125 1544.875 6.295 1545.045 ;
        RECT 6.585 1544.875 6.755 1545.045 ;
        RECT 2906.425 1544.875 2906.595 1545.045 ;
        RECT 2912.865 1544.875 2913.035 1545.045 ;
        RECT 2913.325 1544.875 2913.495 1545.045 ;
        RECT 2913.785 1544.875 2913.955 1545.045 ;
        RECT 5.665 1539.435 5.835 1539.605 ;
        RECT 6.125 1539.435 6.295 1539.605 ;
        RECT 6.585 1539.435 6.755 1539.605 ;
        RECT 2906.425 1539.435 2906.595 1539.605 ;
        RECT 2912.865 1539.435 2913.035 1539.605 ;
        RECT 2913.325 1539.435 2913.495 1539.605 ;
        RECT 2913.785 1539.435 2913.955 1539.605 ;
        RECT 5.665 1533.995 5.835 1534.165 ;
        RECT 6.125 1533.995 6.295 1534.165 ;
        RECT 6.585 1533.995 6.755 1534.165 ;
        RECT 2906.425 1533.995 2906.595 1534.165 ;
        RECT 2912.865 1533.995 2913.035 1534.165 ;
        RECT 2913.325 1533.995 2913.495 1534.165 ;
        RECT 2913.785 1533.995 2913.955 1534.165 ;
        RECT 5.665 1528.555 5.835 1528.725 ;
        RECT 6.125 1528.555 6.295 1528.725 ;
        RECT 6.585 1528.555 6.755 1528.725 ;
        RECT 2906.425 1528.555 2906.595 1528.725 ;
        RECT 2909.185 1528.555 2909.355 1528.725 ;
        RECT 2909.645 1528.555 2909.815 1528.725 ;
        RECT 2910.105 1528.555 2910.275 1528.725 ;
        RECT 2912.865 1528.555 2913.035 1528.725 ;
        RECT 2913.325 1528.555 2913.495 1528.725 ;
        RECT 2913.785 1528.555 2913.955 1528.725 ;
        RECT 5.665 1523.115 5.835 1523.285 ;
        RECT 6.125 1523.115 6.295 1523.285 ;
        RECT 6.585 1523.115 6.755 1523.285 ;
        RECT 2906.425 1523.115 2906.595 1523.285 ;
        RECT 2912.865 1523.115 2913.035 1523.285 ;
        RECT 2913.325 1523.115 2913.495 1523.285 ;
        RECT 2913.785 1523.115 2913.955 1523.285 ;
        RECT 5.665 1517.675 5.835 1517.845 ;
        RECT 6.125 1517.675 6.295 1517.845 ;
        RECT 6.585 1517.675 6.755 1517.845 ;
        RECT 2906.425 1517.675 2906.595 1517.845 ;
        RECT 2909.185 1517.675 2909.355 1517.845 ;
        RECT 2909.645 1517.675 2909.815 1517.845 ;
        RECT 2910.105 1517.675 2910.275 1517.845 ;
        RECT 2912.865 1517.675 2913.035 1517.845 ;
        RECT 2913.325 1517.675 2913.495 1517.845 ;
        RECT 2913.785 1517.675 2913.955 1517.845 ;
        RECT 5.665 1512.235 5.835 1512.405 ;
        RECT 6.125 1512.235 6.295 1512.405 ;
        RECT 6.585 1512.235 6.755 1512.405 ;
        RECT 2906.425 1512.235 2906.595 1512.405 ;
        RECT 2912.865 1512.235 2913.035 1512.405 ;
        RECT 2913.325 1512.235 2913.495 1512.405 ;
        RECT 2913.785 1512.235 2913.955 1512.405 ;
        RECT 5.665 1506.795 5.835 1506.965 ;
        RECT 6.125 1506.795 6.295 1506.965 ;
        RECT 6.585 1506.795 6.755 1506.965 ;
        RECT 2906.425 1506.795 2906.595 1506.965 ;
        RECT 2912.865 1506.795 2913.035 1506.965 ;
        RECT 2913.325 1506.795 2913.495 1506.965 ;
        RECT 2913.785 1506.795 2913.955 1506.965 ;
        RECT 5.665 1501.355 5.835 1501.525 ;
        RECT 6.125 1501.355 6.295 1501.525 ;
        RECT 6.585 1501.355 6.755 1501.525 ;
        RECT 2906.425 1501.355 2906.595 1501.525 ;
        RECT 2912.865 1501.355 2913.035 1501.525 ;
        RECT 2913.325 1501.355 2913.495 1501.525 ;
        RECT 2913.785 1501.355 2913.955 1501.525 ;
        RECT 5.665 1495.915 5.835 1496.085 ;
        RECT 6.125 1495.915 6.295 1496.085 ;
        RECT 6.585 1495.915 6.755 1496.085 ;
        RECT 2906.425 1495.915 2906.595 1496.085 ;
        RECT 2912.865 1495.915 2913.035 1496.085 ;
        RECT 2913.325 1495.915 2913.495 1496.085 ;
        RECT 2913.785 1495.915 2913.955 1496.085 ;
        RECT 5.665 1490.475 5.835 1490.645 ;
        RECT 6.125 1490.475 6.295 1490.645 ;
        RECT 6.585 1490.475 6.755 1490.645 ;
        RECT 2906.425 1490.475 2906.595 1490.645 ;
        RECT 2912.865 1490.475 2913.035 1490.645 ;
        RECT 2913.325 1490.475 2913.495 1490.645 ;
        RECT 2913.785 1490.475 2913.955 1490.645 ;
        RECT 5.665 1485.035 5.835 1485.205 ;
        RECT 6.125 1485.035 6.295 1485.205 ;
        RECT 6.585 1485.035 6.755 1485.205 ;
        RECT 2906.425 1485.035 2906.595 1485.205 ;
        RECT 2912.865 1485.035 2913.035 1485.205 ;
        RECT 2913.325 1485.035 2913.495 1485.205 ;
        RECT 2913.785 1485.035 2913.955 1485.205 ;
        RECT 5.665 1479.595 5.835 1479.765 ;
        RECT 6.125 1479.595 6.295 1479.765 ;
        RECT 6.585 1479.595 6.755 1479.765 ;
        RECT 2906.425 1479.595 2906.595 1479.765 ;
        RECT 2912.865 1479.595 2913.035 1479.765 ;
        RECT 2913.325 1479.595 2913.495 1479.765 ;
        RECT 2913.785 1479.595 2913.955 1479.765 ;
        RECT 5.665 1474.155 5.835 1474.325 ;
        RECT 6.125 1474.155 6.295 1474.325 ;
        RECT 6.585 1474.155 6.755 1474.325 ;
        RECT 2906.425 1474.155 2906.595 1474.325 ;
        RECT 2909.185 1474.155 2909.355 1474.325 ;
        RECT 2909.645 1474.155 2909.815 1474.325 ;
        RECT 2910.105 1474.155 2910.275 1474.325 ;
        RECT 2912.865 1474.155 2913.035 1474.325 ;
        RECT 2913.325 1474.155 2913.495 1474.325 ;
        RECT 2913.785 1474.155 2913.955 1474.325 ;
        RECT 5.665 1468.715 5.835 1468.885 ;
        RECT 6.125 1468.715 6.295 1468.885 ;
        RECT 6.585 1468.715 6.755 1468.885 ;
        RECT 2906.425 1468.715 2906.595 1468.885 ;
        RECT 2912.865 1468.715 2913.035 1468.885 ;
        RECT 2913.325 1468.715 2913.495 1468.885 ;
        RECT 2913.785 1468.715 2913.955 1468.885 ;
        RECT 5.665 1463.275 5.835 1463.445 ;
        RECT 6.125 1463.275 6.295 1463.445 ;
        RECT 6.585 1463.275 6.755 1463.445 ;
        RECT 2906.425 1463.275 2906.595 1463.445 ;
        RECT 2912.865 1463.275 2913.035 1463.445 ;
        RECT 2913.325 1463.275 2913.495 1463.445 ;
        RECT 2913.785 1463.275 2913.955 1463.445 ;
        RECT 5.665 1457.835 5.835 1458.005 ;
        RECT 6.125 1457.835 6.295 1458.005 ;
        RECT 6.585 1457.835 6.755 1458.005 ;
        RECT 2906.425 1457.835 2906.595 1458.005 ;
        RECT 2912.865 1457.835 2913.035 1458.005 ;
        RECT 2913.325 1457.835 2913.495 1458.005 ;
        RECT 2913.785 1457.835 2913.955 1458.005 ;
        RECT 5.665 1452.395 5.835 1452.565 ;
        RECT 6.125 1452.395 6.295 1452.565 ;
        RECT 6.585 1452.395 6.755 1452.565 ;
        RECT 2906.425 1452.395 2906.595 1452.565 ;
        RECT 2912.865 1452.395 2913.035 1452.565 ;
        RECT 2913.325 1452.395 2913.495 1452.565 ;
        RECT 2913.785 1452.395 2913.955 1452.565 ;
        RECT 5.665 1446.955 5.835 1447.125 ;
        RECT 6.125 1446.955 6.295 1447.125 ;
        RECT 6.585 1446.955 6.755 1447.125 ;
        RECT 2906.425 1446.955 2906.595 1447.125 ;
        RECT 2912.865 1446.955 2913.035 1447.125 ;
        RECT 2913.325 1446.955 2913.495 1447.125 ;
        RECT 2913.785 1446.955 2913.955 1447.125 ;
        RECT 5.665 1441.515 5.835 1441.685 ;
        RECT 6.125 1441.515 6.295 1441.685 ;
        RECT 6.585 1441.515 6.755 1441.685 ;
        RECT 2906.425 1441.515 2906.595 1441.685 ;
        RECT 2912.865 1441.515 2913.035 1441.685 ;
        RECT 2913.325 1441.515 2913.495 1441.685 ;
        RECT 2913.785 1441.515 2913.955 1441.685 ;
        RECT 5.665 1436.075 5.835 1436.245 ;
        RECT 6.125 1436.075 6.295 1436.245 ;
        RECT 6.585 1436.075 6.755 1436.245 ;
        RECT 2906.425 1436.075 2906.595 1436.245 ;
        RECT 2912.865 1436.075 2913.035 1436.245 ;
        RECT 2913.325 1436.075 2913.495 1436.245 ;
        RECT 2913.785 1436.075 2913.955 1436.245 ;
        RECT 5.665 1430.635 5.835 1430.805 ;
        RECT 6.125 1430.635 6.295 1430.805 ;
        RECT 6.585 1430.635 6.755 1430.805 ;
        RECT 2906.425 1430.635 2906.595 1430.805 ;
        RECT 2912.865 1430.635 2913.035 1430.805 ;
        RECT 2913.325 1430.635 2913.495 1430.805 ;
        RECT 2913.785 1430.635 2913.955 1430.805 ;
        RECT 5.665 1425.195 5.835 1425.365 ;
        RECT 6.125 1425.195 6.295 1425.365 ;
        RECT 6.585 1425.195 6.755 1425.365 ;
        RECT 2906.425 1425.195 2906.595 1425.365 ;
        RECT 2912.865 1425.195 2913.035 1425.365 ;
        RECT 2913.325 1425.195 2913.495 1425.365 ;
        RECT 2913.785 1425.195 2913.955 1425.365 ;
        RECT 5.665 1419.755 5.835 1419.925 ;
        RECT 6.125 1419.755 6.295 1419.925 ;
        RECT 6.585 1419.755 6.755 1419.925 ;
        RECT 2906.425 1419.755 2906.595 1419.925 ;
        RECT 2912.865 1419.755 2913.035 1419.925 ;
        RECT 2913.325 1419.755 2913.495 1419.925 ;
        RECT 2913.785 1419.755 2913.955 1419.925 ;
        RECT 5.665 1414.315 5.835 1414.485 ;
        RECT 6.125 1414.315 6.295 1414.485 ;
        RECT 6.585 1414.315 6.755 1414.485 ;
        RECT 2906.425 1414.315 2906.595 1414.485 ;
        RECT 2912.865 1414.315 2913.035 1414.485 ;
        RECT 2913.325 1414.315 2913.495 1414.485 ;
        RECT 2913.785 1414.315 2913.955 1414.485 ;
        RECT 5.665 1408.875 5.835 1409.045 ;
        RECT 6.125 1408.875 6.295 1409.045 ;
        RECT 6.585 1408.875 6.755 1409.045 ;
        RECT 2906.425 1408.875 2906.595 1409.045 ;
        RECT 2912.865 1408.875 2913.035 1409.045 ;
        RECT 2913.325 1408.875 2913.495 1409.045 ;
        RECT 2913.785 1408.875 2913.955 1409.045 ;
        RECT 5.665 1403.435 5.835 1403.605 ;
        RECT 6.125 1403.435 6.295 1403.605 ;
        RECT 6.585 1403.435 6.755 1403.605 ;
        RECT 2906.425 1403.435 2906.595 1403.605 ;
        RECT 2912.865 1403.435 2913.035 1403.605 ;
        RECT 2913.325 1403.435 2913.495 1403.605 ;
        RECT 2913.785 1403.435 2913.955 1403.605 ;
        RECT 5.665 1397.995 5.835 1398.165 ;
        RECT 6.125 1397.995 6.295 1398.165 ;
        RECT 6.585 1397.995 6.755 1398.165 ;
        RECT 2906.425 1397.995 2906.595 1398.165 ;
        RECT 2912.865 1397.995 2913.035 1398.165 ;
        RECT 2913.325 1397.995 2913.495 1398.165 ;
        RECT 2913.785 1397.995 2913.955 1398.165 ;
        RECT 5.665 1392.555 5.835 1392.725 ;
        RECT 6.125 1392.555 6.295 1392.725 ;
        RECT 6.585 1392.555 6.755 1392.725 ;
        RECT 2906.425 1392.555 2906.595 1392.725 ;
        RECT 2912.865 1392.555 2913.035 1392.725 ;
        RECT 2913.325 1392.555 2913.495 1392.725 ;
        RECT 2913.785 1392.555 2913.955 1392.725 ;
        RECT 5.665 1387.115 5.835 1387.285 ;
        RECT 6.125 1387.115 6.295 1387.285 ;
        RECT 6.585 1387.115 6.755 1387.285 ;
        RECT 2906.425 1387.115 2906.595 1387.285 ;
        RECT 2912.865 1387.115 2913.035 1387.285 ;
        RECT 2913.325 1387.115 2913.495 1387.285 ;
        RECT 2913.785 1387.115 2913.955 1387.285 ;
        RECT 5.665 1381.675 5.835 1381.845 ;
        RECT 6.125 1381.675 6.295 1381.845 ;
        RECT 6.585 1381.675 6.755 1381.845 ;
        RECT 2906.425 1381.675 2906.595 1381.845 ;
        RECT 2912.865 1381.675 2913.035 1381.845 ;
        RECT 2913.325 1381.675 2913.495 1381.845 ;
        RECT 2913.785 1381.675 2913.955 1381.845 ;
        RECT 5.665 1376.235 5.835 1376.405 ;
        RECT 6.125 1376.235 6.295 1376.405 ;
        RECT 6.585 1376.235 6.755 1376.405 ;
        RECT 2906.425 1376.235 2906.595 1376.405 ;
        RECT 2912.865 1376.235 2913.035 1376.405 ;
        RECT 2913.325 1376.235 2913.495 1376.405 ;
        RECT 2913.785 1376.235 2913.955 1376.405 ;
        RECT 5.665 1370.795 5.835 1370.965 ;
        RECT 6.125 1370.795 6.295 1370.965 ;
        RECT 6.585 1370.795 6.755 1370.965 ;
        RECT 2906.425 1370.795 2906.595 1370.965 ;
        RECT 2912.865 1370.795 2913.035 1370.965 ;
        RECT 2913.325 1370.795 2913.495 1370.965 ;
        RECT 2913.785 1370.795 2913.955 1370.965 ;
        RECT 5.665 1365.355 5.835 1365.525 ;
        RECT 6.125 1365.355 6.295 1365.525 ;
        RECT 6.585 1365.355 6.755 1365.525 ;
        RECT 2906.425 1365.355 2906.595 1365.525 ;
        RECT 2912.865 1365.355 2913.035 1365.525 ;
        RECT 2913.325 1365.355 2913.495 1365.525 ;
        RECT 2913.785 1365.355 2913.955 1365.525 ;
        RECT 5.665 1359.915 5.835 1360.085 ;
        RECT 6.125 1359.915 6.295 1360.085 ;
        RECT 6.585 1359.915 6.755 1360.085 ;
        RECT 2906.425 1359.915 2906.595 1360.085 ;
        RECT 2912.865 1359.915 2913.035 1360.085 ;
        RECT 2913.325 1359.915 2913.495 1360.085 ;
        RECT 2913.785 1359.915 2913.955 1360.085 ;
        RECT 5.665 1354.475 5.835 1354.645 ;
        RECT 6.125 1354.475 6.295 1354.645 ;
        RECT 6.585 1354.475 6.755 1354.645 ;
        RECT 2906.425 1354.475 2906.595 1354.645 ;
        RECT 2912.865 1354.475 2913.035 1354.645 ;
        RECT 2913.325 1354.475 2913.495 1354.645 ;
        RECT 2913.785 1354.475 2913.955 1354.645 ;
        RECT 5.665 1349.035 5.835 1349.205 ;
        RECT 6.125 1349.035 6.295 1349.205 ;
        RECT 6.585 1349.035 6.755 1349.205 ;
        RECT 2906.425 1349.035 2906.595 1349.205 ;
        RECT 2912.865 1349.035 2913.035 1349.205 ;
        RECT 2913.325 1349.035 2913.495 1349.205 ;
        RECT 2913.785 1349.035 2913.955 1349.205 ;
        RECT 5.665 1343.595 5.835 1343.765 ;
        RECT 6.125 1343.595 6.295 1343.765 ;
        RECT 6.585 1343.595 6.755 1343.765 ;
        RECT 2906.425 1343.595 2906.595 1343.765 ;
        RECT 2912.865 1343.595 2913.035 1343.765 ;
        RECT 2913.325 1343.595 2913.495 1343.765 ;
        RECT 2913.785 1343.595 2913.955 1343.765 ;
        RECT 5.665 1338.155 5.835 1338.325 ;
        RECT 6.125 1338.155 6.295 1338.325 ;
        RECT 6.585 1338.155 6.755 1338.325 ;
        RECT 2906.425 1338.155 2906.595 1338.325 ;
        RECT 2912.865 1338.155 2913.035 1338.325 ;
        RECT 2913.325 1338.155 2913.495 1338.325 ;
        RECT 2913.785 1338.155 2913.955 1338.325 ;
        RECT 5.665 1332.715 5.835 1332.885 ;
        RECT 6.125 1332.715 6.295 1332.885 ;
        RECT 6.585 1332.715 6.755 1332.885 ;
        RECT 2906.425 1332.715 2906.595 1332.885 ;
        RECT 2912.865 1332.715 2913.035 1332.885 ;
        RECT 2913.325 1332.715 2913.495 1332.885 ;
        RECT 2913.785 1332.715 2913.955 1332.885 ;
        RECT 5.665 1327.275 5.835 1327.445 ;
        RECT 6.125 1327.275 6.295 1327.445 ;
        RECT 6.585 1327.275 6.755 1327.445 ;
        RECT 8.885 1327.275 9.055 1327.445 ;
        RECT 9.345 1327.275 9.515 1327.445 ;
        RECT 9.805 1327.275 9.975 1327.445 ;
        RECT 2906.425 1327.275 2906.595 1327.445 ;
        RECT 2912.865 1327.275 2913.035 1327.445 ;
        RECT 2913.325 1327.275 2913.495 1327.445 ;
        RECT 2913.785 1327.275 2913.955 1327.445 ;
        RECT 5.665 1321.835 5.835 1322.005 ;
        RECT 6.125 1321.835 6.295 1322.005 ;
        RECT 6.585 1321.835 6.755 1322.005 ;
        RECT 2906.425 1321.835 2906.595 1322.005 ;
        RECT 2912.865 1321.835 2913.035 1322.005 ;
        RECT 2913.325 1321.835 2913.495 1322.005 ;
        RECT 2913.785 1321.835 2913.955 1322.005 ;
        RECT 5.665 1316.395 5.835 1316.565 ;
        RECT 6.125 1316.395 6.295 1316.565 ;
        RECT 6.585 1316.395 6.755 1316.565 ;
        RECT 2906.425 1316.395 2906.595 1316.565 ;
        RECT 2912.865 1316.395 2913.035 1316.565 ;
        RECT 2913.325 1316.395 2913.495 1316.565 ;
        RECT 2913.785 1316.395 2913.955 1316.565 ;
        RECT 5.665 1310.955 5.835 1311.125 ;
        RECT 6.125 1310.955 6.295 1311.125 ;
        RECT 6.585 1310.955 6.755 1311.125 ;
        RECT 2906.425 1310.955 2906.595 1311.125 ;
        RECT 2912.865 1310.955 2913.035 1311.125 ;
        RECT 2913.325 1310.955 2913.495 1311.125 ;
        RECT 2913.785 1310.955 2913.955 1311.125 ;
        RECT 5.665 1305.515 5.835 1305.685 ;
        RECT 6.125 1305.515 6.295 1305.685 ;
        RECT 6.585 1305.515 6.755 1305.685 ;
        RECT 2906.425 1305.515 2906.595 1305.685 ;
        RECT 2912.865 1305.515 2913.035 1305.685 ;
        RECT 2913.325 1305.515 2913.495 1305.685 ;
        RECT 2913.785 1305.515 2913.955 1305.685 ;
        RECT 5.665 1300.075 5.835 1300.245 ;
        RECT 6.125 1300.075 6.295 1300.245 ;
        RECT 6.585 1300.075 6.755 1300.245 ;
        RECT 2906.425 1300.075 2906.595 1300.245 ;
        RECT 2909.185 1300.075 2909.355 1300.245 ;
        RECT 2909.645 1300.075 2909.815 1300.245 ;
        RECT 2910.105 1300.075 2910.275 1300.245 ;
        RECT 2912.865 1300.075 2913.035 1300.245 ;
        RECT 2913.325 1300.075 2913.495 1300.245 ;
        RECT 2913.785 1300.075 2913.955 1300.245 ;
        RECT 5.665 1294.635 5.835 1294.805 ;
        RECT 6.125 1294.635 6.295 1294.805 ;
        RECT 6.585 1294.635 6.755 1294.805 ;
        RECT 2906.425 1294.635 2906.595 1294.805 ;
        RECT 2912.865 1294.635 2913.035 1294.805 ;
        RECT 2913.325 1294.635 2913.495 1294.805 ;
        RECT 2913.785 1294.635 2913.955 1294.805 ;
        RECT 5.665 1289.195 5.835 1289.365 ;
        RECT 6.125 1289.195 6.295 1289.365 ;
        RECT 6.585 1289.195 6.755 1289.365 ;
        RECT 2906.425 1289.195 2906.595 1289.365 ;
        RECT 2912.865 1289.195 2913.035 1289.365 ;
        RECT 2913.325 1289.195 2913.495 1289.365 ;
        RECT 2913.785 1289.195 2913.955 1289.365 ;
        RECT 5.665 1283.755 5.835 1283.925 ;
        RECT 6.125 1283.755 6.295 1283.925 ;
        RECT 6.585 1283.755 6.755 1283.925 ;
        RECT 8.885 1283.755 9.055 1283.925 ;
        RECT 9.345 1283.755 9.515 1283.925 ;
        RECT 9.805 1283.755 9.975 1283.925 ;
        RECT 2906.425 1283.755 2906.595 1283.925 ;
        RECT 2912.865 1283.755 2913.035 1283.925 ;
        RECT 2913.325 1283.755 2913.495 1283.925 ;
        RECT 2913.785 1283.755 2913.955 1283.925 ;
        RECT 5.665 1278.315 5.835 1278.485 ;
        RECT 6.125 1278.315 6.295 1278.485 ;
        RECT 6.585 1278.315 6.755 1278.485 ;
        RECT 2906.425 1278.315 2906.595 1278.485 ;
        RECT 2912.865 1278.315 2913.035 1278.485 ;
        RECT 2913.325 1278.315 2913.495 1278.485 ;
        RECT 2913.785 1278.315 2913.955 1278.485 ;
        RECT 5.665 1272.875 5.835 1273.045 ;
        RECT 6.125 1272.875 6.295 1273.045 ;
        RECT 6.585 1272.875 6.755 1273.045 ;
        RECT 8.885 1272.875 9.055 1273.045 ;
        RECT 9.345 1272.875 9.515 1273.045 ;
        RECT 9.805 1272.875 9.975 1273.045 ;
        RECT 2906.425 1272.875 2906.595 1273.045 ;
        RECT 2912.865 1272.875 2913.035 1273.045 ;
        RECT 2913.325 1272.875 2913.495 1273.045 ;
        RECT 2913.785 1272.875 2913.955 1273.045 ;
        RECT 5.665 1267.435 5.835 1267.605 ;
        RECT 6.125 1267.435 6.295 1267.605 ;
        RECT 6.585 1267.435 6.755 1267.605 ;
        RECT 2906.425 1267.435 2906.595 1267.605 ;
        RECT 2909.185 1267.435 2909.355 1267.605 ;
        RECT 2909.645 1267.435 2909.815 1267.605 ;
        RECT 2910.105 1267.435 2910.275 1267.605 ;
        RECT 2912.865 1267.435 2913.035 1267.605 ;
        RECT 2913.325 1267.435 2913.495 1267.605 ;
        RECT 2913.785 1267.435 2913.955 1267.605 ;
        RECT 5.665 1261.995 5.835 1262.165 ;
        RECT 6.125 1261.995 6.295 1262.165 ;
        RECT 6.585 1261.995 6.755 1262.165 ;
        RECT 2906.425 1261.995 2906.595 1262.165 ;
        RECT 2912.865 1261.995 2913.035 1262.165 ;
        RECT 2913.325 1261.995 2913.495 1262.165 ;
        RECT 2913.785 1261.995 2913.955 1262.165 ;
        RECT 5.665 1256.555 5.835 1256.725 ;
        RECT 6.125 1256.555 6.295 1256.725 ;
        RECT 6.585 1256.555 6.755 1256.725 ;
        RECT 2906.425 1256.555 2906.595 1256.725 ;
        RECT 2912.865 1256.555 2913.035 1256.725 ;
        RECT 2913.325 1256.555 2913.495 1256.725 ;
        RECT 2913.785 1256.555 2913.955 1256.725 ;
        RECT 5.665 1251.115 5.835 1251.285 ;
        RECT 6.125 1251.115 6.295 1251.285 ;
        RECT 6.585 1251.115 6.755 1251.285 ;
        RECT 2906.425 1251.115 2906.595 1251.285 ;
        RECT 2912.865 1251.115 2913.035 1251.285 ;
        RECT 2913.325 1251.115 2913.495 1251.285 ;
        RECT 2913.785 1251.115 2913.955 1251.285 ;
        RECT 5.665 1245.675 5.835 1245.845 ;
        RECT 6.125 1245.675 6.295 1245.845 ;
        RECT 6.585 1245.675 6.755 1245.845 ;
        RECT 2906.425 1245.675 2906.595 1245.845 ;
        RECT 2912.865 1245.675 2913.035 1245.845 ;
        RECT 2913.325 1245.675 2913.495 1245.845 ;
        RECT 2913.785 1245.675 2913.955 1245.845 ;
        RECT 5.665 1240.235 5.835 1240.405 ;
        RECT 6.125 1240.235 6.295 1240.405 ;
        RECT 6.585 1240.235 6.755 1240.405 ;
        RECT 2910.105 1240.235 2910.275 1240.405 ;
        RECT 2912.865 1240.235 2913.035 1240.405 ;
        RECT 2913.325 1240.235 2913.495 1240.405 ;
        RECT 2913.785 1240.235 2913.955 1240.405 ;
        RECT 5.665 1234.795 5.835 1234.965 ;
        RECT 6.125 1234.795 6.295 1234.965 ;
        RECT 6.585 1234.795 6.755 1234.965 ;
        RECT 2910.105 1234.795 2910.275 1234.965 ;
        RECT 2912.865 1234.795 2913.035 1234.965 ;
        RECT 2913.325 1234.795 2913.495 1234.965 ;
        RECT 2913.785 1234.795 2913.955 1234.965 ;
        RECT 5.665 1229.355 5.835 1229.525 ;
        RECT 6.125 1229.355 6.295 1229.525 ;
        RECT 6.585 1229.355 6.755 1229.525 ;
        RECT 2910.105 1229.355 2910.275 1229.525 ;
        RECT 2912.865 1229.355 2913.035 1229.525 ;
        RECT 2913.325 1229.355 2913.495 1229.525 ;
        RECT 2913.785 1229.355 2913.955 1229.525 ;
        RECT 5.665 1223.915 5.835 1224.085 ;
        RECT 6.125 1223.915 6.295 1224.085 ;
        RECT 6.585 1223.915 6.755 1224.085 ;
        RECT 2910.105 1223.915 2910.275 1224.085 ;
        RECT 2912.865 1223.915 2913.035 1224.085 ;
        RECT 2913.325 1223.915 2913.495 1224.085 ;
        RECT 2913.785 1223.915 2913.955 1224.085 ;
        RECT 5.665 1218.475 5.835 1218.645 ;
        RECT 6.125 1218.475 6.295 1218.645 ;
        RECT 6.585 1218.475 6.755 1218.645 ;
        RECT 8.885 1218.475 9.055 1218.645 ;
        RECT 9.345 1218.475 9.515 1218.645 ;
        RECT 9.805 1218.475 9.975 1218.645 ;
        RECT 2910.105 1218.475 2910.275 1218.645 ;
        RECT 2912.865 1218.475 2913.035 1218.645 ;
        RECT 2913.325 1218.475 2913.495 1218.645 ;
        RECT 2913.785 1218.475 2913.955 1218.645 ;
        RECT 5.665 1213.035 5.835 1213.205 ;
        RECT 6.125 1213.035 6.295 1213.205 ;
        RECT 6.585 1213.035 6.755 1213.205 ;
        RECT 2910.105 1213.035 2910.275 1213.205 ;
        RECT 2912.865 1213.035 2913.035 1213.205 ;
        RECT 2913.325 1213.035 2913.495 1213.205 ;
        RECT 2913.785 1213.035 2913.955 1213.205 ;
        RECT 5.665 1207.595 5.835 1207.765 ;
        RECT 6.125 1207.595 6.295 1207.765 ;
        RECT 6.585 1207.595 6.755 1207.765 ;
        RECT 2910.105 1207.595 2910.275 1207.765 ;
        RECT 2912.865 1207.595 2913.035 1207.765 ;
        RECT 2913.325 1207.595 2913.495 1207.765 ;
        RECT 2913.785 1207.595 2913.955 1207.765 ;
        RECT 5.665 1202.155 5.835 1202.325 ;
        RECT 6.125 1202.155 6.295 1202.325 ;
        RECT 6.585 1202.155 6.755 1202.325 ;
        RECT 2910.105 1202.155 2910.275 1202.325 ;
        RECT 2912.865 1202.155 2913.035 1202.325 ;
        RECT 2913.325 1202.155 2913.495 1202.325 ;
        RECT 2913.785 1202.155 2913.955 1202.325 ;
        RECT 5.665 1196.715 5.835 1196.885 ;
        RECT 6.125 1196.715 6.295 1196.885 ;
        RECT 6.585 1196.715 6.755 1196.885 ;
        RECT 2910.105 1196.715 2910.275 1196.885 ;
        RECT 2912.865 1196.715 2913.035 1196.885 ;
        RECT 2913.325 1196.715 2913.495 1196.885 ;
        RECT 2913.785 1196.715 2913.955 1196.885 ;
        RECT 5.665 1191.275 5.835 1191.445 ;
        RECT 6.125 1191.275 6.295 1191.445 ;
        RECT 6.585 1191.275 6.755 1191.445 ;
        RECT 2910.105 1191.275 2910.275 1191.445 ;
        RECT 2912.865 1191.275 2913.035 1191.445 ;
        RECT 2913.325 1191.275 2913.495 1191.445 ;
        RECT 2913.785 1191.275 2913.955 1191.445 ;
        RECT 5.665 1185.835 5.835 1186.005 ;
        RECT 6.125 1185.835 6.295 1186.005 ;
        RECT 6.585 1185.835 6.755 1186.005 ;
        RECT 2910.105 1185.835 2910.275 1186.005 ;
        RECT 2912.865 1185.835 2913.035 1186.005 ;
        RECT 2913.325 1185.835 2913.495 1186.005 ;
        RECT 2913.785 1185.835 2913.955 1186.005 ;
        RECT 5.665 1180.395 5.835 1180.565 ;
        RECT 6.125 1180.395 6.295 1180.565 ;
        RECT 6.585 1180.395 6.755 1180.565 ;
        RECT 2910.105 1180.395 2910.275 1180.565 ;
        RECT 2912.865 1180.395 2913.035 1180.565 ;
        RECT 2913.325 1180.395 2913.495 1180.565 ;
        RECT 2913.785 1180.395 2913.955 1180.565 ;
        RECT 5.665 1174.955 5.835 1175.125 ;
        RECT 6.125 1174.955 6.295 1175.125 ;
        RECT 6.585 1174.955 6.755 1175.125 ;
        RECT 2910.105 1174.955 2910.275 1175.125 ;
        RECT 2912.865 1174.955 2913.035 1175.125 ;
        RECT 2913.325 1174.955 2913.495 1175.125 ;
        RECT 2913.785 1174.955 2913.955 1175.125 ;
        RECT 5.665 1169.515 5.835 1169.685 ;
        RECT 6.125 1169.515 6.295 1169.685 ;
        RECT 6.585 1169.515 6.755 1169.685 ;
        RECT 2910.105 1169.515 2910.275 1169.685 ;
        RECT 2912.865 1169.515 2913.035 1169.685 ;
        RECT 2913.325 1169.515 2913.495 1169.685 ;
        RECT 2913.785 1169.515 2913.955 1169.685 ;
        RECT 5.665 1164.075 5.835 1164.245 ;
        RECT 6.125 1164.075 6.295 1164.245 ;
        RECT 6.585 1164.075 6.755 1164.245 ;
        RECT 2910.105 1164.075 2910.275 1164.245 ;
        RECT 2912.865 1164.075 2913.035 1164.245 ;
        RECT 2913.325 1164.075 2913.495 1164.245 ;
        RECT 2913.785 1164.075 2913.955 1164.245 ;
        RECT 5.665 1158.635 5.835 1158.805 ;
        RECT 6.125 1158.635 6.295 1158.805 ;
        RECT 6.585 1158.635 6.755 1158.805 ;
        RECT 2910.105 1158.635 2910.275 1158.805 ;
        RECT 2912.865 1158.635 2913.035 1158.805 ;
        RECT 2913.325 1158.635 2913.495 1158.805 ;
        RECT 2913.785 1158.635 2913.955 1158.805 ;
        RECT 5.665 1153.195 5.835 1153.365 ;
        RECT 6.125 1153.195 6.295 1153.365 ;
        RECT 6.585 1153.195 6.755 1153.365 ;
        RECT 2910.105 1153.195 2910.275 1153.365 ;
        RECT 2912.865 1153.195 2913.035 1153.365 ;
        RECT 2913.325 1153.195 2913.495 1153.365 ;
        RECT 2913.785 1153.195 2913.955 1153.365 ;
        RECT 5.665 1147.755 5.835 1147.925 ;
        RECT 6.125 1147.755 6.295 1147.925 ;
        RECT 6.585 1147.755 6.755 1147.925 ;
        RECT 2910.105 1147.755 2910.275 1147.925 ;
        RECT 2912.865 1147.755 2913.035 1147.925 ;
        RECT 2913.325 1147.755 2913.495 1147.925 ;
        RECT 2913.785 1147.755 2913.955 1147.925 ;
        RECT 5.665 1142.315 5.835 1142.485 ;
        RECT 6.125 1142.315 6.295 1142.485 ;
        RECT 6.585 1142.315 6.755 1142.485 ;
        RECT 2910.105 1142.315 2910.275 1142.485 ;
        RECT 2912.865 1142.315 2913.035 1142.485 ;
        RECT 2913.325 1142.315 2913.495 1142.485 ;
        RECT 2913.785 1142.315 2913.955 1142.485 ;
        RECT 5.665 1136.875 5.835 1137.045 ;
        RECT 6.125 1136.875 6.295 1137.045 ;
        RECT 6.585 1136.875 6.755 1137.045 ;
        RECT 2910.105 1136.875 2910.275 1137.045 ;
        RECT 2912.865 1136.875 2913.035 1137.045 ;
        RECT 2913.325 1136.875 2913.495 1137.045 ;
        RECT 2913.785 1136.875 2913.955 1137.045 ;
        RECT 5.665 1131.435 5.835 1131.605 ;
        RECT 6.125 1131.435 6.295 1131.605 ;
        RECT 6.585 1131.435 6.755 1131.605 ;
        RECT 2910.105 1131.435 2910.275 1131.605 ;
        RECT 2912.865 1131.435 2913.035 1131.605 ;
        RECT 2913.325 1131.435 2913.495 1131.605 ;
        RECT 2913.785 1131.435 2913.955 1131.605 ;
        RECT 5.665 1125.995 5.835 1126.165 ;
        RECT 6.125 1125.995 6.295 1126.165 ;
        RECT 6.585 1125.995 6.755 1126.165 ;
        RECT 2910.105 1125.995 2910.275 1126.165 ;
        RECT 2912.865 1125.995 2913.035 1126.165 ;
        RECT 2913.325 1125.995 2913.495 1126.165 ;
        RECT 2913.785 1125.995 2913.955 1126.165 ;
        RECT 5.665 1120.555 5.835 1120.725 ;
        RECT 6.125 1120.555 6.295 1120.725 ;
        RECT 6.585 1120.555 6.755 1120.725 ;
        RECT 2910.105 1120.555 2910.275 1120.725 ;
        RECT 2912.865 1120.555 2913.035 1120.725 ;
        RECT 2913.325 1120.555 2913.495 1120.725 ;
        RECT 2913.785 1120.555 2913.955 1120.725 ;
        RECT 5.665 1115.115 5.835 1115.285 ;
        RECT 6.125 1115.115 6.295 1115.285 ;
        RECT 6.585 1115.115 6.755 1115.285 ;
        RECT 2910.105 1115.115 2910.275 1115.285 ;
        RECT 2912.865 1115.115 2913.035 1115.285 ;
        RECT 2913.325 1115.115 2913.495 1115.285 ;
        RECT 2913.785 1115.115 2913.955 1115.285 ;
        RECT 5.665 1109.675 5.835 1109.845 ;
        RECT 6.125 1109.675 6.295 1109.845 ;
        RECT 6.585 1109.675 6.755 1109.845 ;
        RECT 8.885 1109.675 9.055 1109.845 ;
        RECT 9.345 1109.675 9.515 1109.845 ;
        RECT 9.805 1109.675 9.975 1109.845 ;
        RECT 2910.105 1109.675 2910.275 1109.845 ;
        RECT 2912.865 1109.675 2913.035 1109.845 ;
        RECT 2913.325 1109.675 2913.495 1109.845 ;
        RECT 2913.785 1109.675 2913.955 1109.845 ;
        RECT 5.665 1104.235 5.835 1104.405 ;
        RECT 6.125 1104.235 6.295 1104.405 ;
        RECT 6.585 1104.235 6.755 1104.405 ;
        RECT 2910.105 1104.235 2910.275 1104.405 ;
        RECT 2912.865 1104.235 2913.035 1104.405 ;
        RECT 2913.325 1104.235 2913.495 1104.405 ;
        RECT 2913.785 1104.235 2913.955 1104.405 ;
        RECT 5.665 1098.795 5.835 1098.965 ;
        RECT 6.125 1098.795 6.295 1098.965 ;
        RECT 6.585 1098.795 6.755 1098.965 ;
        RECT 2910.105 1098.795 2910.275 1098.965 ;
        RECT 2912.865 1098.795 2913.035 1098.965 ;
        RECT 2913.325 1098.795 2913.495 1098.965 ;
        RECT 2913.785 1098.795 2913.955 1098.965 ;
        RECT 5.665 1093.355 5.835 1093.525 ;
        RECT 6.125 1093.355 6.295 1093.525 ;
        RECT 6.585 1093.355 6.755 1093.525 ;
        RECT 2910.105 1093.355 2910.275 1093.525 ;
        RECT 2912.865 1093.355 2913.035 1093.525 ;
        RECT 2913.325 1093.355 2913.495 1093.525 ;
        RECT 2913.785 1093.355 2913.955 1093.525 ;
        RECT 5.665 1087.915 5.835 1088.085 ;
        RECT 6.125 1087.915 6.295 1088.085 ;
        RECT 6.585 1087.915 6.755 1088.085 ;
        RECT 2910.105 1087.915 2910.275 1088.085 ;
        RECT 2912.865 1087.915 2913.035 1088.085 ;
        RECT 2913.325 1087.915 2913.495 1088.085 ;
        RECT 2913.785 1087.915 2913.955 1088.085 ;
        RECT 5.665 1082.475 5.835 1082.645 ;
        RECT 6.125 1082.475 6.295 1082.645 ;
        RECT 6.585 1082.475 6.755 1082.645 ;
        RECT 2910.105 1082.475 2910.275 1082.645 ;
        RECT 2912.865 1082.475 2913.035 1082.645 ;
        RECT 2913.325 1082.475 2913.495 1082.645 ;
        RECT 2913.785 1082.475 2913.955 1082.645 ;
        RECT 5.665 1077.035 5.835 1077.205 ;
        RECT 6.125 1077.035 6.295 1077.205 ;
        RECT 6.585 1077.035 6.755 1077.205 ;
        RECT 2910.105 1077.035 2910.275 1077.205 ;
        RECT 2912.865 1077.035 2913.035 1077.205 ;
        RECT 2913.325 1077.035 2913.495 1077.205 ;
        RECT 2913.785 1077.035 2913.955 1077.205 ;
        RECT 5.665 1071.595 5.835 1071.765 ;
        RECT 6.125 1071.595 6.295 1071.765 ;
        RECT 6.585 1071.595 6.755 1071.765 ;
        RECT 2910.105 1071.595 2910.275 1071.765 ;
        RECT 2912.865 1071.595 2913.035 1071.765 ;
        RECT 2913.325 1071.595 2913.495 1071.765 ;
        RECT 2913.785 1071.595 2913.955 1071.765 ;
        RECT 5.665 1066.155 5.835 1066.325 ;
        RECT 6.125 1066.155 6.295 1066.325 ;
        RECT 6.585 1066.155 6.755 1066.325 ;
        RECT 2910.105 1066.155 2910.275 1066.325 ;
        RECT 2912.865 1066.155 2913.035 1066.325 ;
        RECT 2913.325 1066.155 2913.495 1066.325 ;
        RECT 2913.785 1066.155 2913.955 1066.325 ;
        RECT 5.665 1060.715 5.835 1060.885 ;
        RECT 6.125 1060.715 6.295 1060.885 ;
        RECT 6.585 1060.715 6.755 1060.885 ;
        RECT 2910.105 1060.715 2910.275 1060.885 ;
        RECT 2912.865 1060.715 2913.035 1060.885 ;
        RECT 2913.325 1060.715 2913.495 1060.885 ;
        RECT 2913.785 1060.715 2913.955 1060.885 ;
        RECT 5.665 1055.275 5.835 1055.445 ;
        RECT 6.125 1055.275 6.295 1055.445 ;
        RECT 6.585 1055.275 6.755 1055.445 ;
        RECT 2910.105 1055.275 2910.275 1055.445 ;
        RECT 2912.865 1055.275 2913.035 1055.445 ;
        RECT 2913.325 1055.275 2913.495 1055.445 ;
        RECT 2913.785 1055.275 2913.955 1055.445 ;
        RECT 5.665 1049.835 5.835 1050.005 ;
        RECT 6.125 1049.835 6.295 1050.005 ;
        RECT 6.585 1049.835 6.755 1050.005 ;
        RECT 2910.105 1049.835 2910.275 1050.005 ;
        RECT 2912.865 1049.835 2913.035 1050.005 ;
        RECT 2913.325 1049.835 2913.495 1050.005 ;
        RECT 2913.785 1049.835 2913.955 1050.005 ;
        RECT 5.665 1044.395 5.835 1044.565 ;
        RECT 6.125 1044.395 6.295 1044.565 ;
        RECT 6.585 1044.395 6.755 1044.565 ;
        RECT 2910.105 1044.395 2910.275 1044.565 ;
        RECT 2912.865 1044.395 2913.035 1044.565 ;
        RECT 2913.325 1044.395 2913.495 1044.565 ;
        RECT 2913.785 1044.395 2913.955 1044.565 ;
        RECT 5.665 1038.955 5.835 1039.125 ;
        RECT 6.125 1038.955 6.295 1039.125 ;
        RECT 6.585 1038.955 6.755 1039.125 ;
        RECT 2910.105 1038.955 2910.275 1039.125 ;
        RECT 2912.865 1038.955 2913.035 1039.125 ;
        RECT 2913.325 1038.955 2913.495 1039.125 ;
        RECT 2913.785 1038.955 2913.955 1039.125 ;
        RECT 5.665 1033.515 5.835 1033.685 ;
        RECT 6.125 1033.515 6.295 1033.685 ;
        RECT 6.585 1033.515 6.755 1033.685 ;
        RECT 8.885 1033.515 9.055 1033.685 ;
        RECT 9.345 1033.515 9.515 1033.685 ;
        RECT 9.805 1033.515 9.975 1033.685 ;
        RECT 2910.105 1033.515 2910.275 1033.685 ;
        RECT 2912.865 1033.515 2913.035 1033.685 ;
        RECT 2913.325 1033.515 2913.495 1033.685 ;
        RECT 2913.785 1033.515 2913.955 1033.685 ;
        RECT 5.665 1028.075 5.835 1028.245 ;
        RECT 6.125 1028.075 6.295 1028.245 ;
        RECT 6.585 1028.075 6.755 1028.245 ;
        RECT 2910.105 1028.075 2910.275 1028.245 ;
        RECT 2912.865 1028.075 2913.035 1028.245 ;
        RECT 2913.325 1028.075 2913.495 1028.245 ;
        RECT 2913.785 1028.075 2913.955 1028.245 ;
        RECT 5.665 1022.635 5.835 1022.805 ;
        RECT 6.125 1022.635 6.295 1022.805 ;
        RECT 6.585 1022.635 6.755 1022.805 ;
        RECT 2910.105 1022.635 2910.275 1022.805 ;
        RECT 2912.865 1022.635 2913.035 1022.805 ;
        RECT 2913.325 1022.635 2913.495 1022.805 ;
        RECT 2913.785 1022.635 2913.955 1022.805 ;
        RECT 5.665 1017.195 5.835 1017.365 ;
        RECT 6.125 1017.195 6.295 1017.365 ;
        RECT 6.585 1017.195 6.755 1017.365 ;
        RECT 2910.105 1017.195 2910.275 1017.365 ;
        RECT 2912.865 1017.195 2913.035 1017.365 ;
        RECT 2913.325 1017.195 2913.495 1017.365 ;
        RECT 2913.785 1017.195 2913.955 1017.365 ;
        RECT 5.665 1011.755 5.835 1011.925 ;
        RECT 6.125 1011.755 6.295 1011.925 ;
        RECT 6.585 1011.755 6.755 1011.925 ;
        RECT 2910.105 1011.755 2910.275 1011.925 ;
        RECT 2912.865 1011.755 2913.035 1011.925 ;
        RECT 2913.325 1011.755 2913.495 1011.925 ;
        RECT 2913.785 1011.755 2913.955 1011.925 ;
        RECT 5.665 1006.315 5.835 1006.485 ;
        RECT 6.125 1006.315 6.295 1006.485 ;
        RECT 6.585 1006.315 6.755 1006.485 ;
        RECT 2909.185 1006.315 2909.355 1006.485 ;
        RECT 2909.645 1006.315 2909.815 1006.485 ;
        RECT 2910.105 1006.315 2910.275 1006.485 ;
        RECT 2912.865 1006.315 2913.035 1006.485 ;
        RECT 2913.325 1006.315 2913.495 1006.485 ;
        RECT 2913.785 1006.315 2913.955 1006.485 ;
        RECT 5.665 1000.875 5.835 1001.045 ;
        RECT 6.125 1000.875 6.295 1001.045 ;
        RECT 6.585 1000.875 6.755 1001.045 ;
        RECT 2910.105 1000.875 2910.275 1001.045 ;
        RECT 2912.865 1000.875 2913.035 1001.045 ;
        RECT 2913.325 1000.875 2913.495 1001.045 ;
        RECT 2913.785 1000.875 2913.955 1001.045 ;
        RECT 5.665 995.435 5.835 995.605 ;
        RECT 6.125 995.435 6.295 995.605 ;
        RECT 6.585 995.435 6.755 995.605 ;
        RECT 2909.185 995.435 2909.355 995.605 ;
        RECT 2909.645 995.435 2909.815 995.605 ;
        RECT 2910.105 995.435 2910.275 995.605 ;
        RECT 2912.865 995.435 2913.035 995.605 ;
        RECT 2913.325 995.435 2913.495 995.605 ;
        RECT 2913.785 995.435 2913.955 995.605 ;
        RECT 5.665 989.995 5.835 990.165 ;
        RECT 6.125 989.995 6.295 990.165 ;
        RECT 6.585 989.995 6.755 990.165 ;
        RECT 2910.105 989.995 2910.275 990.165 ;
        RECT 2912.865 989.995 2913.035 990.165 ;
        RECT 2913.325 989.995 2913.495 990.165 ;
        RECT 2913.785 989.995 2913.955 990.165 ;
        RECT 5.665 984.555 5.835 984.725 ;
        RECT 6.125 984.555 6.295 984.725 ;
        RECT 6.585 984.555 6.755 984.725 ;
        RECT 2910.105 984.555 2910.275 984.725 ;
        RECT 2912.865 984.555 2913.035 984.725 ;
        RECT 2913.325 984.555 2913.495 984.725 ;
        RECT 2913.785 984.555 2913.955 984.725 ;
        RECT 5.665 979.115 5.835 979.285 ;
        RECT 6.125 979.115 6.295 979.285 ;
        RECT 6.585 979.115 6.755 979.285 ;
        RECT 2910.105 979.115 2910.275 979.285 ;
        RECT 2912.865 979.115 2913.035 979.285 ;
        RECT 2913.325 979.115 2913.495 979.285 ;
        RECT 2913.785 979.115 2913.955 979.285 ;
        RECT 5.665 973.675 5.835 973.845 ;
        RECT 6.125 973.675 6.295 973.845 ;
        RECT 6.585 973.675 6.755 973.845 ;
        RECT 2910.105 973.675 2910.275 973.845 ;
        RECT 2912.865 973.675 2913.035 973.845 ;
        RECT 2913.325 973.675 2913.495 973.845 ;
        RECT 2913.785 973.675 2913.955 973.845 ;
        RECT 5.665 968.235 5.835 968.405 ;
        RECT 6.125 968.235 6.295 968.405 ;
        RECT 6.585 968.235 6.755 968.405 ;
        RECT 2910.105 968.235 2910.275 968.405 ;
        RECT 2912.865 968.235 2913.035 968.405 ;
        RECT 2913.325 968.235 2913.495 968.405 ;
        RECT 2913.785 968.235 2913.955 968.405 ;
        RECT 5.665 962.795 5.835 962.965 ;
        RECT 6.125 962.795 6.295 962.965 ;
        RECT 6.585 962.795 6.755 962.965 ;
        RECT 2910.105 962.795 2910.275 962.965 ;
        RECT 2912.865 962.795 2913.035 962.965 ;
        RECT 2913.325 962.795 2913.495 962.965 ;
        RECT 2913.785 962.795 2913.955 962.965 ;
        RECT 5.665 957.355 5.835 957.525 ;
        RECT 6.125 957.355 6.295 957.525 ;
        RECT 6.585 957.355 6.755 957.525 ;
        RECT 2910.105 957.355 2910.275 957.525 ;
        RECT 2912.865 957.355 2913.035 957.525 ;
        RECT 2913.325 957.355 2913.495 957.525 ;
        RECT 2913.785 957.355 2913.955 957.525 ;
        RECT 5.665 951.915 5.835 952.085 ;
        RECT 6.125 951.915 6.295 952.085 ;
        RECT 6.585 951.915 6.755 952.085 ;
        RECT 2910.105 951.915 2910.275 952.085 ;
        RECT 2912.865 951.915 2913.035 952.085 ;
        RECT 2913.325 951.915 2913.495 952.085 ;
        RECT 2913.785 951.915 2913.955 952.085 ;
        RECT 5.665 946.475 5.835 946.645 ;
        RECT 6.125 946.475 6.295 946.645 ;
        RECT 6.585 946.475 6.755 946.645 ;
        RECT 2910.105 946.475 2910.275 946.645 ;
        RECT 2912.865 946.475 2913.035 946.645 ;
        RECT 2913.325 946.475 2913.495 946.645 ;
        RECT 2913.785 946.475 2913.955 946.645 ;
        RECT 5.665 941.035 5.835 941.205 ;
        RECT 6.125 941.035 6.295 941.205 ;
        RECT 6.585 941.035 6.755 941.205 ;
        RECT 2910.105 941.035 2910.275 941.205 ;
        RECT 2912.865 941.035 2913.035 941.205 ;
        RECT 2913.325 941.035 2913.495 941.205 ;
        RECT 2913.785 941.035 2913.955 941.205 ;
        RECT 5.665 935.595 5.835 935.765 ;
        RECT 6.125 935.595 6.295 935.765 ;
        RECT 6.585 935.595 6.755 935.765 ;
        RECT 2910.105 935.595 2910.275 935.765 ;
        RECT 2912.865 935.595 2913.035 935.765 ;
        RECT 2913.325 935.595 2913.495 935.765 ;
        RECT 2913.785 935.595 2913.955 935.765 ;
        RECT 5.665 930.155 5.835 930.325 ;
        RECT 6.125 930.155 6.295 930.325 ;
        RECT 6.585 930.155 6.755 930.325 ;
        RECT 2910.105 930.155 2910.275 930.325 ;
        RECT 2912.865 930.155 2913.035 930.325 ;
        RECT 2913.325 930.155 2913.495 930.325 ;
        RECT 2913.785 930.155 2913.955 930.325 ;
        RECT 5.665 924.715 5.835 924.885 ;
        RECT 6.125 924.715 6.295 924.885 ;
        RECT 6.585 924.715 6.755 924.885 ;
        RECT 2910.105 924.715 2910.275 924.885 ;
        RECT 2912.865 924.715 2913.035 924.885 ;
        RECT 2913.325 924.715 2913.495 924.885 ;
        RECT 2913.785 924.715 2913.955 924.885 ;
        RECT 5.665 919.275 5.835 919.445 ;
        RECT 6.125 919.275 6.295 919.445 ;
        RECT 6.585 919.275 6.755 919.445 ;
        RECT 2910.105 919.275 2910.275 919.445 ;
        RECT 2912.865 919.275 2913.035 919.445 ;
        RECT 2913.325 919.275 2913.495 919.445 ;
        RECT 2913.785 919.275 2913.955 919.445 ;
        RECT 5.665 913.835 5.835 914.005 ;
        RECT 6.125 913.835 6.295 914.005 ;
        RECT 6.585 913.835 6.755 914.005 ;
        RECT 2910.105 913.835 2910.275 914.005 ;
        RECT 2912.865 913.835 2913.035 914.005 ;
        RECT 2913.325 913.835 2913.495 914.005 ;
        RECT 2913.785 913.835 2913.955 914.005 ;
        RECT 5.665 908.395 5.835 908.565 ;
        RECT 6.125 908.395 6.295 908.565 ;
        RECT 6.585 908.395 6.755 908.565 ;
        RECT 2910.105 908.395 2910.275 908.565 ;
        RECT 2912.865 908.395 2913.035 908.565 ;
        RECT 2913.325 908.395 2913.495 908.565 ;
        RECT 2913.785 908.395 2913.955 908.565 ;
        RECT 5.665 902.955 5.835 903.125 ;
        RECT 6.125 902.955 6.295 903.125 ;
        RECT 6.585 902.955 6.755 903.125 ;
        RECT 2910.105 902.955 2910.275 903.125 ;
        RECT 2912.865 902.955 2913.035 903.125 ;
        RECT 2913.325 902.955 2913.495 903.125 ;
        RECT 2913.785 902.955 2913.955 903.125 ;
        RECT 5.665 897.515 5.835 897.685 ;
        RECT 6.125 897.515 6.295 897.685 ;
        RECT 6.585 897.515 6.755 897.685 ;
        RECT 2910.105 897.515 2910.275 897.685 ;
        RECT 2912.865 897.515 2913.035 897.685 ;
        RECT 2913.325 897.515 2913.495 897.685 ;
        RECT 2913.785 897.515 2913.955 897.685 ;
        RECT 5.665 892.075 5.835 892.245 ;
        RECT 6.125 892.075 6.295 892.245 ;
        RECT 6.585 892.075 6.755 892.245 ;
        RECT 2910.105 892.075 2910.275 892.245 ;
        RECT 2912.865 892.075 2913.035 892.245 ;
        RECT 2913.325 892.075 2913.495 892.245 ;
        RECT 2913.785 892.075 2913.955 892.245 ;
        RECT 5.665 886.635 5.835 886.805 ;
        RECT 6.125 886.635 6.295 886.805 ;
        RECT 6.585 886.635 6.755 886.805 ;
        RECT 2910.105 886.635 2910.275 886.805 ;
        RECT 2912.865 886.635 2913.035 886.805 ;
        RECT 2913.325 886.635 2913.495 886.805 ;
        RECT 2913.785 886.635 2913.955 886.805 ;
        RECT 5.665 881.195 5.835 881.365 ;
        RECT 6.125 881.195 6.295 881.365 ;
        RECT 6.585 881.195 6.755 881.365 ;
        RECT 2910.105 881.195 2910.275 881.365 ;
        RECT 2912.865 881.195 2913.035 881.365 ;
        RECT 2913.325 881.195 2913.495 881.365 ;
        RECT 2913.785 881.195 2913.955 881.365 ;
        RECT 5.665 875.755 5.835 875.925 ;
        RECT 6.125 875.755 6.295 875.925 ;
        RECT 6.585 875.755 6.755 875.925 ;
        RECT 2910.105 875.755 2910.275 875.925 ;
        RECT 2912.865 875.755 2913.035 875.925 ;
        RECT 2913.325 875.755 2913.495 875.925 ;
        RECT 2913.785 875.755 2913.955 875.925 ;
        RECT 5.665 870.315 5.835 870.485 ;
        RECT 6.125 870.315 6.295 870.485 ;
        RECT 6.585 870.315 6.755 870.485 ;
        RECT 2910.105 870.315 2910.275 870.485 ;
        RECT 2912.865 870.315 2913.035 870.485 ;
        RECT 2913.325 870.315 2913.495 870.485 ;
        RECT 2913.785 870.315 2913.955 870.485 ;
        RECT 5.665 864.875 5.835 865.045 ;
        RECT 6.125 864.875 6.295 865.045 ;
        RECT 6.585 864.875 6.755 865.045 ;
        RECT 2910.105 864.875 2910.275 865.045 ;
        RECT 2912.865 864.875 2913.035 865.045 ;
        RECT 2913.325 864.875 2913.495 865.045 ;
        RECT 2913.785 864.875 2913.955 865.045 ;
        RECT 5.665 859.435 5.835 859.605 ;
        RECT 6.125 859.435 6.295 859.605 ;
        RECT 6.585 859.435 6.755 859.605 ;
        RECT 2910.105 859.435 2910.275 859.605 ;
        RECT 2912.865 859.435 2913.035 859.605 ;
        RECT 2913.325 859.435 2913.495 859.605 ;
        RECT 2913.785 859.435 2913.955 859.605 ;
        RECT 5.665 853.995 5.835 854.165 ;
        RECT 6.125 853.995 6.295 854.165 ;
        RECT 6.585 853.995 6.755 854.165 ;
        RECT 2910.105 853.995 2910.275 854.165 ;
        RECT 2912.865 853.995 2913.035 854.165 ;
        RECT 2913.325 853.995 2913.495 854.165 ;
        RECT 2913.785 853.995 2913.955 854.165 ;
        RECT 5.665 848.555 5.835 848.725 ;
        RECT 6.125 848.555 6.295 848.725 ;
        RECT 6.585 848.555 6.755 848.725 ;
        RECT 2910.105 848.555 2910.275 848.725 ;
        RECT 2912.865 848.555 2913.035 848.725 ;
        RECT 2913.325 848.555 2913.495 848.725 ;
        RECT 2913.785 848.555 2913.955 848.725 ;
        RECT 5.665 843.115 5.835 843.285 ;
        RECT 6.125 843.115 6.295 843.285 ;
        RECT 6.585 843.115 6.755 843.285 ;
        RECT 2910.105 843.115 2910.275 843.285 ;
        RECT 2912.865 843.115 2913.035 843.285 ;
        RECT 2913.325 843.115 2913.495 843.285 ;
        RECT 2913.785 843.115 2913.955 843.285 ;
        RECT 5.665 837.675 5.835 837.845 ;
        RECT 6.125 837.675 6.295 837.845 ;
        RECT 6.585 837.675 6.755 837.845 ;
        RECT 2910.105 837.675 2910.275 837.845 ;
        RECT 2912.865 837.675 2913.035 837.845 ;
        RECT 2913.325 837.675 2913.495 837.845 ;
        RECT 2913.785 837.675 2913.955 837.845 ;
        RECT 5.665 832.235 5.835 832.405 ;
        RECT 6.125 832.235 6.295 832.405 ;
        RECT 6.585 832.235 6.755 832.405 ;
        RECT 2910.105 832.235 2910.275 832.405 ;
        RECT 2912.865 832.235 2913.035 832.405 ;
        RECT 2913.325 832.235 2913.495 832.405 ;
        RECT 2913.785 832.235 2913.955 832.405 ;
        RECT 5.665 826.795 5.835 826.965 ;
        RECT 6.125 826.795 6.295 826.965 ;
        RECT 6.585 826.795 6.755 826.965 ;
        RECT 2910.105 826.795 2910.275 826.965 ;
        RECT 2912.865 826.795 2913.035 826.965 ;
        RECT 2913.325 826.795 2913.495 826.965 ;
        RECT 2913.785 826.795 2913.955 826.965 ;
        RECT 5.665 821.355 5.835 821.525 ;
        RECT 6.125 821.355 6.295 821.525 ;
        RECT 6.585 821.355 6.755 821.525 ;
        RECT 2910.105 821.355 2910.275 821.525 ;
        RECT 2912.865 821.355 2913.035 821.525 ;
        RECT 2913.325 821.355 2913.495 821.525 ;
        RECT 2913.785 821.355 2913.955 821.525 ;
        RECT 5.665 815.915 5.835 816.085 ;
        RECT 6.125 815.915 6.295 816.085 ;
        RECT 6.585 815.915 6.755 816.085 ;
        RECT 2910.105 815.915 2910.275 816.085 ;
        RECT 2912.865 815.915 2913.035 816.085 ;
        RECT 2913.325 815.915 2913.495 816.085 ;
        RECT 2913.785 815.915 2913.955 816.085 ;
        RECT 5.665 810.475 5.835 810.645 ;
        RECT 6.125 810.475 6.295 810.645 ;
        RECT 6.585 810.475 6.755 810.645 ;
        RECT 2909.185 810.475 2909.355 810.645 ;
        RECT 2909.645 810.475 2909.815 810.645 ;
        RECT 2910.105 810.475 2910.275 810.645 ;
        RECT 2912.865 810.475 2913.035 810.645 ;
        RECT 2913.325 810.475 2913.495 810.645 ;
        RECT 2913.785 810.475 2913.955 810.645 ;
        RECT 5.665 805.035 5.835 805.205 ;
        RECT 6.125 805.035 6.295 805.205 ;
        RECT 6.585 805.035 6.755 805.205 ;
        RECT 2910.105 805.035 2910.275 805.205 ;
        RECT 2912.865 805.035 2913.035 805.205 ;
        RECT 2913.325 805.035 2913.495 805.205 ;
        RECT 2913.785 805.035 2913.955 805.205 ;
        RECT 5.665 799.595 5.835 799.765 ;
        RECT 6.125 799.595 6.295 799.765 ;
        RECT 6.585 799.595 6.755 799.765 ;
        RECT 2910.105 799.595 2910.275 799.765 ;
        RECT 2912.865 799.595 2913.035 799.765 ;
        RECT 2913.325 799.595 2913.495 799.765 ;
        RECT 2913.785 799.595 2913.955 799.765 ;
        RECT 5.665 794.155 5.835 794.325 ;
        RECT 6.125 794.155 6.295 794.325 ;
        RECT 6.585 794.155 6.755 794.325 ;
        RECT 2910.105 794.155 2910.275 794.325 ;
        RECT 2912.865 794.155 2913.035 794.325 ;
        RECT 2913.325 794.155 2913.495 794.325 ;
        RECT 2913.785 794.155 2913.955 794.325 ;
        RECT 5.665 788.715 5.835 788.885 ;
        RECT 6.125 788.715 6.295 788.885 ;
        RECT 6.585 788.715 6.755 788.885 ;
        RECT 2910.105 788.715 2910.275 788.885 ;
        RECT 2912.865 788.715 2913.035 788.885 ;
        RECT 2913.325 788.715 2913.495 788.885 ;
        RECT 2913.785 788.715 2913.955 788.885 ;
        RECT 5.665 783.275 5.835 783.445 ;
        RECT 6.125 783.275 6.295 783.445 ;
        RECT 6.585 783.275 6.755 783.445 ;
        RECT 2910.105 783.275 2910.275 783.445 ;
        RECT 2912.865 783.275 2913.035 783.445 ;
        RECT 2913.325 783.275 2913.495 783.445 ;
        RECT 2913.785 783.275 2913.955 783.445 ;
        RECT 5.665 777.835 5.835 778.005 ;
        RECT 6.125 777.835 6.295 778.005 ;
        RECT 6.585 777.835 6.755 778.005 ;
        RECT 2910.105 777.835 2910.275 778.005 ;
        RECT 2912.865 777.835 2913.035 778.005 ;
        RECT 2913.325 777.835 2913.495 778.005 ;
        RECT 2913.785 777.835 2913.955 778.005 ;
        RECT 5.665 772.395 5.835 772.565 ;
        RECT 6.125 772.395 6.295 772.565 ;
        RECT 6.585 772.395 6.755 772.565 ;
        RECT 2910.105 772.395 2910.275 772.565 ;
        RECT 2912.865 772.395 2913.035 772.565 ;
        RECT 2913.325 772.395 2913.495 772.565 ;
        RECT 2913.785 772.395 2913.955 772.565 ;
        RECT 5.665 766.955 5.835 767.125 ;
        RECT 6.125 766.955 6.295 767.125 ;
        RECT 6.585 766.955 6.755 767.125 ;
        RECT 2910.105 766.955 2910.275 767.125 ;
        RECT 2912.865 766.955 2913.035 767.125 ;
        RECT 2913.325 766.955 2913.495 767.125 ;
        RECT 2913.785 766.955 2913.955 767.125 ;
        RECT 5.665 761.515 5.835 761.685 ;
        RECT 6.125 761.515 6.295 761.685 ;
        RECT 6.585 761.515 6.755 761.685 ;
        RECT 2910.105 761.515 2910.275 761.685 ;
        RECT 2912.865 761.515 2913.035 761.685 ;
        RECT 2913.325 761.515 2913.495 761.685 ;
        RECT 2913.785 761.515 2913.955 761.685 ;
        RECT 5.665 756.075 5.835 756.245 ;
        RECT 6.125 756.075 6.295 756.245 ;
        RECT 6.585 756.075 6.755 756.245 ;
        RECT 2910.105 756.075 2910.275 756.245 ;
        RECT 2912.865 756.075 2913.035 756.245 ;
        RECT 2913.325 756.075 2913.495 756.245 ;
        RECT 2913.785 756.075 2913.955 756.245 ;
        RECT 5.665 750.635 5.835 750.805 ;
        RECT 6.125 750.635 6.295 750.805 ;
        RECT 6.585 750.635 6.755 750.805 ;
        RECT 2910.105 750.635 2910.275 750.805 ;
        RECT 2912.865 750.635 2913.035 750.805 ;
        RECT 2913.325 750.635 2913.495 750.805 ;
        RECT 2913.785 750.635 2913.955 750.805 ;
        RECT 5.665 745.195 5.835 745.365 ;
        RECT 6.125 745.195 6.295 745.365 ;
        RECT 6.585 745.195 6.755 745.365 ;
        RECT 2910.105 745.195 2910.275 745.365 ;
        RECT 2912.865 745.195 2913.035 745.365 ;
        RECT 2913.325 745.195 2913.495 745.365 ;
        RECT 2913.785 745.195 2913.955 745.365 ;
        RECT 5.665 739.755 5.835 739.925 ;
        RECT 6.125 739.755 6.295 739.925 ;
        RECT 6.585 739.755 6.755 739.925 ;
        RECT 2910.105 739.755 2910.275 739.925 ;
        RECT 2912.865 739.755 2913.035 739.925 ;
        RECT 2913.325 739.755 2913.495 739.925 ;
        RECT 2913.785 739.755 2913.955 739.925 ;
        RECT 5.665 734.315 5.835 734.485 ;
        RECT 6.125 734.315 6.295 734.485 ;
        RECT 6.585 734.315 6.755 734.485 ;
        RECT 2909.185 734.315 2909.355 734.485 ;
        RECT 2909.645 734.315 2909.815 734.485 ;
        RECT 2910.105 734.315 2910.275 734.485 ;
        RECT 2912.865 734.315 2913.035 734.485 ;
        RECT 2913.325 734.315 2913.495 734.485 ;
        RECT 2913.785 734.315 2913.955 734.485 ;
        RECT 5.665 728.875 5.835 729.045 ;
        RECT 6.125 728.875 6.295 729.045 ;
        RECT 6.585 728.875 6.755 729.045 ;
        RECT 2910.105 728.875 2910.275 729.045 ;
        RECT 2912.865 728.875 2913.035 729.045 ;
        RECT 2913.325 728.875 2913.495 729.045 ;
        RECT 2913.785 728.875 2913.955 729.045 ;
        RECT 5.665 723.435 5.835 723.605 ;
        RECT 6.125 723.435 6.295 723.605 ;
        RECT 6.585 723.435 6.755 723.605 ;
        RECT 8.885 723.435 9.055 723.605 ;
        RECT 9.345 723.435 9.515 723.605 ;
        RECT 9.805 723.435 9.975 723.605 ;
        RECT 2910.105 723.435 2910.275 723.605 ;
        RECT 2912.865 723.435 2913.035 723.605 ;
        RECT 2913.325 723.435 2913.495 723.605 ;
        RECT 2913.785 723.435 2913.955 723.605 ;
        RECT 5.665 717.995 5.835 718.165 ;
        RECT 6.125 717.995 6.295 718.165 ;
        RECT 6.585 717.995 6.755 718.165 ;
        RECT 2910.105 717.995 2910.275 718.165 ;
        RECT 2912.865 717.995 2913.035 718.165 ;
        RECT 2913.325 717.995 2913.495 718.165 ;
        RECT 2913.785 717.995 2913.955 718.165 ;
        RECT 5.665 712.555 5.835 712.725 ;
        RECT 6.125 712.555 6.295 712.725 ;
        RECT 6.585 712.555 6.755 712.725 ;
        RECT 2910.105 712.555 2910.275 712.725 ;
        RECT 2912.865 712.555 2913.035 712.725 ;
        RECT 2913.325 712.555 2913.495 712.725 ;
        RECT 2913.785 712.555 2913.955 712.725 ;
        RECT 5.665 707.115 5.835 707.285 ;
        RECT 6.125 707.115 6.295 707.285 ;
        RECT 6.585 707.115 6.755 707.285 ;
        RECT 2910.105 707.115 2910.275 707.285 ;
        RECT 2912.865 707.115 2913.035 707.285 ;
        RECT 2913.325 707.115 2913.495 707.285 ;
        RECT 2913.785 707.115 2913.955 707.285 ;
        RECT 5.665 701.675 5.835 701.845 ;
        RECT 6.125 701.675 6.295 701.845 ;
        RECT 6.585 701.675 6.755 701.845 ;
        RECT 2910.105 701.675 2910.275 701.845 ;
        RECT 2912.865 701.675 2913.035 701.845 ;
        RECT 2913.325 701.675 2913.495 701.845 ;
        RECT 2913.785 701.675 2913.955 701.845 ;
        RECT 5.665 696.235 5.835 696.405 ;
        RECT 6.125 696.235 6.295 696.405 ;
        RECT 6.585 696.235 6.755 696.405 ;
        RECT 2910.105 696.235 2910.275 696.405 ;
        RECT 2912.865 696.235 2913.035 696.405 ;
        RECT 2913.325 696.235 2913.495 696.405 ;
        RECT 2913.785 696.235 2913.955 696.405 ;
        RECT 5.665 690.795 5.835 690.965 ;
        RECT 6.125 690.795 6.295 690.965 ;
        RECT 6.585 690.795 6.755 690.965 ;
        RECT 2910.105 690.795 2910.275 690.965 ;
        RECT 2912.865 690.795 2913.035 690.965 ;
        RECT 2913.325 690.795 2913.495 690.965 ;
        RECT 2913.785 690.795 2913.955 690.965 ;
        RECT 5.665 685.355 5.835 685.525 ;
        RECT 6.125 685.355 6.295 685.525 ;
        RECT 6.585 685.355 6.755 685.525 ;
        RECT 2910.105 685.355 2910.275 685.525 ;
        RECT 2912.865 685.355 2913.035 685.525 ;
        RECT 2913.325 685.355 2913.495 685.525 ;
        RECT 2913.785 685.355 2913.955 685.525 ;
        RECT 5.665 679.915 5.835 680.085 ;
        RECT 6.125 679.915 6.295 680.085 ;
        RECT 6.585 679.915 6.755 680.085 ;
        RECT 2910.105 679.915 2910.275 680.085 ;
        RECT 2912.865 679.915 2913.035 680.085 ;
        RECT 2913.325 679.915 2913.495 680.085 ;
        RECT 2913.785 679.915 2913.955 680.085 ;
        RECT 5.665 674.475 5.835 674.645 ;
        RECT 6.125 674.475 6.295 674.645 ;
        RECT 6.585 674.475 6.755 674.645 ;
        RECT 2910.105 674.475 2910.275 674.645 ;
        RECT 2912.865 674.475 2913.035 674.645 ;
        RECT 2913.325 674.475 2913.495 674.645 ;
        RECT 2913.785 674.475 2913.955 674.645 ;
        RECT 5.665 669.035 5.835 669.205 ;
        RECT 6.125 669.035 6.295 669.205 ;
        RECT 6.585 669.035 6.755 669.205 ;
        RECT 2910.105 669.035 2910.275 669.205 ;
        RECT 2912.865 669.035 2913.035 669.205 ;
        RECT 2913.325 669.035 2913.495 669.205 ;
        RECT 2913.785 669.035 2913.955 669.205 ;
        RECT 5.665 663.595 5.835 663.765 ;
        RECT 6.125 663.595 6.295 663.765 ;
        RECT 6.585 663.595 6.755 663.765 ;
        RECT 2910.105 663.595 2910.275 663.765 ;
        RECT 2912.865 663.595 2913.035 663.765 ;
        RECT 2913.325 663.595 2913.495 663.765 ;
        RECT 2913.785 663.595 2913.955 663.765 ;
        RECT 5.665 658.155 5.835 658.325 ;
        RECT 6.125 658.155 6.295 658.325 ;
        RECT 6.585 658.155 6.755 658.325 ;
        RECT 2910.105 658.155 2910.275 658.325 ;
        RECT 2912.865 658.155 2913.035 658.325 ;
        RECT 2913.325 658.155 2913.495 658.325 ;
        RECT 2913.785 658.155 2913.955 658.325 ;
        RECT 5.665 652.715 5.835 652.885 ;
        RECT 6.125 652.715 6.295 652.885 ;
        RECT 6.585 652.715 6.755 652.885 ;
        RECT 2910.105 652.715 2910.275 652.885 ;
        RECT 2912.865 652.715 2913.035 652.885 ;
        RECT 2913.325 652.715 2913.495 652.885 ;
        RECT 2913.785 652.715 2913.955 652.885 ;
        RECT 5.665 647.275 5.835 647.445 ;
        RECT 6.125 647.275 6.295 647.445 ;
        RECT 6.585 647.275 6.755 647.445 ;
        RECT 2910.105 647.275 2910.275 647.445 ;
        RECT 2912.865 647.275 2913.035 647.445 ;
        RECT 2913.325 647.275 2913.495 647.445 ;
        RECT 2913.785 647.275 2913.955 647.445 ;
        RECT 5.665 641.835 5.835 642.005 ;
        RECT 6.125 641.835 6.295 642.005 ;
        RECT 6.585 641.835 6.755 642.005 ;
        RECT 2910.105 641.835 2910.275 642.005 ;
        RECT 2912.865 641.835 2913.035 642.005 ;
        RECT 2913.325 641.835 2913.495 642.005 ;
        RECT 2913.785 641.835 2913.955 642.005 ;
        RECT 5.665 636.395 5.835 636.565 ;
        RECT 6.125 636.395 6.295 636.565 ;
        RECT 6.585 636.395 6.755 636.565 ;
        RECT 2910.105 636.395 2910.275 636.565 ;
        RECT 2912.865 636.395 2913.035 636.565 ;
        RECT 2913.325 636.395 2913.495 636.565 ;
        RECT 2913.785 636.395 2913.955 636.565 ;
        RECT 5.665 630.955 5.835 631.125 ;
        RECT 6.125 630.955 6.295 631.125 ;
        RECT 6.585 630.955 6.755 631.125 ;
        RECT 8.885 630.955 9.055 631.125 ;
        RECT 9.345 630.955 9.515 631.125 ;
        RECT 9.805 630.955 9.975 631.125 ;
        RECT 2910.105 630.955 2910.275 631.125 ;
        RECT 2912.865 630.955 2913.035 631.125 ;
        RECT 2913.325 630.955 2913.495 631.125 ;
        RECT 2913.785 630.955 2913.955 631.125 ;
        RECT 5.665 625.515 5.835 625.685 ;
        RECT 6.125 625.515 6.295 625.685 ;
        RECT 6.585 625.515 6.755 625.685 ;
        RECT 2910.105 625.515 2910.275 625.685 ;
        RECT 2912.865 625.515 2913.035 625.685 ;
        RECT 2913.325 625.515 2913.495 625.685 ;
        RECT 2913.785 625.515 2913.955 625.685 ;
        RECT 5.665 620.075 5.835 620.245 ;
        RECT 6.125 620.075 6.295 620.245 ;
        RECT 6.585 620.075 6.755 620.245 ;
        RECT 2910.105 620.075 2910.275 620.245 ;
        RECT 2912.865 620.075 2913.035 620.245 ;
        RECT 2913.325 620.075 2913.495 620.245 ;
        RECT 2913.785 620.075 2913.955 620.245 ;
        RECT 5.665 614.635 5.835 614.805 ;
        RECT 6.125 614.635 6.295 614.805 ;
        RECT 6.585 614.635 6.755 614.805 ;
        RECT 2910.105 614.635 2910.275 614.805 ;
        RECT 2912.865 614.635 2913.035 614.805 ;
        RECT 2913.325 614.635 2913.495 614.805 ;
        RECT 2913.785 614.635 2913.955 614.805 ;
        RECT 5.665 609.195 5.835 609.365 ;
        RECT 6.125 609.195 6.295 609.365 ;
        RECT 6.585 609.195 6.755 609.365 ;
        RECT 2910.105 609.195 2910.275 609.365 ;
        RECT 2912.865 609.195 2913.035 609.365 ;
        RECT 2913.325 609.195 2913.495 609.365 ;
        RECT 2913.785 609.195 2913.955 609.365 ;
        RECT 5.665 603.755 5.835 603.925 ;
        RECT 6.125 603.755 6.295 603.925 ;
        RECT 6.585 603.755 6.755 603.925 ;
        RECT 8.885 603.755 9.055 603.925 ;
        RECT 9.345 603.755 9.515 603.925 ;
        RECT 9.805 603.755 9.975 603.925 ;
        RECT 2910.105 603.755 2910.275 603.925 ;
        RECT 2912.865 603.755 2913.035 603.925 ;
        RECT 2913.325 603.755 2913.495 603.925 ;
        RECT 2913.785 603.755 2913.955 603.925 ;
        RECT 5.665 598.315 5.835 598.485 ;
        RECT 6.125 598.315 6.295 598.485 ;
        RECT 6.585 598.315 6.755 598.485 ;
        RECT 2910.105 598.315 2910.275 598.485 ;
        RECT 2912.865 598.315 2913.035 598.485 ;
        RECT 2913.325 598.315 2913.495 598.485 ;
        RECT 2913.785 598.315 2913.955 598.485 ;
        RECT 5.665 592.875 5.835 593.045 ;
        RECT 6.125 592.875 6.295 593.045 ;
        RECT 6.585 592.875 6.755 593.045 ;
        RECT 2910.105 592.875 2910.275 593.045 ;
        RECT 2912.865 592.875 2913.035 593.045 ;
        RECT 2913.325 592.875 2913.495 593.045 ;
        RECT 2913.785 592.875 2913.955 593.045 ;
        RECT 5.665 587.435 5.835 587.605 ;
        RECT 6.125 587.435 6.295 587.605 ;
        RECT 6.585 587.435 6.755 587.605 ;
        RECT 2910.105 587.435 2910.275 587.605 ;
        RECT 2912.865 587.435 2913.035 587.605 ;
        RECT 2913.325 587.435 2913.495 587.605 ;
        RECT 2913.785 587.435 2913.955 587.605 ;
        RECT 5.665 581.995 5.835 582.165 ;
        RECT 6.125 581.995 6.295 582.165 ;
        RECT 6.585 581.995 6.755 582.165 ;
        RECT 2910.105 581.995 2910.275 582.165 ;
        RECT 2912.865 581.995 2913.035 582.165 ;
        RECT 2913.325 581.995 2913.495 582.165 ;
        RECT 2913.785 581.995 2913.955 582.165 ;
        RECT 5.665 576.555 5.835 576.725 ;
        RECT 6.125 576.555 6.295 576.725 ;
        RECT 6.585 576.555 6.755 576.725 ;
        RECT 2910.105 576.555 2910.275 576.725 ;
        RECT 2912.865 576.555 2913.035 576.725 ;
        RECT 2913.325 576.555 2913.495 576.725 ;
        RECT 2913.785 576.555 2913.955 576.725 ;
        RECT 5.665 571.115 5.835 571.285 ;
        RECT 6.125 571.115 6.295 571.285 ;
        RECT 6.585 571.115 6.755 571.285 ;
        RECT 2910.105 571.115 2910.275 571.285 ;
        RECT 2912.865 571.115 2913.035 571.285 ;
        RECT 2913.325 571.115 2913.495 571.285 ;
        RECT 2913.785 571.115 2913.955 571.285 ;
        RECT 5.665 565.675 5.835 565.845 ;
        RECT 6.125 565.675 6.295 565.845 ;
        RECT 6.585 565.675 6.755 565.845 ;
        RECT 2910.105 565.675 2910.275 565.845 ;
        RECT 2912.865 565.675 2913.035 565.845 ;
        RECT 2913.325 565.675 2913.495 565.845 ;
        RECT 2913.785 565.675 2913.955 565.845 ;
        RECT 5.665 560.235 5.835 560.405 ;
        RECT 6.125 560.235 6.295 560.405 ;
        RECT 6.585 560.235 6.755 560.405 ;
        RECT 2910.105 560.235 2910.275 560.405 ;
        RECT 2912.865 560.235 2913.035 560.405 ;
        RECT 2913.325 560.235 2913.495 560.405 ;
        RECT 2913.785 560.235 2913.955 560.405 ;
        RECT 5.665 554.795 5.835 554.965 ;
        RECT 6.125 554.795 6.295 554.965 ;
        RECT 6.585 554.795 6.755 554.965 ;
        RECT 2910.105 554.795 2910.275 554.965 ;
        RECT 2912.865 554.795 2913.035 554.965 ;
        RECT 2913.325 554.795 2913.495 554.965 ;
        RECT 2913.785 554.795 2913.955 554.965 ;
        RECT 5.665 549.355 5.835 549.525 ;
        RECT 6.125 549.355 6.295 549.525 ;
        RECT 6.585 549.355 6.755 549.525 ;
        RECT 2910.105 549.355 2910.275 549.525 ;
        RECT 2912.865 549.355 2913.035 549.525 ;
        RECT 2913.325 549.355 2913.495 549.525 ;
        RECT 2913.785 549.355 2913.955 549.525 ;
        RECT 5.665 543.915 5.835 544.085 ;
        RECT 6.125 543.915 6.295 544.085 ;
        RECT 6.585 543.915 6.755 544.085 ;
        RECT 2910.105 543.915 2910.275 544.085 ;
        RECT 2912.865 543.915 2913.035 544.085 ;
        RECT 2913.325 543.915 2913.495 544.085 ;
        RECT 2913.785 543.915 2913.955 544.085 ;
        RECT 5.665 538.475 5.835 538.645 ;
        RECT 6.125 538.475 6.295 538.645 ;
        RECT 6.585 538.475 6.755 538.645 ;
        RECT 2910.105 538.475 2910.275 538.645 ;
        RECT 2912.865 538.475 2913.035 538.645 ;
        RECT 2913.325 538.475 2913.495 538.645 ;
        RECT 2913.785 538.475 2913.955 538.645 ;
        RECT 5.665 533.035 5.835 533.205 ;
        RECT 6.125 533.035 6.295 533.205 ;
        RECT 6.585 533.035 6.755 533.205 ;
        RECT 2910.105 533.035 2910.275 533.205 ;
        RECT 2912.865 533.035 2913.035 533.205 ;
        RECT 2913.325 533.035 2913.495 533.205 ;
        RECT 2913.785 533.035 2913.955 533.205 ;
        RECT 5.665 527.595 5.835 527.765 ;
        RECT 6.125 527.595 6.295 527.765 ;
        RECT 6.585 527.595 6.755 527.765 ;
        RECT 2910.105 527.595 2910.275 527.765 ;
        RECT 2912.865 527.595 2913.035 527.765 ;
        RECT 2913.325 527.595 2913.495 527.765 ;
        RECT 2913.785 527.595 2913.955 527.765 ;
        RECT 5.665 522.155 5.835 522.325 ;
        RECT 6.125 522.155 6.295 522.325 ;
        RECT 6.585 522.155 6.755 522.325 ;
        RECT 2910.105 522.155 2910.275 522.325 ;
        RECT 2912.865 522.155 2913.035 522.325 ;
        RECT 2913.325 522.155 2913.495 522.325 ;
        RECT 2913.785 522.155 2913.955 522.325 ;
        RECT 5.665 516.715 5.835 516.885 ;
        RECT 6.125 516.715 6.295 516.885 ;
        RECT 6.585 516.715 6.755 516.885 ;
        RECT 2910.105 516.715 2910.275 516.885 ;
        RECT 2912.865 516.715 2913.035 516.885 ;
        RECT 2913.325 516.715 2913.495 516.885 ;
        RECT 2913.785 516.715 2913.955 516.885 ;
        RECT 5.665 511.275 5.835 511.445 ;
        RECT 6.125 511.275 6.295 511.445 ;
        RECT 6.585 511.275 6.755 511.445 ;
        RECT 2910.105 511.275 2910.275 511.445 ;
        RECT 2912.865 511.275 2913.035 511.445 ;
        RECT 2913.325 511.275 2913.495 511.445 ;
        RECT 2913.785 511.275 2913.955 511.445 ;
        RECT 5.665 505.835 5.835 506.005 ;
        RECT 6.125 505.835 6.295 506.005 ;
        RECT 6.585 505.835 6.755 506.005 ;
        RECT 2910.105 505.835 2910.275 506.005 ;
        RECT 2912.865 505.835 2913.035 506.005 ;
        RECT 2913.325 505.835 2913.495 506.005 ;
        RECT 2913.785 505.835 2913.955 506.005 ;
        RECT 5.665 500.395 5.835 500.565 ;
        RECT 6.125 500.395 6.295 500.565 ;
        RECT 6.585 500.395 6.755 500.565 ;
        RECT 2910.105 500.395 2910.275 500.565 ;
        RECT 2912.865 500.395 2913.035 500.565 ;
        RECT 2913.325 500.395 2913.495 500.565 ;
        RECT 2913.785 500.395 2913.955 500.565 ;
        RECT 5.665 494.955 5.835 495.125 ;
        RECT 6.125 494.955 6.295 495.125 ;
        RECT 6.585 494.955 6.755 495.125 ;
        RECT 2910.105 494.955 2910.275 495.125 ;
        RECT 2912.865 494.955 2913.035 495.125 ;
        RECT 2913.325 494.955 2913.495 495.125 ;
        RECT 2913.785 494.955 2913.955 495.125 ;
        RECT 5.665 489.515 5.835 489.685 ;
        RECT 6.125 489.515 6.295 489.685 ;
        RECT 6.585 489.515 6.755 489.685 ;
        RECT 2910.105 489.515 2910.275 489.685 ;
        RECT 2912.865 489.515 2913.035 489.685 ;
        RECT 2913.325 489.515 2913.495 489.685 ;
        RECT 2913.785 489.515 2913.955 489.685 ;
        RECT 5.665 484.075 5.835 484.245 ;
        RECT 6.125 484.075 6.295 484.245 ;
        RECT 6.585 484.075 6.755 484.245 ;
        RECT 2910.105 484.075 2910.275 484.245 ;
        RECT 2912.865 484.075 2913.035 484.245 ;
        RECT 2913.325 484.075 2913.495 484.245 ;
        RECT 2913.785 484.075 2913.955 484.245 ;
        RECT 5.665 478.635 5.835 478.805 ;
        RECT 6.125 478.635 6.295 478.805 ;
        RECT 6.585 478.635 6.755 478.805 ;
        RECT 2910.105 478.635 2910.275 478.805 ;
        RECT 2912.865 478.635 2913.035 478.805 ;
        RECT 2913.325 478.635 2913.495 478.805 ;
        RECT 2913.785 478.635 2913.955 478.805 ;
        RECT 5.665 473.195 5.835 473.365 ;
        RECT 6.125 473.195 6.295 473.365 ;
        RECT 6.585 473.195 6.755 473.365 ;
        RECT 2910.105 473.195 2910.275 473.365 ;
        RECT 2912.865 473.195 2913.035 473.365 ;
        RECT 2913.325 473.195 2913.495 473.365 ;
        RECT 2913.785 473.195 2913.955 473.365 ;
        RECT 5.665 467.755 5.835 467.925 ;
        RECT 6.125 467.755 6.295 467.925 ;
        RECT 6.585 467.755 6.755 467.925 ;
        RECT 2909.185 467.755 2909.355 467.925 ;
        RECT 2909.645 467.755 2909.815 467.925 ;
        RECT 2910.105 467.755 2910.275 467.925 ;
        RECT 2912.865 467.755 2913.035 467.925 ;
        RECT 2913.325 467.755 2913.495 467.925 ;
        RECT 2913.785 467.755 2913.955 467.925 ;
        RECT 5.665 462.315 5.835 462.485 ;
        RECT 6.125 462.315 6.295 462.485 ;
        RECT 6.585 462.315 6.755 462.485 ;
        RECT 2910.105 462.315 2910.275 462.485 ;
        RECT 2912.865 462.315 2913.035 462.485 ;
        RECT 2913.325 462.315 2913.495 462.485 ;
        RECT 2913.785 462.315 2913.955 462.485 ;
        RECT 5.665 456.875 5.835 457.045 ;
        RECT 6.125 456.875 6.295 457.045 ;
        RECT 6.585 456.875 6.755 457.045 ;
        RECT 2910.105 456.875 2910.275 457.045 ;
        RECT 2912.865 456.875 2913.035 457.045 ;
        RECT 2913.325 456.875 2913.495 457.045 ;
        RECT 2913.785 456.875 2913.955 457.045 ;
        RECT 5.665 451.435 5.835 451.605 ;
        RECT 6.125 451.435 6.295 451.605 ;
        RECT 6.585 451.435 6.755 451.605 ;
        RECT 2910.105 451.435 2910.275 451.605 ;
        RECT 2910.565 451.435 2910.735 451.605 ;
        RECT 2911.025 451.435 2911.195 451.605 ;
        RECT 2911.485 451.435 2911.655 451.605 ;
        RECT 2912.865 451.435 2913.035 451.605 ;
        RECT 2913.325 451.435 2913.495 451.605 ;
        RECT 2913.785 451.435 2913.955 451.605 ;
        RECT 5.665 445.995 5.835 446.165 ;
        RECT 6.125 445.995 6.295 446.165 ;
        RECT 6.585 445.995 6.755 446.165 ;
        RECT 2910.105 445.995 2910.275 446.165 ;
        RECT 2912.865 445.995 2913.035 446.165 ;
        RECT 2913.325 445.995 2913.495 446.165 ;
        RECT 2913.785 445.995 2913.955 446.165 ;
        RECT 5.665 440.555 5.835 440.725 ;
        RECT 6.125 440.555 6.295 440.725 ;
        RECT 6.585 440.555 6.755 440.725 ;
        RECT 8.885 440.555 9.055 440.725 ;
        RECT 9.345 440.555 9.515 440.725 ;
        RECT 9.805 440.555 9.975 440.725 ;
        RECT 2910.105 440.555 2910.275 440.725 ;
        RECT 2912.865 440.555 2913.035 440.725 ;
        RECT 2913.325 440.555 2913.495 440.725 ;
        RECT 2913.785 440.555 2913.955 440.725 ;
        RECT 5.665 435.115 5.835 435.285 ;
        RECT 6.125 435.115 6.295 435.285 ;
        RECT 6.585 435.115 6.755 435.285 ;
        RECT 2910.105 435.115 2910.275 435.285 ;
        RECT 2912.865 435.115 2913.035 435.285 ;
        RECT 2913.325 435.115 2913.495 435.285 ;
        RECT 2913.785 435.115 2913.955 435.285 ;
        RECT 5.665 429.675 5.835 429.845 ;
        RECT 6.125 429.675 6.295 429.845 ;
        RECT 6.585 429.675 6.755 429.845 ;
        RECT 2910.105 429.675 2910.275 429.845 ;
        RECT 2912.865 429.675 2913.035 429.845 ;
        RECT 2913.325 429.675 2913.495 429.845 ;
        RECT 2913.785 429.675 2913.955 429.845 ;
        RECT 5.665 424.235 5.835 424.405 ;
        RECT 6.125 424.235 6.295 424.405 ;
        RECT 6.585 424.235 6.755 424.405 ;
        RECT 2910.105 424.235 2910.275 424.405 ;
        RECT 2912.865 424.235 2913.035 424.405 ;
        RECT 2913.325 424.235 2913.495 424.405 ;
        RECT 2913.785 424.235 2913.955 424.405 ;
        RECT 5.665 418.795 5.835 418.965 ;
        RECT 6.125 418.795 6.295 418.965 ;
        RECT 6.585 418.795 6.755 418.965 ;
        RECT 2910.105 418.795 2910.275 418.965 ;
        RECT 2912.865 418.795 2913.035 418.965 ;
        RECT 2913.325 418.795 2913.495 418.965 ;
        RECT 2913.785 418.795 2913.955 418.965 ;
        RECT 5.665 413.355 5.835 413.525 ;
        RECT 6.125 413.355 6.295 413.525 ;
        RECT 6.585 413.355 6.755 413.525 ;
        RECT 2910.105 413.355 2910.275 413.525 ;
        RECT 2912.865 413.355 2913.035 413.525 ;
        RECT 2913.325 413.355 2913.495 413.525 ;
        RECT 2913.785 413.355 2913.955 413.525 ;
        RECT 5.665 407.915 5.835 408.085 ;
        RECT 6.125 407.915 6.295 408.085 ;
        RECT 6.585 407.915 6.755 408.085 ;
        RECT 2910.105 407.915 2910.275 408.085 ;
        RECT 2912.865 407.915 2913.035 408.085 ;
        RECT 2913.325 407.915 2913.495 408.085 ;
        RECT 2913.785 407.915 2913.955 408.085 ;
        RECT 5.665 402.475 5.835 402.645 ;
        RECT 6.125 402.475 6.295 402.645 ;
        RECT 6.585 402.475 6.755 402.645 ;
        RECT 8.885 402.475 9.055 402.645 ;
        RECT 9.345 402.475 9.515 402.645 ;
        RECT 9.805 402.475 9.975 402.645 ;
        RECT 2910.105 402.475 2910.275 402.645 ;
        RECT 2912.865 402.475 2913.035 402.645 ;
        RECT 2913.325 402.475 2913.495 402.645 ;
        RECT 2913.785 402.475 2913.955 402.645 ;
        RECT 5.665 397.035 5.835 397.205 ;
        RECT 6.125 397.035 6.295 397.205 ;
        RECT 6.585 397.035 6.755 397.205 ;
        RECT 2910.105 397.035 2910.275 397.205 ;
        RECT 2912.865 397.035 2913.035 397.205 ;
        RECT 2913.325 397.035 2913.495 397.205 ;
        RECT 2913.785 397.035 2913.955 397.205 ;
        RECT 5.665 391.595 5.835 391.765 ;
        RECT 6.125 391.595 6.295 391.765 ;
        RECT 6.585 391.595 6.755 391.765 ;
        RECT 8.885 391.595 9.055 391.765 ;
        RECT 9.345 391.595 9.515 391.765 ;
        RECT 9.805 391.595 9.975 391.765 ;
        RECT 2910.105 391.595 2910.275 391.765 ;
        RECT 2912.865 391.595 2913.035 391.765 ;
        RECT 2913.325 391.595 2913.495 391.765 ;
        RECT 2913.785 391.595 2913.955 391.765 ;
        RECT 5.665 386.155 5.835 386.325 ;
        RECT 6.125 386.155 6.295 386.325 ;
        RECT 6.585 386.155 6.755 386.325 ;
        RECT 2910.105 386.155 2910.275 386.325 ;
        RECT 2912.865 386.155 2913.035 386.325 ;
        RECT 2913.325 386.155 2913.495 386.325 ;
        RECT 2913.785 386.155 2913.955 386.325 ;
        RECT 5.665 380.715 5.835 380.885 ;
        RECT 6.125 380.715 6.295 380.885 ;
        RECT 6.585 380.715 6.755 380.885 ;
        RECT 2910.105 380.715 2910.275 380.885 ;
        RECT 2912.865 380.715 2913.035 380.885 ;
        RECT 2913.325 380.715 2913.495 380.885 ;
        RECT 2913.785 380.715 2913.955 380.885 ;
        RECT 5.665 375.275 5.835 375.445 ;
        RECT 6.125 375.275 6.295 375.445 ;
        RECT 6.585 375.275 6.755 375.445 ;
        RECT 2910.105 375.275 2910.275 375.445 ;
        RECT 2912.865 375.275 2913.035 375.445 ;
        RECT 2913.325 375.275 2913.495 375.445 ;
        RECT 2913.785 375.275 2913.955 375.445 ;
        RECT 5.665 369.835 5.835 370.005 ;
        RECT 6.125 369.835 6.295 370.005 ;
        RECT 6.585 369.835 6.755 370.005 ;
        RECT 2910.105 369.835 2910.275 370.005 ;
        RECT 2912.865 369.835 2913.035 370.005 ;
        RECT 2913.325 369.835 2913.495 370.005 ;
        RECT 2913.785 369.835 2913.955 370.005 ;
        RECT 5.665 364.395 5.835 364.565 ;
        RECT 6.125 364.395 6.295 364.565 ;
        RECT 6.585 364.395 6.755 364.565 ;
        RECT 2910.105 364.395 2910.275 364.565 ;
        RECT 2912.865 364.395 2913.035 364.565 ;
        RECT 2913.325 364.395 2913.495 364.565 ;
        RECT 2913.785 364.395 2913.955 364.565 ;
        RECT 5.665 358.955 5.835 359.125 ;
        RECT 6.125 358.955 6.295 359.125 ;
        RECT 6.585 358.955 6.755 359.125 ;
        RECT 2910.105 358.955 2910.275 359.125 ;
        RECT 2912.865 358.955 2913.035 359.125 ;
        RECT 2913.325 358.955 2913.495 359.125 ;
        RECT 2913.785 358.955 2913.955 359.125 ;
        RECT 5.665 353.515 5.835 353.685 ;
        RECT 6.125 353.515 6.295 353.685 ;
        RECT 6.585 353.515 6.755 353.685 ;
        RECT 2910.105 353.515 2910.275 353.685 ;
        RECT 2912.865 353.515 2913.035 353.685 ;
        RECT 2913.325 353.515 2913.495 353.685 ;
        RECT 2913.785 353.515 2913.955 353.685 ;
        RECT 5.665 348.075 5.835 348.245 ;
        RECT 6.125 348.075 6.295 348.245 ;
        RECT 6.585 348.075 6.755 348.245 ;
        RECT 2910.105 348.075 2910.275 348.245 ;
        RECT 2912.865 348.075 2913.035 348.245 ;
        RECT 2913.325 348.075 2913.495 348.245 ;
        RECT 2913.785 348.075 2913.955 348.245 ;
        RECT 5.665 342.635 5.835 342.805 ;
        RECT 6.125 342.635 6.295 342.805 ;
        RECT 6.585 342.635 6.755 342.805 ;
        RECT 2910.105 342.635 2910.275 342.805 ;
        RECT 2912.865 342.635 2913.035 342.805 ;
        RECT 2913.325 342.635 2913.495 342.805 ;
        RECT 2913.785 342.635 2913.955 342.805 ;
        RECT 5.665 337.195 5.835 337.365 ;
        RECT 6.125 337.195 6.295 337.365 ;
        RECT 6.585 337.195 6.755 337.365 ;
        RECT 2910.105 337.195 2910.275 337.365 ;
        RECT 2912.865 337.195 2913.035 337.365 ;
        RECT 2913.325 337.195 2913.495 337.365 ;
        RECT 2913.785 337.195 2913.955 337.365 ;
        RECT 5.665 331.755 5.835 331.925 ;
        RECT 6.125 331.755 6.295 331.925 ;
        RECT 6.585 331.755 6.755 331.925 ;
        RECT 2910.105 331.755 2910.275 331.925 ;
        RECT 2912.865 331.755 2913.035 331.925 ;
        RECT 2913.325 331.755 2913.495 331.925 ;
        RECT 2913.785 331.755 2913.955 331.925 ;
        RECT 5.665 326.315 5.835 326.485 ;
        RECT 6.125 326.315 6.295 326.485 ;
        RECT 6.585 326.315 6.755 326.485 ;
        RECT 2910.105 326.315 2910.275 326.485 ;
        RECT 2912.865 326.315 2913.035 326.485 ;
        RECT 2913.325 326.315 2913.495 326.485 ;
        RECT 2913.785 326.315 2913.955 326.485 ;
        RECT 5.665 320.875 5.835 321.045 ;
        RECT 6.125 320.875 6.295 321.045 ;
        RECT 6.585 320.875 6.755 321.045 ;
        RECT 2910.105 320.875 2910.275 321.045 ;
        RECT 2912.865 320.875 2913.035 321.045 ;
        RECT 2913.325 320.875 2913.495 321.045 ;
        RECT 2913.785 320.875 2913.955 321.045 ;
        RECT 5.665 315.435 5.835 315.605 ;
        RECT 6.125 315.435 6.295 315.605 ;
        RECT 6.585 315.435 6.755 315.605 ;
        RECT 8.885 315.435 9.055 315.605 ;
        RECT 9.345 315.435 9.515 315.605 ;
        RECT 9.805 315.435 9.975 315.605 ;
        RECT 2910.105 315.435 2910.275 315.605 ;
        RECT 2912.865 315.435 2913.035 315.605 ;
        RECT 2913.325 315.435 2913.495 315.605 ;
        RECT 2913.785 315.435 2913.955 315.605 ;
        RECT 5.665 309.995 5.835 310.165 ;
        RECT 6.125 309.995 6.295 310.165 ;
        RECT 6.585 309.995 6.755 310.165 ;
        RECT 2910.105 309.995 2910.275 310.165 ;
        RECT 2912.865 309.995 2913.035 310.165 ;
        RECT 2913.325 309.995 2913.495 310.165 ;
        RECT 2913.785 309.995 2913.955 310.165 ;
        RECT 5.665 304.555 5.835 304.725 ;
        RECT 6.125 304.555 6.295 304.725 ;
        RECT 6.585 304.555 6.755 304.725 ;
        RECT 2910.105 304.555 2910.275 304.725 ;
        RECT 2912.865 304.555 2913.035 304.725 ;
        RECT 2913.325 304.555 2913.495 304.725 ;
        RECT 2913.785 304.555 2913.955 304.725 ;
        RECT 5.665 299.115 5.835 299.285 ;
        RECT 6.125 299.115 6.295 299.285 ;
        RECT 6.585 299.115 6.755 299.285 ;
        RECT 2910.105 299.115 2910.275 299.285 ;
        RECT 2912.865 299.115 2913.035 299.285 ;
        RECT 2913.325 299.115 2913.495 299.285 ;
        RECT 2913.785 299.115 2913.955 299.285 ;
        RECT 5.665 293.675 5.835 293.845 ;
        RECT 6.125 293.675 6.295 293.845 ;
        RECT 6.585 293.675 6.755 293.845 ;
        RECT 2910.105 293.675 2910.275 293.845 ;
        RECT 2912.865 293.675 2913.035 293.845 ;
        RECT 2913.325 293.675 2913.495 293.845 ;
        RECT 2913.785 293.675 2913.955 293.845 ;
        RECT 5.665 288.235 5.835 288.405 ;
        RECT 6.125 288.235 6.295 288.405 ;
        RECT 6.585 288.235 6.755 288.405 ;
        RECT 2909.185 288.235 2909.355 288.405 ;
        RECT 2909.645 288.235 2909.815 288.405 ;
        RECT 2910.105 288.235 2910.275 288.405 ;
        RECT 2912.865 288.235 2913.035 288.405 ;
        RECT 2913.325 288.235 2913.495 288.405 ;
        RECT 2913.785 288.235 2913.955 288.405 ;
        RECT 5.665 282.795 5.835 282.965 ;
        RECT 6.125 282.795 6.295 282.965 ;
        RECT 6.585 282.795 6.755 282.965 ;
        RECT 2910.105 282.795 2910.275 282.965 ;
        RECT 2912.865 282.795 2913.035 282.965 ;
        RECT 2913.325 282.795 2913.495 282.965 ;
        RECT 2913.785 282.795 2913.955 282.965 ;
        RECT 5.665 277.355 5.835 277.525 ;
        RECT 6.125 277.355 6.295 277.525 ;
        RECT 6.585 277.355 6.755 277.525 ;
        RECT 2910.105 277.355 2910.275 277.525 ;
        RECT 2912.865 277.355 2913.035 277.525 ;
        RECT 2913.325 277.355 2913.495 277.525 ;
        RECT 2913.785 277.355 2913.955 277.525 ;
        RECT 5.665 271.915 5.835 272.085 ;
        RECT 6.125 271.915 6.295 272.085 ;
        RECT 6.585 271.915 6.755 272.085 ;
        RECT 2910.105 271.915 2910.275 272.085 ;
        RECT 2912.865 271.915 2913.035 272.085 ;
        RECT 2913.325 271.915 2913.495 272.085 ;
        RECT 2913.785 271.915 2913.955 272.085 ;
        RECT 5.665 266.475 5.835 266.645 ;
        RECT 6.125 266.475 6.295 266.645 ;
        RECT 6.585 266.475 6.755 266.645 ;
        RECT 2910.105 266.475 2910.275 266.645 ;
        RECT 2912.865 266.475 2913.035 266.645 ;
        RECT 2913.325 266.475 2913.495 266.645 ;
        RECT 2913.785 266.475 2913.955 266.645 ;
        RECT 5.665 261.035 5.835 261.205 ;
        RECT 6.125 261.035 6.295 261.205 ;
        RECT 6.585 261.035 6.755 261.205 ;
        RECT 2910.105 261.035 2910.275 261.205 ;
        RECT 2912.865 261.035 2913.035 261.205 ;
        RECT 2913.325 261.035 2913.495 261.205 ;
        RECT 2913.785 261.035 2913.955 261.205 ;
        RECT 5.665 255.595 5.835 255.765 ;
        RECT 6.125 255.595 6.295 255.765 ;
        RECT 6.585 255.595 6.755 255.765 ;
        RECT 2910.105 255.595 2910.275 255.765 ;
        RECT 2912.865 255.595 2913.035 255.765 ;
        RECT 2913.325 255.595 2913.495 255.765 ;
        RECT 2913.785 255.595 2913.955 255.765 ;
        RECT 5.665 250.155 5.835 250.325 ;
        RECT 6.125 250.155 6.295 250.325 ;
        RECT 6.585 250.155 6.755 250.325 ;
        RECT 2910.105 250.155 2910.275 250.325 ;
        RECT 2912.865 250.155 2913.035 250.325 ;
        RECT 2913.325 250.155 2913.495 250.325 ;
        RECT 2913.785 250.155 2913.955 250.325 ;
        RECT 5.665 244.715 5.835 244.885 ;
        RECT 6.125 244.715 6.295 244.885 ;
        RECT 6.585 244.715 6.755 244.885 ;
        RECT 2910.105 244.715 2910.275 244.885 ;
        RECT 2912.865 244.715 2913.035 244.885 ;
        RECT 2913.325 244.715 2913.495 244.885 ;
        RECT 2913.785 244.715 2913.955 244.885 ;
        RECT 5.665 239.275 5.835 239.445 ;
        RECT 6.125 239.275 6.295 239.445 ;
        RECT 6.585 239.275 6.755 239.445 ;
        RECT 2910.105 239.275 2910.275 239.445 ;
        RECT 2912.865 239.275 2913.035 239.445 ;
        RECT 2913.325 239.275 2913.495 239.445 ;
        RECT 2913.785 239.275 2913.955 239.445 ;
        RECT 5.665 233.835 5.835 234.005 ;
        RECT 6.125 233.835 6.295 234.005 ;
        RECT 6.585 233.835 6.755 234.005 ;
        RECT 2910.105 233.835 2910.275 234.005 ;
        RECT 2910.565 233.835 2910.735 234.005 ;
        RECT 2911.025 233.835 2911.195 234.005 ;
        RECT 2911.485 233.835 2911.655 234.005 ;
        RECT 2912.865 233.835 2913.035 234.005 ;
        RECT 2913.325 233.835 2913.495 234.005 ;
        RECT 2913.785 233.835 2913.955 234.005 ;
        RECT 5.665 228.395 5.835 228.565 ;
        RECT 6.125 228.395 6.295 228.565 ;
        RECT 6.585 228.395 6.755 228.565 ;
        RECT 2910.105 228.395 2910.275 228.565 ;
        RECT 2912.865 228.395 2913.035 228.565 ;
        RECT 2913.325 228.395 2913.495 228.565 ;
        RECT 2913.785 228.395 2913.955 228.565 ;
        RECT 5.665 222.955 5.835 223.125 ;
        RECT 6.125 222.955 6.295 223.125 ;
        RECT 6.585 222.955 6.755 223.125 ;
        RECT 2910.105 222.955 2910.275 223.125 ;
        RECT 2912.865 222.955 2913.035 223.125 ;
        RECT 2913.325 222.955 2913.495 223.125 ;
        RECT 2913.785 222.955 2913.955 223.125 ;
        RECT 5.665 217.515 5.835 217.685 ;
        RECT 6.125 217.515 6.295 217.685 ;
        RECT 6.585 217.515 6.755 217.685 ;
        RECT 2910.105 217.515 2910.275 217.685 ;
        RECT 2912.865 217.515 2913.035 217.685 ;
        RECT 2913.325 217.515 2913.495 217.685 ;
        RECT 2913.785 217.515 2913.955 217.685 ;
        RECT 5.665 212.075 5.835 212.245 ;
        RECT 6.125 212.075 6.295 212.245 ;
        RECT 6.585 212.075 6.755 212.245 ;
        RECT 2910.105 212.075 2910.275 212.245 ;
        RECT 2912.865 212.075 2913.035 212.245 ;
        RECT 2913.325 212.075 2913.495 212.245 ;
        RECT 2913.785 212.075 2913.955 212.245 ;
        RECT 5.665 206.635 5.835 206.805 ;
        RECT 6.125 206.635 6.295 206.805 ;
        RECT 6.585 206.635 6.755 206.805 ;
        RECT 2910.105 206.635 2910.275 206.805 ;
        RECT 2912.865 206.635 2913.035 206.805 ;
        RECT 2913.325 206.635 2913.495 206.805 ;
        RECT 2913.785 206.635 2913.955 206.805 ;
        RECT 5.665 201.195 5.835 201.365 ;
        RECT 6.125 201.195 6.295 201.365 ;
        RECT 6.585 201.195 6.755 201.365 ;
        RECT 2910.105 201.195 2910.275 201.365 ;
        RECT 2912.865 201.195 2913.035 201.365 ;
        RECT 2913.325 201.195 2913.495 201.365 ;
        RECT 2913.785 201.195 2913.955 201.365 ;
        RECT 5.665 195.755 5.835 195.925 ;
        RECT 6.125 195.755 6.295 195.925 ;
        RECT 6.585 195.755 6.755 195.925 ;
        RECT 2910.105 195.755 2910.275 195.925 ;
        RECT 2912.865 195.755 2913.035 195.925 ;
        RECT 2913.325 195.755 2913.495 195.925 ;
        RECT 2913.785 195.755 2913.955 195.925 ;
        RECT 5.665 190.315 5.835 190.485 ;
        RECT 6.125 190.315 6.295 190.485 ;
        RECT 6.585 190.315 6.755 190.485 ;
        RECT 2910.105 190.315 2910.275 190.485 ;
        RECT 2912.865 190.315 2913.035 190.485 ;
        RECT 2913.325 190.315 2913.495 190.485 ;
        RECT 2913.785 190.315 2913.955 190.485 ;
        RECT 5.665 184.875 5.835 185.045 ;
        RECT 6.125 184.875 6.295 185.045 ;
        RECT 6.585 184.875 6.755 185.045 ;
        RECT 2910.105 184.875 2910.275 185.045 ;
        RECT 2912.865 184.875 2913.035 185.045 ;
        RECT 2913.325 184.875 2913.495 185.045 ;
        RECT 2913.785 184.875 2913.955 185.045 ;
        RECT 5.665 179.435 5.835 179.605 ;
        RECT 6.125 179.435 6.295 179.605 ;
        RECT 6.585 179.435 6.755 179.605 ;
        RECT 2910.105 179.435 2910.275 179.605 ;
        RECT 2912.865 179.435 2913.035 179.605 ;
        RECT 2913.325 179.435 2913.495 179.605 ;
        RECT 2913.785 179.435 2913.955 179.605 ;
        RECT 5.665 173.995 5.835 174.165 ;
        RECT 6.125 173.995 6.295 174.165 ;
        RECT 6.585 173.995 6.755 174.165 ;
        RECT 2910.105 173.995 2910.275 174.165 ;
        RECT 2912.865 173.995 2913.035 174.165 ;
        RECT 2913.325 173.995 2913.495 174.165 ;
        RECT 2913.785 173.995 2913.955 174.165 ;
        RECT 5.665 168.555 5.835 168.725 ;
        RECT 6.125 168.555 6.295 168.725 ;
        RECT 6.585 168.555 6.755 168.725 ;
        RECT 2910.105 168.555 2910.275 168.725 ;
        RECT 2912.865 168.555 2913.035 168.725 ;
        RECT 2913.325 168.555 2913.495 168.725 ;
        RECT 2913.785 168.555 2913.955 168.725 ;
        RECT 5.665 163.115 5.835 163.285 ;
        RECT 6.125 163.115 6.295 163.285 ;
        RECT 6.585 163.115 6.755 163.285 ;
        RECT 2910.105 163.115 2910.275 163.285 ;
        RECT 2912.865 163.115 2913.035 163.285 ;
        RECT 2913.325 163.115 2913.495 163.285 ;
        RECT 2913.785 163.115 2913.955 163.285 ;
        RECT 5.665 157.675 5.835 157.845 ;
        RECT 6.125 157.675 6.295 157.845 ;
        RECT 6.585 157.675 6.755 157.845 ;
        RECT 2910.105 157.675 2910.275 157.845 ;
        RECT 2912.865 157.675 2913.035 157.845 ;
        RECT 2913.325 157.675 2913.495 157.845 ;
        RECT 2913.785 157.675 2913.955 157.845 ;
        RECT 5.665 152.235 5.835 152.405 ;
        RECT 6.125 152.235 6.295 152.405 ;
        RECT 6.585 152.235 6.755 152.405 ;
        RECT 2910.105 152.235 2910.275 152.405 ;
        RECT 2912.865 152.235 2913.035 152.405 ;
        RECT 2913.325 152.235 2913.495 152.405 ;
        RECT 2913.785 152.235 2913.955 152.405 ;
        RECT 5.665 146.795 5.835 146.965 ;
        RECT 6.125 146.795 6.295 146.965 ;
        RECT 6.585 146.795 6.755 146.965 ;
        RECT 2910.105 146.795 2910.275 146.965 ;
        RECT 2912.865 146.795 2913.035 146.965 ;
        RECT 2913.325 146.795 2913.495 146.965 ;
        RECT 2913.785 146.795 2913.955 146.965 ;
        RECT 5.665 141.355 5.835 141.525 ;
        RECT 6.125 141.355 6.295 141.525 ;
        RECT 6.585 141.355 6.755 141.525 ;
        RECT 2910.105 141.355 2910.275 141.525 ;
        RECT 2912.865 141.355 2913.035 141.525 ;
        RECT 2913.325 141.355 2913.495 141.525 ;
        RECT 2913.785 141.355 2913.955 141.525 ;
        RECT 5.665 135.915 5.835 136.085 ;
        RECT 6.125 135.915 6.295 136.085 ;
        RECT 6.585 135.915 6.755 136.085 ;
        RECT 2910.105 135.915 2910.275 136.085 ;
        RECT 2912.865 135.915 2913.035 136.085 ;
        RECT 2913.325 135.915 2913.495 136.085 ;
        RECT 2913.785 135.915 2913.955 136.085 ;
        RECT 5.665 130.475 5.835 130.645 ;
        RECT 6.125 130.475 6.295 130.645 ;
        RECT 6.585 130.475 6.755 130.645 ;
        RECT 2910.105 130.475 2910.275 130.645 ;
        RECT 2912.865 130.475 2913.035 130.645 ;
        RECT 2913.325 130.475 2913.495 130.645 ;
        RECT 2913.785 130.475 2913.955 130.645 ;
        RECT 5.665 125.035 5.835 125.205 ;
        RECT 6.125 125.035 6.295 125.205 ;
        RECT 6.585 125.035 6.755 125.205 ;
        RECT 7.045 125.035 7.215 125.205 ;
        RECT 7.505 125.035 7.675 125.205 ;
        RECT 7.965 125.035 8.135 125.205 ;
        RECT 8.425 125.035 8.595 125.205 ;
        RECT 8.885 125.035 9.055 125.205 ;
        RECT 9.345 125.035 9.515 125.205 ;
        RECT 9.805 125.035 9.975 125.205 ;
        RECT 10.265 125.035 10.435 125.205 ;
        RECT 10.725 125.035 10.895 125.205 ;
        RECT 11.185 125.035 11.355 125.205 ;
        RECT 11.645 125.035 11.815 125.205 ;
        RECT 12.105 125.035 12.275 125.205 ;
        RECT 12.565 125.035 12.735 125.205 ;
        RECT 13.025 125.035 13.195 125.205 ;
        RECT 13.485 125.035 13.655 125.205 ;
        RECT 2910.105 125.035 2910.275 125.205 ;
        RECT 2912.865 125.035 2913.035 125.205 ;
        RECT 2913.325 125.035 2913.495 125.205 ;
        RECT 2913.785 125.035 2913.955 125.205 ;
        RECT 5.665 119.595 5.835 119.765 ;
        RECT 6.125 119.595 6.295 119.765 ;
        RECT 6.585 119.595 6.755 119.765 ;
        RECT 2910.105 119.595 2910.275 119.765 ;
        RECT 2912.865 119.595 2913.035 119.765 ;
        RECT 2913.325 119.595 2913.495 119.765 ;
        RECT 2913.785 119.595 2913.955 119.765 ;
        RECT 5.665 114.155 5.835 114.325 ;
        RECT 6.125 114.155 6.295 114.325 ;
        RECT 6.585 114.155 6.755 114.325 ;
        RECT 2910.105 114.155 2910.275 114.325 ;
        RECT 2912.865 114.155 2913.035 114.325 ;
        RECT 2913.325 114.155 2913.495 114.325 ;
        RECT 2913.785 114.155 2913.955 114.325 ;
        RECT 5.665 108.715 5.835 108.885 ;
        RECT 6.125 108.715 6.295 108.885 ;
        RECT 6.585 108.715 6.755 108.885 ;
        RECT 2910.105 108.715 2910.275 108.885 ;
        RECT 2912.865 108.715 2913.035 108.885 ;
        RECT 2913.325 108.715 2913.495 108.885 ;
        RECT 2913.785 108.715 2913.955 108.885 ;
        RECT 5.665 103.275 5.835 103.445 ;
        RECT 6.125 103.275 6.295 103.445 ;
        RECT 6.585 103.275 6.755 103.445 ;
        RECT 8.885 103.275 9.055 103.445 ;
        RECT 9.345 103.275 9.515 103.445 ;
        RECT 9.805 103.275 9.975 103.445 ;
        RECT 2910.105 103.275 2910.275 103.445 ;
        RECT 2912.865 103.275 2913.035 103.445 ;
        RECT 2913.325 103.275 2913.495 103.445 ;
        RECT 2913.785 103.275 2913.955 103.445 ;
        RECT 5.665 97.835 5.835 98.005 ;
        RECT 6.125 97.835 6.295 98.005 ;
        RECT 6.585 97.835 6.755 98.005 ;
        RECT 2910.105 97.835 2910.275 98.005 ;
        RECT 2912.865 97.835 2913.035 98.005 ;
        RECT 2913.325 97.835 2913.495 98.005 ;
        RECT 2913.785 97.835 2913.955 98.005 ;
        RECT 5.665 92.395 5.835 92.565 ;
        RECT 6.125 92.395 6.295 92.565 ;
        RECT 6.585 92.395 6.755 92.565 ;
        RECT 2910.105 92.395 2910.275 92.565 ;
        RECT 2912.865 92.395 2913.035 92.565 ;
        RECT 2913.325 92.395 2913.495 92.565 ;
        RECT 2913.785 92.395 2913.955 92.565 ;
        RECT 5.665 86.955 5.835 87.125 ;
        RECT 6.125 86.955 6.295 87.125 ;
        RECT 6.585 86.955 6.755 87.125 ;
        RECT 2910.105 86.955 2910.275 87.125 ;
        RECT 2912.865 86.955 2913.035 87.125 ;
        RECT 2913.325 86.955 2913.495 87.125 ;
        RECT 2913.785 86.955 2913.955 87.125 ;
        RECT 5.665 81.515 5.835 81.685 ;
        RECT 6.125 81.515 6.295 81.685 ;
        RECT 6.585 81.515 6.755 81.685 ;
        RECT 2910.105 81.515 2910.275 81.685 ;
        RECT 2912.865 81.515 2913.035 81.685 ;
        RECT 2913.325 81.515 2913.495 81.685 ;
        RECT 2913.785 81.515 2913.955 81.685 ;
        RECT 5.665 76.075 5.835 76.245 ;
        RECT 6.125 76.075 6.295 76.245 ;
        RECT 6.585 76.075 6.755 76.245 ;
        RECT 2910.105 76.075 2910.275 76.245 ;
        RECT 2912.865 76.075 2913.035 76.245 ;
        RECT 2913.325 76.075 2913.495 76.245 ;
        RECT 2913.785 76.075 2913.955 76.245 ;
        RECT 5.665 70.635 5.835 70.805 ;
        RECT 6.125 70.635 6.295 70.805 ;
        RECT 6.585 70.635 6.755 70.805 ;
        RECT 2910.105 70.635 2910.275 70.805 ;
        RECT 2912.865 70.635 2913.035 70.805 ;
        RECT 2913.325 70.635 2913.495 70.805 ;
        RECT 2913.785 70.635 2913.955 70.805 ;
        RECT 5.665 65.195 5.835 65.365 ;
        RECT 6.125 65.195 6.295 65.365 ;
        RECT 6.585 65.195 6.755 65.365 ;
        RECT 2910.105 65.195 2910.275 65.365 ;
        RECT 2912.865 65.195 2913.035 65.365 ;
        RECT 2913.325 65.195 2913.495 65.365 ;
        RECT 2913.785 65.195 2913.955 65.365 ;
        RECT 5.665 59.755 5.835 59.925 ;
        RECT 6.125 59.755 6.295 59.925 ;
        RECT 6.585 59.755 6.755 59.925 ;
        RECT 2909.185 59.755 2909.355 59.925 ;
        RECT 2909.645 59.755 2909.815 59.925 ;
        RECT 2910.105 59.755 2910.275 59.925 ;
        RECT 2912.865 59.755 2913.035 59.925 ;
        RECT 2913.325 59.755 2913.495 59.925 ;
        RECT 2913.785 59.755 2913.955 59.925 ;
        RECT 5.665 54.315 5.835 54.485 ;
        RECT 6.125 54.315 6.295 54.485 ;
        RECT 6.585 54.315 6.755 54.485 ;
        RECT 2910.105 54.315 2910.275 54.485 ;
        RECT 2912.865 54.315 2913.035 54.485 ;
        RECT 2913.325 54.315 2913.495 54.485 ;
        RECT 2913.785 54.315 2913.955 54.485 ;
        RECT 5.665 48.875 5.835 49.045 ;
        RECT 6.125 48.875 6.295 49.045 ;
        RECT 6.585 48.875 6.755 49.045 ;
        RECT 2910.105 48.875 2910.275 49.045 ;
        RECT 2912.865 48.875 2913.035 49.045 ;
        RECT 2913.325 48.875 2913.495 49.045 ;
        RECT 2913.785 48.875 2913.955 49.045 ;
        RECT 5.665 43.435 5.835 43.605 ;
        RECT 6.125 43.435 6.295 43.605 ;
        RECT 6.585 43.435 6.755 43.605 ;
        RECT 7.045 43.435 7.215 43.605 ;
        RECT 7.505 43.435 7.675 43.605 ;
        RECT 7.965 43.435 8.135 43.605 ;
        RECT 8.425 43.435 8.595 43.605 ;
        RECT 8.885 43.435 9.055 43.605 ;
        RECT 9.345 43.435 9.515 43.605 ;
        RECT 9.805 43.435 9.975 43.605 ;
        RECT 10.265 43.435 10.435 43.605 ;
        RECT 10.725 43.435 10.895 43.605 ;
        RECT 11.185 43.435 11.355 43.605 ;
        RECT 11.645 43.435 11.815 43.605 ;
        RECT 12.105 43.435 12.275 43.605 ;
        RECT 12.565 43.435 12.735 43.605 ;
        RECT 13.025 43.435 13.195 43.605 ;
        RECT 13.485 43.435 13.655 43.605 ;
        RECT 2910.105 43.435 2910.275 43.605 ;
        RECT 2912.865 43.435 2913.035 43.605 ;
        RECT 2913.325 43.435 2913.495 43.605 ;
        RECT 2913.785 43.435 2913.955 43.605 ;
        RECT 5.665 37.995 5.835 38.165 ;
        RECT 6.125 37.995 6.295 38.165 ;
        RECT 6.585 37.995 6.755 38.165 ;
        RECT 2910.105 37.995 2910.275 38.165 ;
        RECT 2912.865 37.995 2913.035 38.165 ;
        RECT 2913.325 37.995 2913.495 38.165 ;
        RECT 2913.785 37.995 2913.955 38.165 ;
        RECT 5.665 32.555 5.835 32.725 ;
        RECT 6.125 32.555 6.295 32.725 ;
        RECT 6.585 32.555 6.755 32.725 ;
        RECT 2910.105 32.555 2910.275 32.725 ;
        RECT 2912.865 32.555 2913.035 32.725 ;
        RECT 2913.325 32.555 2913.495 32.725 ;
        RECT 2913.785 32.555 2913.955 32.725 ;
        RECT 5.665 27.115 5.835 27.285 ;
        RECT 6.125 27.115 6.295 27.285 ;
        RECT 6.585 27.115 6.755 27.285 ;
        RECT 2910.105 27.115 2910.275 27.285 ;
        RECT 2912.865 27.115 2913.035 27.285 ;
        RECT 2913.325 27.115 2913.495 27.285 ;
        RECT 2913.785 27.115 2913.955 27.285 ;
        RECT 5.665 21.675 5.835 21.845 ;
        RECT 6.125 21.675 6.295 21.845 ;
        RECT 6.585 21.675 6.755 21.845 ;
        RECT 7.045 21.675 7.215 21.845 ;
        RECT 7.505 21.675 7.675 21.845 ;
        RECT 7.965 21.675 8.135 21.845 ;
        RECT 8.425 21.675 8.595 21.845 ;
        RECT 8.885 21.675 9.055 21.845 ;
        RECT 9.345 21.675 9.515 21.845 ;
        RECT 9.805 21.675 9.975 21.845 ;
        RECT 10.265 21.675 10.435 21.845 ;
        RECT 10.725 21.675 10.895 21.845 ;
        RECT 11.185 21.675 11.355 21.845 ;
        RECT 11.645 21.675 11.815 21.845 ;
        RECT 12.105 21.675 12.275 21.845 ;
        RECT 12.565 21.675 12.735 21.845 ;
        RECT 13.025 21.675 13.195 21.845 ;
        RECT 13.485 21.675 13.655 21.845 ;
        RECT 2910.105 21.675 2910.275 21.845 ;
        RECT 2912.865 21.675 2913.035 21.845 ;
        RECT 2913.325 21.675 2913.495 21.845 ;
        RECT 2913.785 21.675 2913.955 21.845 ;
        RECT 5.665 16.235 5.835 16.405 ;
        RECT 6.125 16.235 6.295 16.405 ;
        RECT 6.585 16.235 6.755 16.405 ;
        RECT 7.045 16.235 7.215 16.405 ;
        RECT 7.505 16.235 7.675 16.405 ;
        RECT 7.965 16.235 8.135 16.405 ;
        RECT 8.425 16.235 8.595 16.405 ;
        RECT 8.885 16.235 9.055 16.405 ;
        RECT 9.345 16.235 9.515 16.405 ;
        RECT 9.805 16.235 9.975 16.405 ;
        RECT 10.265 16.235 10.435 16.405 ;
        RECT 10.725 16.235 10.895 16.405 ;
        RECT 11.185 16.235 11.355 16.405 ;
        RECT 11.645 16.235 11.815 16.405 ;
        RECT 12.105 16.235 12.275 16.405 ;
        RECT 12.565 16.235 12.735 16.405 ;
        RECT 13.025 16.235 13.195 16.405 ;
        RECT 13.485 16.235 13.655 16.405 ;
        RECT 2907.345 16.235 2907.515 16.405 ;
        RECT 2907.805 16.235 2907.975 16.405 ;
        RECT 2908.265 16.235 2908.435 16.405 ;
        RECT 2908.725 16.235 2908.895 16.405 ;
        RECT 2909.185 16.235 2909.355 16.405 ;
        RECT 2909.645 16.235 2909.815 16.405 ;
        RECT 2910.105 16.235 2910.275 16.405 ;
        RECT 2910.565 16.235 2910.735 16.405 ;
        RECT 2911.025 16.235 2911.195 16.405 ;
        RECT 2911.485 16.235 2911.655 16.405 ;
        RECT 2912.865 16.235 2913.035 16.405 ;
        RECT 2913.325 16.235 2913.495 16.405 ;
        RECT 2913.785 16.235 2913.955 16.405 ;
        RECT 5.665 10.795 5.835 10.965 ;
        RECT 6.125 10.795 6.295 10.965 ;
        RECT 6.585 10.795 6.755 10.965 ;
        RECT 8.885 10.795 9.055 10.965 ;
        RECT 9.345 10.795 9.515 10.965 ;
        RECT 9.805 10.795 9.975 10.965 ;
        RECT 10.265 10.795 10.435 10.965 ;
        RECT 10.725 10.795 10.895 10.965 ;
        RECT 11.185 10.795 11.355 10.965 ;
        RECT 19.925 10.795 20.095 10.965 ;
        RECT 34.185 10.795 34.355 10.965 ;
        RECT 48.445 10.795 48.615 10.965 ;
        RECT 62.705 10.795 62.875 10.965 ;
        RECT 76.965 10.795 77.135 10.965 ;
        RECT 82.025 10.795 82.195 10.965 ;
        RECT 82.485 10.795 82.655 10.965 ;
        RECT 82.945 10.795 83.115 10.965 ;
        RECT 83.405 10.795 83.575 10.965 ;
        RECT 83.865 10.795 84.035 10.965 ;
        RECT 84.325 10.795 84.495 10.965 ;
        RECT 84.785 10.795 84.955 10.965 ;
        RECT 85.245 10.795 85.415 10.965 ;
        RECT 85.705 10.795 85.875 10.965 ;
        RECT 86.165 10.795 86.335 10.965 ;
        RECT 86.625 10.795 86.795 10.965 ;
        RECT 87.085 10.795 87.255 10.965 ;
        RECT 87.545 10.795 87.715 10.965 ;
        RECT 88.005 10.795 88.175 10.965 ;
        RECT 88.465 10.795 88.635 10.965 ;
        RECT 88.925 10.795 89.095 10.965 ;
        RECT 89.385 10.795 89.555 10.965 ;
        RECT 89.845 10.795 90.015 10.965 ;
        RECT 90.305 10.795 90.475 10.965 ;
        RECT 91.225 10.795 91.395 10.965 ;
        RECT 105.485 10.795 105.655 10.965 ;
        RECT 119.745 10.795 119.915 10.965 ;
        RECT 134.005 10.795 134.175 10.965 ;
        RECT 148.265 10.795 148.435 10.965 ;
        RECT 162.525 10.795 162.695 10.965 ;
        RECT 176.785 10.795 176.955 10.965 ;
        RECT 191.045 10.795 191.215 10.965 ;
        RECT 205.305 10.795 205.475 10.965 ;
        RECT 205.765 10.795 205.935 10.965 ;
        RECT 206.225 10.795 206.395 10.965 ;
        RECT 206.685 10.795 206.855 10.965 ;
        RECT 207.145 10.795 207.315 10.965 ;
        RECT 207.605 10.795 207.775 10.965 ;
        RECT 208.065 10.795 208.235 10.965 ;
        RECT 208.525 10.795 208.695 10.965 ;
        RECT 208.985 10.795 209.155 10.965 ;
        RECT 209.445 10.795 209.615 10.965 ;
        RECT 209.905 10.795 210.075 10.965 ;
        RECT 210.365 10.795 210.535 10.965 ;
        RECT 210.825 10.795 210.995 10.965 ;
        RECT 211.285 10.795 211.455 10.965 ;
        RECT 211.745 10.795 211.915 10.965 ;
        RECT 212.205 10.795 212.375 10.965 ;
        RECT 212.665 10.795 212.835 10.965 ;
        RECT 219.565 10.795 219.735 10.965 ;
        RECT 225.545 10.795 225.715 10.965 ;
        RECT 226.005 10.795 226.175 10.965 ;
        RECT 226.465 10.795 226.635 10.965 ;
        RECT 226.925 10.795 227.095 10.965 ;
        RECT 227.385 10.795 227.555 10.965 ;
        RECT 227.845 10.795 228.015 10.965 ;
        RECT 228.305 10.795 228.475 10.965 ;
        RECT 228.765 10.795 228.935 10.965 ;
        RECT 229.225 10.795 229.395 10.965 ;
        RECT 229.685 10.795 229.855 10.965 ;
        RECT 230.145 10.795 230.315 10.965 ;
        RECT 230.605 10.795 230.775 10.965 ;
        RECT 231.065 10.795 231.235 10.965 ;
        RECT 231.525 10.795 231.695 10.965 ;
        RECT 233.825 10.795 233.995 10.965 ;
        RECT 240.265 10.795 240.435 10.965 ;
        RECT 240.725 10.795 240.895 10.965 ;
        RECT 241.185 10.795 241.355 10.965 ;
        RECT 241.645 10.795 241.815 10.965 ;
        RECT 242.105 10.795 242.275 10.965 ;
        RECT 242.565 10.795 242.735 10.965 ;
        RECT 243.025 10.795 243.195 10.965 ;
        RECT 243.485 10.795 243.655 10.965 ;
        RECT 243.945 10.795 244.115 10.965 ;
        RECT 248.085 10.795 248.255 10.965 ;
        RECT 262.345 10.795 262.515 10.965 ;
        RECT 262.805 10.795 262.975 10.965 ;
        RECT 263.265 10.795 263.435 10.965 ;
        RECT 263.725 10.795 263.895 10.965 ;
        RECT 264.185 10.795 264.355 10.965 ;
        RECT 264.645 10.795 264.815 10.965 ;
        RECT 265.105 10.795 265.275 10.965 ;
        RECT 265.565 10.795 265.735 10.965 ;
        RECT 266.025 10.795 266.195 10.965 ;
        RECT 266.485 10.795 266.655 10.965 ;
        RECT 266.945 10.795 267.115 10.965 ;
        RECT 267.405 10.795 267.575 10.965 ;
        RECT 267.865 10.795 268.035 10.965 ;
        RECT 268.325 10.795 268.495 10.965 ;
        RECT 268.785 10.795 268.955 10.965 ;
        RECT 276.605 10.795 276.775 10.965 ;
        RECT 290.865 10.795 291.035 10.965 ;
        RECT 305.125 10.795 305.295 10.965 ;
        RECT 319.385 10.795 319.555 10.965 ;
        RECT 333.645 10.795 333.815 10.965 ;
        RECT 347.905 10.795 348.075 10.965 ;
        RECT 352.505 10.795 352.675 10.965 ;
        RECT 352.965 10.795 353.135 10.965 ;
        RECT 353.425 10.795 353.595 10.965 ;
        RECT 362.165 10.795 362.335 10.965 ;
        RECT 376.425 10.795 376.595 10.965 ;
        RECT 390.685 10.795 390.855 10.965 ;
        RECT 391.145 10.795 391.315 10.965 ;
        RECT 391.605 10.795 391.775 10.965 ;
        RECT 392.065 10.795 392.235 10.965 ;
        RECT 392.525 10.795 392.695 10.965 ;
        RECT 392.985 10.795 393.155 10.965 ;
        RECT 393.445 10.795 393.615 10.965 ;
        RECT 393.905 10.795 394.075 10.965 ;
        RECT 394.365 10.795 394.535 10.965 ;
        RECT 394.825 10.795 394.995 10.965 ;
        RECT 395.285 10.795 395.455 10.965 ;
        RECT 395.745 10.795 395.915 10.965 ;
        RECT 396.205 10.795 396.375 10.965 ;
        RECT 396.665 10.795 396.835 10.965 ;
        RECT 397.125 10.795 397.295 10.965 ;
        RECT 397.585 10.795 397.755 10.965 ;
        RECT 398.045 10.795 398.215 10.965 ;
        RECT 398.505 10.795 398.675 10.965 ;
        RECT 398.965 10.795 399.135 10.965 ;
        RECT 399.425 10.795 399.595 10.965 ;
        RECT 399.885 10.795 400.055 10.965 ;
        RECT 400.345 10.795 400.515 10.965 ;
        RECT 400.805 10.795 400.975 10.965 ;
        RECT 404.945 10.795 405.115 10.965 ;
        RECT 419.205 10.795 419.375 10.965 ;
        RECT 433.465 10.795 433.635 10.965 ;
        RECT 447.725 10.795 447.895 10.965 ;
        RECT 450.945 10.795 451.115 10.965 ;
        RECT 451.405 10.795 451.575 10.965 ;
        RECT 451.865 10.795 452.035 10.965 ;
        RECT 452.325 10.795 452.495 10.965 ;
        RECT 452.785 10.795 452.955 10.965 ;
        RECT 453.245 10.795 453.415 10.965 ;
        RECT 453.705 10.795 453.875 10.965 ;
        RECT 454.165 10.795 454.335 10.965 ;
        RECT 454.625 10.795 454.795 10.965 ;
        RECT 455.085 10.795 455.255 10.965 ;
        RECT 455.545 10.795 455.715 10.965 ;
        RECT 456.005 10.795 456.175 10.965 ;
        RECT 456.465 10.795 456.635 10.965 ;
        RECT 456.925 10.795 457.095 10.965 ;
        RECT 461.985 10.795 462.155 10.965 ;
        RECT 476.245 10.795 476.415 10.965 ;
        RECT 490.505 10.795 490.675 10.965 ;
        RECT 504.765 10.795 504.935 10.965 ;
        RECT 519.025 10.795 519.195 10.965 ;
        RECT 533.285 10.795 533.455 10.965 ;
        RECT 547.545 10.795 547.715 10.965 ;
        RECT 561.805 10.795 561.975 10.965 ;
        RECT 576.065 10.795 576.235 10.965 ;
        RECT 590.325 10.795 590.495 10.965 ;
        RECT 604.585 10.795 604.755 10.965 ;
        RECT 618.845 10.795 619.015 10.965 ;
        RECT 633.105 10.795 633.275 10.965 ;
        RECT 647.365 10.795 647.535 10.965 ;
        RECT 661.625 10.795 661.795 10.965 ;
        RECT 675.885 10.795 676.055 10.965 ;
        RECT 690.145 10.795 690.315 10.965 ;
        RECT 704.405 10.795 704.575 10.965 ;
        RECT 718.665 10.795 718.835 10.965 ;
        RECT 732.925 10.795 733.095 10.965 ;
        RECT 747.185 10.795 747.355 10.965 ;
        RECT 761.445 10.795 761.615 10.965 ;
        RECT 775.705 10.795 775.875 10.965 ;
        RECT 789.965 10.795 790.135 10.965 ;
        RECT 804.225 10.795 804.395 10.965 ;
        RECT 818.485 10.795 818.655 10.965 ;
        RECT 832.745 10.795 832.915 10.965 ;
        RECT 847.005 10.795 847.175 10.965 ;
        RECT 861.265 10.795 861.435 10.965 ;
        RECT 875.525 10.795 875.695 10.965 ;
        RECT 889.785 10.795 889.955 10.965 ;
        RECT 904.045 10.795 904.215 10.965 ;
        RECT 918.305 10.795 918.475 10.965 ;
        RECT 932.565 10.795 932.735 10.965 ;
        RECT 946.825 10.795 946.995 10.965 ;
        RECT 961.085 10.795 961.255 10.965 ;
        RECT 975.345 10.795 975.515 10.965 ;
        RECT 989.605 10.795 989.775 10.965 ;
        RECT 1003.865 10.795 1004.035 10.965 ;
        RECT 1018.125 10.795 1018.295 10.965 ;
        RECT 1032.385 10.795 1032.555 10.965 ;
        RECT 1046.645 10.795 1046.815 10.965 ;
        RECT 1060.905 10.795 1061.075 10.965 ;
        RECT 1075.165 10.795 1075.335 10.965 ;
        RECT 1089.425 10.795 1089.595 10.965 ;
        RECT 1103.685 10.795 1103.855 10.965 ;
        RECT 1117.945 10.795 1118.115 10.965 ;
        RECT 1132.205 10.795 1132.375 10.965 ;
        RECT 1146.465 10.795 1146.635 10.965 ;
        RECT 1160.725 10.795 1160.895 10.965 ;
        RECT 1174.985 10.795 1175.155 10.965 ;
        RECT 1189.245 10.795 1189.415 10.965 ;
        RECT 1203.505 10.795 1203.675 10.965 ;
        RECT 1217.765 10.795 1217.935 10.965 ;
        RECT 1232.025 10.795 1232.195 10.965 ;
        RECT 1246.285 10.795 1246.455 10.965 ;
        RECT 1260.545 10.795 1260.715 10.965 ;
        RECT 1274.805 10.795 1274.975 10.965 ;
        RECT 1289.065 10.795 1289.235 10.965 ;
        RECT 1303.325 10.795 1303.495 10.965 ;
        RECT 1317.585 10.795 1317.755 10.965 ;
        RECT 1331.845 10.795 1332.015 10.965 ;
        RECT 1346.105 10.795 1346.275 10.965 ;
        RECT 1360.365 10.795 1360.535 10.965 ;
        RECT 1374.625 10.795 1374.795 10.965 ;
        RECT 1388.885 10.795 1389.055 10.965 ;
        RECT 1403.145 10.795 1403.315 10.965 ;
        RECT 1417.405 10.795 1417.575 10.965 ;
        RECT 1431.665 10.795 1431.835 10.965 ;
        RECT 1445.925 10.795 1446.095 10.965 ;
        RECT 1460.185 10.795 1460.355 10.965 ;
        RECT 1474.445 10.795 1474.615 10.965 ;
        RECT 1488.705 10.795 1488.875 10.965 ;
        RECT 1502.965 10.795 1503.135 10.965 ;
        RECT 1517.225 10.795 1517.395 10.965 ;
        RECT 1531.485 10.795 1531.655 10.965 ;
        RECT 1545.745 10.795 1545.915 10.965 ;
        RECT 1560.005 10.795 1560.175 10.965 ;
        RECT 1574.265 10.795 1574.435 10.965 ;
        RECT 1588.525 10.795 1588.695 10.965 ;
        RECT 1602.785 10.795 1602.955 10.965 ;
        RECT 1617.045 10.795 1617.215 10.965 ;
        RECT 1631.305 10.795 1631.475 10.965 ;
        RECT 1645.565 10.795 1645.735 10.965 ;
        RECT 1659.825 10.795 1659.995 10.965 ;
        RECT 1674.085 10.795 1674.255 10.965 ;
        RECT 1688.345 10.795 1688.515 10.965 ;
        RECT 1702.605 10.795 1702.775 10.965 ;
        RECT 1716.865 10.795 1717.035 10.965 ;
        RECT 1731.125 10.795 1731.295 10.965 ;
        RECT 1745.385 10.795 1745.555 10.965 ;
        RECT 1759.645 10.795 1759.815 10.965 ;
        RECT 1773.905 10.795 1774.075 10.965 ;
        RECT 1788.165 10.795 1788.335 10.965 ;
        RECT 1802.425 10.795 1802.595 10.965 ;
        RECT 1816.685 10.795 1816.855 10.965 ;
        RECT 1830.945 10.795 1831.115 10.965 ;
        RECT 1845.205 10.795 1845.375 10.965 ;
        RECT 1859.465 10.795 1859.635 10.965 ;
        RECT 1873.725 10.795 1873.895 10.965 ;
        RECT 1887.985 10.795 1888.155 10.965 ;
        RECT 1902.245 10.795 1902.415 10.965 ;
        RECT 1916.505 10.795 1916.675 10.965 ;
        RECT 1930.765 10.795 1930.935 10.965 ;
        RECT 1945.025 10.795 1945.195 10.965 ;
        RECT 1959.285 10.795 1959.455 10.965 ;
        RECT 1973.545 10.795 1973.715 10.965 ;
        RECT 1987.805 10.795 1987.975 10.965 ;
        RECT 2002.065 10.795 2002.235 10.965 ;
        RECT 2016.325 10.795 2016.495 10.965 ;
        RECT 2030.585 10.795 2030.755 10.965 ;
        RECT 2044.845 10.795 2045.015 10.965 ;
        RECT 2059.105 10.795 2059.275 10.965 ;
        RECT 2073.365 10.795 2073.535 10.965 ;
        RECT 2087.625 10.795 2087.795 10.965 ;
        RECT 2101.885 10.795 2102.055 10.965 ;
        RECT 2116.145 10.795 2116.315 10.965 ;
        RECT 2130.405 10.795 2130.575 10.965 ;
        RECT 2144.665 10.795 2144.835 10.965 ;
        RECT 2158.925 10.795 2159.095 10.965 ;
        RECT 2173.185 10.795 2173.355 10.965 ;
        RECT 2187.445 10.795 2187.615 10.965 ;
        RECT 2201.705 10.795 2201.875 10.965 ;
        RECT 2215.965 10.795 2216.135 10.965 ;
        RECT 2230.225 10.795 2230.395 10.965 ;
        RECT 2244.485 10.795 2244.655 10.965 ;
        RECT 2258.745 10.795 2258.915 10.965 ;
        RECT 2273.005 10.795 2273.175 10.965 ;
        RECT 2287.265 10.795 2287.435 10.965 ;
        RECT 2301.525 10.795 2301.695 10.965 ;
        RECT 2315.785 10.795 2315.955 10.965 ;
        RECT 2330.045 10.795 2330.215 10.965 ;
        RECT 2344.305 10.795 2344.475 10.965 ;
        RECT 2358.565 10.795 2358.735 10.965 ;
        RECT 2372.825 10.795 2372.995 10.965 ;
        RECT 2387.085 10.795 2387.255 10.965 ;
        RECT 2401.345 10.795 2401.515 10.965 ;
        RECT 2415.605 10.795 2415.775 10.965 ;
        RECT 2429.865 10.795 2430.035 10.965 ;
        RECT 2444.125 10.795 2444.295 10.965 ;
        RECT 2458.385 10.795 2458.555 10.965 ;
        RECT 2472.645 10.795 2472.815 10.965 ;
        RECT 2486.905 10.795 2487.075 10.965 ;
        RECT 2501.165 10.795 2501.335 10.965 ;
        RECT 2515.425 10.795 2515.595 10.965 ;
        RECT 2529.685 10.795 2529.855 10.965 ;
        RECT 2543.945 10.795 2544.115 10.965 ;
        RECT 2558.205 10.795 2558.375 10.965 ;
        RECT 2572.465 10.795 2572.635 10.965 ;
        RECT 2586.725 10.795 2586.895 10.965 ;
        RECT 2600.985 10.795 2601.155 10.965 ;
        RECT 2615.245 10.795 2615.415 10.965 ;
        RECT 2629.505 10.795 2629.675 10.965 ;
        RECT 2643.765 10.795 2643.935 10.965 ;
        RECT 2658.025 10.795 2658.195 10.965 ;
        RECT 2672.285 10.795 2672.455 10.965 ;
        RECT 2686.545 10.795 2686.715 10.965 ;
        RECT 2700.805 10.795 2700.975 10.965 ;
        RECT 2715.065 10.795 2715.235 10.965 ;
        RECT 2729.325 10.795 2729.495 10.965 ;
        RECT 2743.585 10.795 2743.755 10.965 ;
        RECT 2757.845 10.795 2758.015 10.965 ;
        RECT 2772.105 10.795 2772.275 10.965 ;
        RECT 2786.365 10.795 2786.535 10.965 ;
        RECT 2800.625 10.795 2800.795 10.965 ;
        RECT 2814.885 10.795 2815.055 10.965 ;
        RECT 2829.145 10.795 2829.315 10.965 ;
        RECT 2843.405 10.795 2843.575 10.965 ;
        RECT 2857.665 10.795 2857.835 10.965 ;
        RECT 2871.925 10.795 2872.095 10.965 ;
        RECT 2886.185 10.795 2886.355 10.965 ;
        RECT 2900.445 10.795 2900.615 10.965 ;
        RECT 2909.185 10.795 2909.355 10.965 ;
        RECT 2909.645 10.795 2909.815 10.965 ;
        RECT 2910.105 10.795 2910.275 10.965 ;
        RECT 2912.865 10.795 2913.035 10.965 ;
        RECT 2913.325 10.795 2913.495 10.965 ;
        RECT 2913.785 10.795 2913.955 10.965 ;
      LAYER met1 ;
        RECT 5.520 3508.560 2914.100 3509.040 ;
        RECT 5.520 3503.120 13.700 3503.600 ;
        RECT 2906.300 3503.120 2914.100 3503.600 ;
        RECT 5.520 3497.680 13.700 3498.160 ;
        RECT 2906.300 3497.680 2914.100 3498.160 ;
        RECT 5.520 3492.240 13.700 3492.720 ;
        RECT 2906.300 3492.240 2914.100 3492.720 ;
        RECT 5.520 3486.800 13.700 3487.280 ;
        RECT 2906.300 3486.800 2914.100 3487.280 ;
        RECT 5.520 3481.360 13.700 3481.840 ;
        RECT 2906.300 3481.360 2914.100 3481.840 ;
        RECT 5.520 3475.920 13.700 3476.400 ;
        RECT 2906.300 3475.920 2914.100 3476.400 ;
        RECT 5.520 3470.480 13.700 3470.960 ;
        RECT 2906.300 3470.480 2914.100 3470.960 ;
        RECT 5.520 3465.040 13.700 3465.520 ;
        RECT 2906.300 3465.040 2914.100 3465.520 ;
        RECT 5.520 3459.600 13.700 3460.080 ;
        RECT 2906.300 3459.600 2914.100 3460.080 ;
        RECT 5.520 3454.160 13.700 3454.640 ;
        RECT 2906.300 3454.160 2914.100 3454.640 ;
        RECT 5.520 3448.720 13.700 3449.200 ;
        RECT 2906.300 3448.720 2914.100 3449.200 ;
        RECT 5.520 3443.280 13.700 3443.760 ;
        RECT 2906.300 3443.280 2914.100 3443.760 ;
        RECT 5.520 3437.840 13.700 3438.320 ;
        RECT 2906.300 3437.840 2914.100 3438.320 ;
        RECT 5.520 3432.400 13.700 3432.880 ;
        RECT 2906.300 3432.400 2914.100 3432.880 ;
        RECT 5.520 3426.960 13.700 3427.440 ;
        RECT 2906.300 3426.960 2914.100 3427.440 ;
        RECT 5.520 3421.520 13.700 3422.000 ;
        RECT 2906.300 3421.520 2914.100 3422.000 ;
        RECT 5.520 3416.080 13.700 3416.560 ;
        RECT 2906.300 3416.080 2914.100 3416.560 ;
        RECT 5.520 3410.640 13.700 3411.120 ;
        RECT 2906.300 3410.640 2914.100 3411.120 ;
        RECT 5.520 3405.200 13.700 3405.680 ;
        RECT 2906.300 3405.200 2914.100 3405.680 ;
        RECT 5.520 3399.760 13.700 3400.240 ;
        RECT 2906.300 3399.760 2914.100 3400.240 ;
        RECT 5.520 3394.320 13.700 3394.800 ;
        RECT 2906.300 3394.320 2914.100 3394.800 ;
        RECT 5.520 3388.880 13.700 3389.360 ;
        RECT 2906.300 3388.880 2914.100 3389.360 ;
        RECT 5.520 3383.440 13.700 3383.920 ;
        RECT 2906.300 3383.440 2914.100 3383.920 ;
        RECT 5.520 3378.000 13.700 3378.480 ;
        RECT 2906.300 3378.000 2914.100 3378.480 ;
        RECT 5.520 3372.560 13.700 3373.040 ;
        RECT 2906.300 3372.560 2914.100 3373.040 ;
        RECT 5.520 3367.120 13.700 3367.600 ;
        RECT 2906.300 3367.120 2914.100 3367.600 ;
        RECT 5.520 3361.680 13.700 3362.160 ;
        RECT 2906.300 3361.680 2914.100 3362.160 ;
        RECT 5.520 3356.240 13.700 3356.720 ;
        RECT 2906.300 3356.240 2914.100 3356.720 ;
        RECT 5.520 3350.800 13.700 3351.280 ;
        RECT 2906.300 3350.800 2914.100 3351.280 ;
        RECT 5.520 3345.360 13.700 3345.840 ;
        RECT 2906.300 3345.360 2914.100 3345.840 ;
        RECT 5.520 3339.920 13.700 3340.400 ;
        RECT 2906.300 3339.920 2914.100 3340.400 ;
        RECT 5.520 3334.480 13.700 3334.960 ;
        RECT 2906.300 3334.480 2914.100 3334.960 ;
        RECT 5.520 3329.040 13.700 3329.520 ;
        RECT 2906.300 3329.040 2914.100 3329.520 ;
        RECT 5.520 3323.600 13.700 3324.080 ;
        RECT 2906.300 3323.600 2914.100 3324.080 ;
        RECT 5.520 3318.160 13.700 3318.640 ;
        RECT 2906.300 3318.160 2914.100 3318.640 ;
        RECT 5.520 3312.720 13.700 3313.200 ;
        RECT 2906.300 3312.720 2914.100 3313.200 ;
        RECT 5.520 3307.280 13.700 3307.760 ;
        RECT 2906.300 3307.280 2914.100 3307.760 ;
        RECT 5.520 3301.840 13.700 3302.320 ;
        RECT 2906.300 3301.840 2914.100 3302.320 ;
        RECT 5.520 3296.400 13.700 3296.880 ;
        RECT 2906.300 3296.400 2914.100 3296.880 ;
        RECT 5.520 3290.960 13.700 3291.440 ;
        RECT 2906.300 3290.960 2914.100 3291.440 ;
        RECT 5.520 3285.520 13.700 3286.000 ;
        RECT 2906.300 3285.520 2914.100 3286.000 ;
        RECT 5.520 3280.080 13.700 3280.560 ;
        RECT 2906.300 3280.080 2914.100 3280.560 ;
        RECT 5.520 3274.640 13.700 3275.120 ;
        RECT 2906.300 3274.640 2914.100 3275.120 ;
        RECT 5.520 3269.200 13.700 3269.680 ;
        RECT 2906.300 3269.200 2914.100 3269.680 ;
        RECT 5.520 3263.760 13.700 3264.240 ;
        RECT 2906.300 3263.760 2914.100 3264.240 ;
        RECT 5.520 3258.320 13.700 3258.800 ;
        RECT 2906.300 3258.320 2914.100 3258.800 ;
        RECT 5.520 3252.880 13.700 3253.360 ;
        RECT 2906.300 3252.880 2914.100 3253.360 ;
        RECT 5.520 3247.440 13.700 3247.920 ;
        RECT 2906.300 3247.440 2914.100 3247.920 ;
        RECT 5.520 3242.000 13.700 3242.480 ;
        RECT 2906.300 3242.000 2914.100 3242.480 ;
        RECT 5.520 3236.560 13.700 3237.040 ;
        RECT 2906.300 3236.560 2914.100 3237.040 ;
        RECT 5.520 3231.120 13.700 3231.600 ;
        RECT 2906.300 3231.120 2914.100 3231.600 ;
        RECT 5.520 3225.680 13.700 3226.160 ;
        RECT 2906.300 3225.680 2914.100 3226.160 ;
        RECT 5.520 3220.240 13.700 3220.720 ;
        RECT 2906.300 3220.240 2914.100 3220.720 ;
        RECT 5.520 3214.800 13.700 3215.280 ;
        RECT 2906.300 3214.800 2914.100 3215.280 ;
        RECT 5.520 3209.360 13.700 3209.840 ;
        RECT 2906.300 3209.360 2914.100 3209.840 ;
        RECT 5.520 3203.920 13.700 3204.400 ;
        RECT 2906.300 3203.920 2914.100 3204.400 ;
        RECT 5.520 3198.480 13.700 3198.960 ;
        RECT 2906.300 3198.480 2914.100 3198.960 ;
        RECT 5.520 3193.040 13.700 3193.520 ;
        RECT 2906.300 3193.040 2914.100 3193.520 ;
        RECT 5.520 3187.600 13.700 3188.080 ;
        RECT 2906.300 3187.600 2914.100 3188.080 ;
        RECT 5.520 3182.160 13.700 3182.640 ;
        RECT 2906.300 3182.160 2914.100 3182.640 ;
        RECT 5.520 3176.720 13.700 3177.200 ;
        RECT 2906.300 3176.720 2914.100 3177.200 ;
        RECT 5.520 3171.280 13.700 3171.760 ;
        RECT 2906.300 3171.280 2914.100 3171.760 ;
        RECT 5.520 3165.840 13.700 3166.320 ;
        RECT 2906.300 3165.840 2914.100 3166.320 ;
        RECT 5.520 3160.400 13.700 3160.880 ;
        RECT 2906.300 3160.400 2914.100 3160.880 ;
        RECT 5.520 3154.960 13.700 3155.440 ;
        RECT 2906.300 3154.960 2914.100 3155.440 ;
        RECT 5.520 3149.520 13.700 3150.000 ;
        RECT 2906.300 3149.520 2914.100 3150.000 ;
        RECT 5.520 3144.080 13.700 3144.560 ;
        RECT 2906.300 3144.080 2914.100 3144.560 ;
        RECT 5.520 3138.640 13.700 3139.120 ;
        RECT 2906.300 3138.640 2914.100 3139.120 ;
        RECT 5.520 3133.200 13.700 3133.680 ;
        RECT 2906.300 3133.200 2914.100 3133.680 ;
        RECT 5.520 3127.760 13.700 3128.240 ;
        RECT 2906.300 3127.760 2914.100 3128.240 ;
        RECT 5.520 3122.320 13.700 3122.800 ;
        RECT 2906.300 3122.320 2914.100 3122.800 ;
        RECT 5.520 3116.880 13.700 3117.360 ;
        RECT 2906.300 3116.880 2914.100 3117.360 ;
        RECT 5.520 3111.440 13.700 3111.920 ;
        RECT 2906.300 3111.440 2914.100 3111.920 ;
        RECT 5.520 3106.000 13.700 3106.480 ;
        RECT 2906.300 3106.000 2914.100 3106.480 ;
        RECT 5.520 3100.560 13.700 3101.040 ;
        RECT 2906.300 3100.560 2914.100 3101.040 ;
        RECT 5.520 3095.120 13.700 3095.600 ;
        RECT 2906.300 3095.120 2914.100 3095.600 ;
        RECT 5.520 3089.680 13.700 3090.160 ;
        RECT 2906.300 3089.680 2914.100 3090.160 ;
        RECT 5.520 3084.240 13.700 3084.720 ;
        RECT 2906.300 3084.240 2914.100 3084.720 ;
        RECT 5.520 3078.800 13.700 3079.280 ;
        RECT 2906.300 3078.800 2914.100 3079.280 ;
        RECT 5.520 3073.360 13.700 3073.840 ;
        RECT 2906.300 3073.360 2914.100 3073.840 ;
        RECT 5.520 3067.920 13.700 3068.400 ;
        RECT 2906.300 3067.920 2914.100 3068.400 ;
        RECT 5.520 3062.480 13.700 3062.960 ;
        RECT 2906.300 3062.480 2914.100 3062.960 ;
        RECT 5.520 3057.040 13.700 3057.520 ;
        RECT 2906.300 3057.040 2914.100 3057.520 ;
        RECT 5.520 3051.600 13.700 3052.080 ;
        RECT 2906.300 3051.600 2914.100 3052.080 ;
        RECT 5.520 3046.160 13.700 3046.640 ;
        RECT 2906.300 3046.160 2914.100 3046.640 ;
        RECT 5.520 3040.720 13.700 3041.200 ;
        RECT 2906.300 3040.720 2914.100 3041.200 ;
        RECT 5.520 3035.280 13.700 3035.760 ;
        RECT 2906.300 3035.280 2914.100 3035.760 ;
        RECT 5.520 3029.840 13.700 3030.320 ;
        RECT 2906.300 3029.840 2914.100 3030.320 ;
        RECT 5.520 3024.400 13.700 3024.880 ;
        RECT 2906.300 3024.400 2914.100 3024.880 ;
        RECT 5.520 3018.960 13.700 3019.440 ;
        RECT 2906.300 3018.960 2914.100 3019.440 ;
        RECT 5.520 3013.520 13.700 3014.000 ;
        RECT 2906.300 3013.520 2914.100 3014.000 ;
        RECT 5.520 3008.080 13.700 3008.560 ;
        RECT 2906.300 3008.080 2914.100 3008.560 ;
        RECT 5.520 3002.640 13.700 3003.120 ;
        RECT 2906.300 3002.640 2914.100 3003.120 ;
        RECT 5.520 2997.200 13.700 2997.680 ;
        RECT 2906.300 2997.200 2914.100 2997.680 ;
        RECT 5.520 2991.760 13.700 2992.240 ;
        RECT 2906.300 2991.760 2914.100 2992.240 ;
        RECT 5.520 2986.320 13.700 2986.800 ;
        RECT 2906.300 2986.320 2914.100 2986.800 ;
        RECT 5.520 2980.880 13.700 2981.360 ;
        RECT 2906.300 2980.880 2914.100 2981.360 ;
        RECT 5.520 2975.440 13.700 2975.920 ;
        RECT 2906.300 2975.440 2914.100 2975.920 ;
        RECT 5.520 2970.000 13.700 2970.480 ;
        RECT 2906.300 2970.000 2914.100 2970.480 ;
        RECT 5.520 2964.560 13.700 2965.040 ;
        RECT 2906.300 2964.560 2914.100 2965.040 ;
        RECT 5.520 2959.120 13.700 2959.600 ;
        RECT 2906.300 2959.120 2914.100 2959.600 ;
        RECT 5.520 2953.680 13.700 2954.160 ;
        RECT 2906.300 2953.680 2914.100 2954.160 ;
        RECT 5.520 2948.240 13.700 2948.720 ;
        RECT 2906.300 2948.240 2914.100 2948.720 ;
        RECT 5.520 2942.800 13.700 2943.280 ;
        RECT 2906.300 2942.800 2914.100 2943.280 ;
        RECT 5.520 2937.360 13.700 2937.840 ;
        RECT 2906.300 2937.360 2914.100 2937.840 ;
        RECT 5.520 2931.920 13.700 2932.400 ;
        RECT 2906.300 2931.920 2914.100 2932.400 ;
        RECT 5.520 2926.480 13.700 2926.960 ;
        RECT 2906.300 2926.480 2914.100 2926.960 ;
        RECT 5.520 2921.040 13.700 2921.520 ;
        RECT 2906.300 2921.040 2914.100 2921.520 ;
        RECT 5.520 2915.600 13.700 2916.080 ;
        RECT 2906.300 2915.600 2914.100 2916.080 ;
        RECT 5.520 2910.160 13.700 2910.640 ;
        RECT 2906.300 2910.160 2914.100 2910.640 ;
        RECT 5.520 2904.720 13.700 2905.200 ;
        RECT 2906.300 2904.720 2914.100 2905.200 ;
        RECT 5.520 2899.280 13.700 2899.760 ;
        RECT 2906.300 2899.280 2914.100 2899.760 ;
        RECT 5.520 2893.840 13.700 2894.320 ;
        RECT 2906.300 2893.840 2914.100 2894.320 ;
        RECT 5.520 2888.400 13.700 2888.880 ;
        RECT 2906.300 2888.400 2914.100 2888.880 ;
        RECT 5.520 2882.960 13.700 2883.440 ;
        RECT 2906.300 2882.960 2914.100 2883.440 ;
        RECT 5.520 2877.520 13.700 2878.000 ;
        RECT 2906.300 2877.520 2914.100 2878.000 ;
        RECT 5.520 2872.080 13.700 2872.560 ;
        RECT 2906.300 2872.080 2914.100 2872.560 ;
        RECT 5.520 2866.640 13.700 2867.120 ;
        RECT 2906.300 2866.640 2914.100 2867.120 ;
        RECT 5.520 2861.200 13.700 2861.680 ;
        RECT 2906.300 2861.200 2914.100 2861.680 ;
        RECT 5.520 2855.760 13.700 2856.240 ;
        RECT 2906.300 2855.760 2914.100 2856.240 ;
        RECT 5.520 2850.320 13.700 2850.800 ;
        RECT 2906.300 2850.320 2914.100 2850.800 ;
        RECT 5.520 2844.880 13.700 2845.360 ;
        RECT 2906.300 2844.880 2914.100 2845.360 ;
        RECT 5.520 2839.440 13.700 2839.920 ;
        RECT 2906.300 2839.440 2914.100 2839.920 ;
        RECT 5.520 2834.000 13.700 2834.480 ;
        RECT 2906.300 2834.000 2914.100 2834.480 ;
        RECT 5.520 2828.560 13.700 2829.040 ;
        RECT 2906.300 2828.560 2914.100 2829.040 ;
        RECT 5.520 2823.120 13.700 2823.600 ;
        RECT 2906.300 2823.120 2914.100 2823.600 ;
        RECT 5.520 2817.680 13.700 2818.160 ;
        RECT 2906.300 2817.680 2914.100 2818.160 ;
        RECT 5.520 2812.240 13.700 2812.720 ;
        RECT 2906.300 2812.240 2914.100 2812.720 ;
        RECT 5.520 2806.800 13.700 2807.280 ;
        RECT 2906.300 2806.800 2914.100 2807.280 ;
        RECT 5.520 2801.360 13.700 2801.840 ;
        RECT 2906.300 2801.360 2914.100 2801.840 ;
        RECT 5.520 2795.920 13.700 2796.400 ;
        RECT 2906.300 2795.920 2914.100 2796.400 ;
        RECT 5.520 2790.480 13.700 2790.960 ;
        RECT 2906.300 2790.480 2914.100 2790.960 ;
        RECT 5.520 2785.040 13.700 2785.520 ;
        RECT 2906.300 2785.040 2914.100 2785.520 ;
        RECT 5.520 2779.600 13.700 2780.080 ;
        RECT 2906.300 2779.600 2914.100 2780.080 ;
        RECT 5.520 2774.160 13.700 2774.640 ;
        RECT 2906.300 2774.160 2914.100 2774.640 ;
        RECT 5.520 2768.720 13.700 2769.200 ;
        RECT 2906.300 2768.720 2914.100 2769.200 ;
        RECT 5.520 2763.280 13.700 2763.760 ;
        RECT 2906.300 2763.280 2914.100 2763.760 ;
        RECT 5.520 2757.840 13.700 2758.320 ;
        RECT 2906.300 2757.840 2914.100 2758.320 ;
        RECT 5.520 2752.400 13.700 2752.880 ;
        RECT 2906.300 2752.400 2914.100 2752.880 ;
        RECT 5.520 2746.960 13.700 2747.440 ;
        RECT 2906.300 2746.960 2914.100 2747.440 ;
        RECT 5.520 2741.520 13.700 2742.000 ;
        RECT 2906.300 2741.520 2914.100 2742.000 ;
        RECT 5.520 2736.080 13.700 2736.560 ;
        RECT 2906.300 2736.080 2914.100 2736.560 ;
        RECT 5.520 2730.640 13.700 2731.120 ;
        RECT 2906.300 2730.640 2914.100 2731.120 ;
        RECT 5.520 2725.200 13.700 2725.680 ;
        RECT 2906.300 2725.200 2914.100 2725.680 ;
        RECT 5.520 2719.760 13.700 2720.240 ;
        RECT 2906.300 2719.760 2914.100 2720.240 ;
        RECT 5.520 2714.320 13.700 2714.800 ;
        RECT 2906.300 2714.320 2914.100 2714.800 ;
        RECT 5.520 2708.880 13.700 2709.360 ;
        RECT 2906.300 2708.880 2914.100 2709.360 ;
        RECT 5.520 2703.440 13.700 2703.920 ;
        RECT 2906.300 2703.440 2914.100 2703.920 ;
        RECT 5.520 2698.000 13.700 2698.480 ;
        RECT 2906.300 2698.000 2914.100 2698.480 ;
        RECT 5.520 2692.560 13.700 2693.040 ;
        RECT 2906.300 2692.560 2914.100 2693.040 ;
        RECT 5.520 2687.120 13.700 2687.600 ;
        RECT 2906.300 2687.120 2914.100 2687.600 ;
        RECT 5.520 2681.680 13.700 2682.160 ;
        RECT 2906.300 2681.680 2914.100 2682.160 ;
        RECT 5.520 2676.240 13.700 2676.720 ;
        RECT 2906.300 2676.240 2914.100 2676.720 ;
        RECT 5.520 2670.800 13.700 2671.280 ;
        RECT 2906.300 2670.800 2914.100 2671.280 ;
        RECT 5.520 2665.360 13.700 2665.840 ;
        RECT 2906.300 2665.360 2914.100 2665.840 ;
        RECT 5.520 2659.920 13.700 2660.400 ;
        RECT 2906.300 2659.920 2914.100 2660.400 ;
        RECT 5.520 2654.480 13.700 2654.960 ;
        RECT 2906.300 2654.480 2914.100 2654.960 ;
        RECT 5.520 2649.040 13.700 2649.520 ;
        RECT 2906.300 2649.040 2914.100 2649.520 ;
        RECT 5.520 2643.600 13.700 2644.080 ;
        RECT 2906.300 2643.600 2914.100 2644.080 ;
        RECT 5.520 2638.160 13.700 2638.640 ;
        RECT 2906.300 2638.160 2914.100 2638.640 ;
        RECT 5.520 2632.720 13.700 2633.200 ;
        RECT 2906.300 2632.720 2914.100 2633.200 ;
        RECT 5.520 2627.280 13.700 2627.760 ;
        RECT 2906.300 2627.280 2914.100 2627.760 ;
        RECT 5.520 2621.840 13.700 2622.320 ;
        RECT 2906.300 2621.840 2914.100 2622.320 ;
        RECT 5.520 2616.400 13.700 2616.880 ;
        RECT 2906.300 2616.400 2914.100 2616.880 ;
        RECT 5.520 2610.960 13.700 2611.440 ;
        RECT 2906.300 2610.960 2914.100 2611.440 ;
        RECT 5.520 2605.520 13.700 2606.000 ;
        RECT 2906.300 2605.520 2914.100 2606.000 ;
        RECT 5.520 2600.080 13.700 2600.560 ;
        RECT 2906.300 2600.080 2914.100 2600.560 ;
        RECT 5.520 2594.640 13.700 2595.120 ;
        RECT 2906.300 2594.640 2914.100 2595.120 ;
        RECT 5.520 2589.200 13.700 2589.680 ;
        RECT 2906.300 2589.200 2914.100 2589.680 ;
        RECT 5.520 2583.760 13.700 2584.240 ;
        RECT 2906.300 2583.760 2914.100 2584.240 ;
        RECT 5.520 2578.320 13.700 2578.800 ;
        RECT 2906.300 2578.320 2914.100 2578.800 ;
        RECT 5.520 2572.880 13.700 2573.360 ;
        RECT 2906.300 2572.880 2914.100 2573.360 ;
        RECT 5.520 2567.440 13.700 2567.920 ;
        RECT 2906.300 2567.440 2914.100 2567.920 ;
        RECT 5.520 2562.000 13.700 2562.480 ;
        RECT 2906.300 2562.000 2914.100 2562.480 ;
        RECT 5.520 2556.560 13.700 2557.040 ;
        RECT 2906.300 2556.560 2914.100 2557.040 ;
        RECT 5.520 2551.120 13.700 2551.600 ;
        RECT 2906.300 2551.120 2914.100 2551.600 ;
        RECT 5.520 2545.680 13.700 2546.160 ;
        RECT 2906.300 2545.680 2914.100 2546.160 ;
        RECT 5.520 2540.240 13.700 2540.720 ;
        RECT 2906.300 2540.240 2914.100 2540.720 ;
        RECT 5.520 2534.800 13.700 2535.280 ;
        RECT 2906.300 2534.800 2914.100 2535.280 ;
        RECT 5.520 2529.360 13.700 2529.840 ;
        RECT 2906.300 2529.360 2914.100 2529.840 ;
        RECT 5.520 2523.920 13.700 2524.400 ;
        RECT 2906.300 2523.920 2914.100 2524.400 ;
        RECT 5.520 2518.480 13.700 2518.960 ;
        RECT 2906.300 2518.480 2914.100 2518.960 ;
        RECT 5.520 2513.040 13.700 2513.520 ;
        RECT 2906.300 2513.040 2914.100 2513.520 ;
        RECT 5.520 2507.600 13.700 2508.080 ;
        RECT 2906.300 2507.600 2914.100 2508.080 ;
        RECT 5.520 2502.160 13.700 2502.640 ;
        RECT 2906.300 2502.160 2914.100 2502.640 ;
        RECT 5.520 2496.720 13.700 2497.200 ;
        RECT 2906.300 2496.720 2914.100 2497.200 ;
        RECT 5.520 2491.280 13.700 2491.760 ;
        RECT 2906.300 2491.280 2914.100 2491.760 ;
        RECT 5.520 2485.840 13.700 2486.320 ;
        RECT 2906.300 2485.840 2914.100 2486.320 ;
        RECT 5.520 2480.400 13.700 2480.880 ;
        RECT 2906.300 2480.400 2914.100 2480.880 ;
        RECT 5.520 2474.960 13.700 2475.440 ;
        RECT 2906.300 2474.960 2914.100 2475.440 ;
        RECT 5.520 2469.520 13.700 2470.000 ;
        RECT 2906.300 2469.520 2914.100 2470.000 ;
        RECT 5.520 2464.080 13.700 2464.560 ;
        RECT 2906.300 2464.080 2914.100 2464.560 ;
        RECT 5.520 2458.640 13.700 2459.120 ;
        RECT 2906.300 2458.640 2914.100 2459.120 ;
        RECT 5.520 2453.200 13.700 2453.680 ;
        RECT 2906.300 2453.200 2914.100 2453.680 ;
        RECT 5.520 2447.760 13.700 2448.240 ;
        RECT 2906.300 2447.760 2914.100 2448.240 ;
        RECT 5.520 2442.320 13.700 2442.800 ;
        RECT 2906.300 2442.320 2914.100 2442.800 ;
        RECT 5.520 2436.880 13.700 2437.360 ;
        RECT 2906.300 2436.880 2914.100 2437.360 ;
        RECT 5.520 2431.440 13.700 2431.920 ;
        RECT 2906.300 2431.440 2914.100 2431.920 ;
        RECT 5.520 2426.000 13.700 2426.480 ;
        RECT 2906.300 2426.000 2914.100 2426.480 ;
        RECT 5.520 2420.560 13.700 2421.040 ;
        RECT 2906.300 2420.560 2914.100 2421.040 ;
        RECT 5.520 2415.120 13.700 2415.600 ;
        RECT 2906.300 2415.120 2914.100 2415.600 ;
        RECT 5.520 2409.680 13.700 2410.160 ;
        RECT 2906.300 2409.680 2914.100 2410.160 ;
        RECT 5.520 2404.240 13.700 2404.720 ;
        RECT 2906.300 2404.240 2914.100 2404.720 ;
        RECT 5.520 2398.800 13.700 2399.280 ;
        RECT 2906.300 2398.800 2914.100 2399.280 ;
        RECT 5.520 2393.360 13.700 2393.840 ;
        RECT 2906.300 2393.360 2914.100 2393.840 ;
        RECT 5.520 2387.920 13.700 2388.400 ;
        RECT 2906.300 2387.920 2914.100 2388.400 ;
        RECT 5.520 2382.480 13.700 2382.960 ;
        RECT 2906.300 2382.480 2914.100 2382.960 ;
        RECT 5.520 2377.040 13.700 2377.520 ;
        RECT 2906.300 2377.040 2914.100 2377.520 ;
        RECT 5.520 2371.600 13.700 2372.080 ;
        RECT 2906.300 2371.600 2914.100 2372.080 ;
        RECT 5.520 2366.160 13.700 2366.640 ;
        RECT 2906.300 2366.160 2914.100 2366.640 ;
        RECT 5.520 2360.720 13.700 2361.200 ;
        RECT 2906.300 2360.720 2914.100 2361.200 ;
        RECT 5.520 2355.280 13.700 2355.760 ;
        RECT 2906.300 2355.280 2914.100 2355.760 ;
        RECT 5.520 2349.840 13.700 2350.320 ;
        RECT 2906.300 2349.840 2914.100 2350.320 ;
        RECT 5.520 2344.400 13.700 2344.880 ;
        RECT 2906.300 2344.400 2914.100 2344.880 ;
        RECT 5.520 2338.960 13.700 2339.440 ;
        RECT 2906.300 2338.960 2914.100 2339.440 ;
        RECT 5.520 2333.520 13.700 2334.000 ;
        RECT 2906.300 2333.520 2914.100 2334.000 ;
        RECT 5.520 2328.080 13.700 2328.560 ;
        RECT 2906.300 2328.080 2914.100 2328.560 ;
        RECT 5.520 2322.640 13.700 2323.120 ;
        RECT 2906.300 2322.640 2914.100 2323.120 ;
        RECT 5.520 2317.200 13.700 2317.680 ;
        RECT 2906.300 2317.200 2914.100 2317.680 ;
        RECT 5.520 2311.760 13.700 2312.240 ;
        RECT 2906.300 2311.760 2914.100 2312.240 ;
        RECT 5.520 2306.320 13.700 2306.800 ;
        RECT 2906.300 2306.320 2914.100 2306.800 ;
        RECT 5.520 2300.880 13.700 2301.360 ;
        RECT 2906.300 2300.880 2914.100 2301.360 ;
        RECT 5.520 2295.440 13.700 2295.920 ;
        RECT 2906.300 2295.440 2914.100 2295.920 ;
        RECT 5.520 2290.000 13.700 2290.480 ;
        RECT 2906.300 2290.000 2914.100 2290.480 ;
        RECT 5.520 2284.560 13.700 2285.040 ;
        RECT 2906.300 2284.560 2914.100 2285.040 ;
        RECT 5.520 2279.120 13.700 2279.600 ;
        RECT 2906.300 2279.120 2914.100 2279.600 ;
        RECT 5.520 2273.680 13.700 2274.160 ;
        RECT 2906.300 2273.680 2914.100 2274.160 ;
        RECT 5.520 2268.240 13.700 2268.720 ;
        RECT 2906.300 2268.240 2914.100 2268.720 ;
        RECT 5.520 2262.800 13.700 2263.280 ;
        RECT 2906.300 2262.800 2914.100 2263.280 ;
        RECT 5.520 2257.360 13.700 2257.840 ;
        RECT 2906.300 2257.360 2914.100 2257.840 ;
        RECT 5.520 2251.920 13.700 2252.400 ;
        RECT 2906.300 2251.920 2914.100 2252.400 ;
        RECT 5.520 2246.480 13.700 2246.960 ;
        RECT 2906.300 2246.480 2914.100 2246.960 ;
        RECT 5.520 2241.040 13.700 2241.520 ;
        RECT 2906.300 2241.040 2914.100 2241.520 ;
        RECT 5.520 2235.600 13.700 2236.080 ;
        RECT 2906.300 2235.600 2914.100 2236.080 ;
        RECT 5.520 2230.160 13.700 2230.640 ;
        RECT 2906.300 2230.160 2914.100 2230.640 ;
        RECT 5.520 2224.720 13.700 2225.200 ;
        RECT 2906.300 2224.720 2914.100 2225.200 ;
        RECT 5.520 2219.280 13.700 2219.760 ;
        RECT 2906.300 2219.280 2914.100 2219.760 ;
        RECT 5.520 2213.840 13.700 2214.320 ;
        RECT 2906.300 2213.840 2914.100 2214.320 ;
        RECT 5.520 2208.400 13.700 2208.880 ;
        RECT 2906.300 2208.400 2914.100 2208.880 ;
        RECT 5.520 2202.960 13.700 2203.440 ;
        RECT 2906.300 2202.960 2914.100 2203.440 ;
        RECT 5.520 2197.520 13.700 2198.000 ;
        RECT 2906.300 2197.520 2914.100 2198.000 ;
        RECT 5.520 2192.080 13.700 2192.560 ;
        RECT 2906.300 2192.080 2914.100 2192.560 ;
        RECT 5.520 2186.640 13.700 2187.120 ;
        RECT 2906.300 2186.640 2914.100 2187.120 ;
        RECT 5.520 2181.200 13.700 2181.680 ;
        RECT 2906.300 2181.200 2914.100 2181.680 ;
        RECT 5.520 2175.760 13.700 2176.240 ;
        RECT 2906.300 2175.760 2914.100 2176.240 ;
        RECT 5.520 2170.320 13.700 2170.800 ;
        RECT 2906.300 2170.320 2914.100 2170.800 ;
        RECT 5.520 2164.880 13.700 2165.360 ;
        RECT 2906.300 2164.880 2914.100 2165.360 ;
        RECT 5.520 2159.440 13.700 2159.920 ;
        RECT 2906.300 2159.440 2914.100 2159.920 ;
        RECT 5.520 2154.000 13.700 2154.480 ;
        RECT 2906.300 2154.000 2914.100 2154.480 ;
        RECT 5.520 2148.560 13.700 2149.040 ;
        RECT 2906.300 2148.560 2914.100 2149.040 ;
        RECT 5.520 2143.120 13.700 2143.600 ;
        RECT 2906.300 2143.120 2914.100 2143.600 ;
        RECT 5.520 2137.680 13.700 2138.160 ;
        RECT 2906.300 2137.680 2914.100 2138.160 ;
        RECT 5.520 2132.240 13.700 2132.720 ;
        RECT 2906.300 2132.240 2914.100 2132.720 ;
        RECT 5.520 2126.800 13.700 2127.280 ;
        RECT 2906.300 2126.800 2914.100 2127.280 ;
        RECT 5.520 2121.360 13.700 2121.840 ;
        RECT 2906.300 2121.360 2914.100 2121.840 ;
        RECT 5.520 2115.920 13.700 2116.400 ;
        RECT 2906.300 2115.920 2914.100 2116.400 ;
        RECT 5.520 2110.480 13.700 2110.960 ;
        RECT 2906.300 2110.480 2914.100 2110.960 ;
        RECT 5.520 2105.040 13.700 2105.520 ;
        RECT 2906.300 2105.040 2914.100 2105.520 ;
        RECT 5.520 2099.600 13.700 2100.080 ;
        RECT 2906.300 2099.600 2914.100 2100.080 ;
        RECT 5.520 2094.160 13.700 2094.640 ;
        RECT 2906.300 2094.160 2914.100 2094.640 ;
        RECT 5.520 2088.720 13.700 2089.200 ;
        RECT 2906.300 2088.720 2914.100 2089.200 ;
        RECT 5.520 2083.280 13.700 2083.760 ;
        RECT 2906.300 2083.280 2914.100 2083.760 ;
        RECT 5.520 2077.840 13.700 2078.320 ;
        RECT 2906.300 2077.840 2914.100 2078.320 ;
        RECT 5.520 2072.400 13.700 2072.880 ;
        RECT 2906.300 2072.400 2914.100 2072.880 ;
        RECT 5.520 2066.960 13.700 2067.440 ;
        RECT 2906.300 2066.960 2914.100 2067.440 ;
        RECT 5.520 2061.520 13.700 2062.000 ;
        RECT 2906.300 2061.520 2914.100 2062.000 ;
        RECT 5.520 2056.080 13.700 2056.560 ;
        RECT 2906.300 2056.080 2914.100 2056.560 ;
        RECT 5.520 2050.640 13.700 2051.120 ;
        RECT 2906.300 2050.640 2914.100 2051.120 ;
        RECT 5.520 2045.200 13.700 2045.680 ;
        RECT 2906.300 2045.200 2914.100 2045.680 ;
        RECT 5.520 2039.760 13.700 2040.240 ;
        RECT 2906.300 2039.760 2914.100 2040.240 ;
        RECT 5.520 2034.320 13.700 2034.800 ;
        RECT 2906.300 2034.320 2914.100 2034.800 ;
        RECT 5.520 2028.880 13.700 2029.360 ;
        RECT 2906.300 2028.880 2914.100 2029.360 ;
        RECT 5.520 2023.440 13.700 2023.920 ;
        RECT 2906.300 2023.440 2914.100 2023.920 ;
        RECT 5.520 2018.000 13.700 2018.480 ;
        RECT 2906.300 2018.000 2914.100 2018.480 ;
        RECT 5.520 2012.560 13.700 2013.040 ;
        RECT 2906.300 2012.560 2914.100 2013.040 ;
        RECT 5.520 2007.120 13.700 2007.600 ;
        RECT 2906.300 2007.120 2914.100 2007.600 ;
        RECT 5.520 2001.680 13.700 2002.160 ;
        RECT 2906.300 2001.680 2914.100 2002.160 ;
        RECT 5.520 1996.240 13.700 1996.720 ;
        RECT 2906.300 1996.240 2914.100 1996.720 ;
        RECT 5.520 1990.800 13.700 1991.280 ;
        RECT 2906.300 1990.800 2914.100 1991.280 ;
        RECT 5.520 1985.360 13.700 1985.840 ;
        RECT 2906.300 1985.360 2914.100 1985.840 ;
        RECT 5.520 1979.920 13.700 1980.400 ;
        RECT 2906.300 1979.920 2914.100 1980.400 ;
        RECT 5.520 1974.480 13.700 1974.960 ;
        RECT 2906.300 1974.480 2914.100 1974.960 ;
        RECT 5.520 1969.040 13.700 1969.520 ;
        RECT 2906.300 1969.040 2914.100 1969.520 ;
        RECT 5.520 1963.600 13.700 1964.080 ;
        RECT 2906.300 1963.600 2914.100 1964.080 ;
        RECT 5.520 1958.160 13.700 1958.640 ;
        RECT 2906.300 1958.160 2914.100 1958.640 ;
        RECT 5.520 1952.720 13.700 1953.200 ;
        RECT 2906.300 1952.720 2914.100 1953.200 ;
        RECT 5.520 1947.280 13.700 1947.760 ;
        RECT 2906.300 1947.280 2914.100 1947.760 ;
        RECT 5.520 1941.840 13.700 1942.320 ;
        RECT 2906.300 1941.840 2914.100 1942.320 ;
        RECT 5.520 1936.400 13.700 1936.880 ;
        RECT 2906.300 1936.400 2914.100 1936.880 ;
        RECT 5.520 1930.960 13.700 1931.440 ;
        RECT 2906.300 1930.960 2914.100 1931.440 ;
        RECT 5.520 1925.520 13.700 1926.000 ;
        RECT 2906.300 1925.520 2914.100 1926.000 ;
        RECT 5.520 1920.080 13.700 1920.560 ;
        RECT 2906.300 1920.080 2914.100 1920.560 ;
        RECT 5.520 1914.640 13.700 1915.120 ;
        RECT 2906.300 1914.640 2914.100 1915.120 ;
        RECT 5.520 1909.200 13.700 1909.680 ;
        RECT 2906.300 1909.200 2914.100 1909.680 ;
        RECT 5.520 1903.760 13.700 1904.240 ;
        RECT 2906.300 1903.760 2914.100 1904.240 ;
        RECT 5.520 1898.320 13.700 1898.800 ;
        RECT 2906.300 1898.320 2914.100 1898.800 ;
        RECT 5.520 1892.880 13.700 1893.360 ;
        RECT 2906.300 1892.880 2914.100 1893.360 ;
        RECT 5.520 1887.440 13.700 1887.920 ;
        RECT 2906.300 1887.440 2914.100 1887.920 ;
        RECT 5.520 1882.000 13.700 1882.480 ;
        RECT 2906.300 1882.000 2914.100 1882.480 ;
        RECT 5.520 1876.560 13.700 1877.040 ;
        RECT 2906.300 1876.560 2914.100 1877.040 ;
        RECT 5.520 1871.120 13.700 1871.600 ;
        RECT 2906.300 1871.120 2914.100 1871.600 ;
        RECT 5.520 1865.680 13.700 1866.160 ;
        RECT 2906.300 1865.680 2914.100 1866.160 ;
        RECT 5.520 1860.240 13.700 1860.720 ;
        RECT 2906.300 1860.240 2914.100 1860.720 ;
        RECT 5.520 1854.800 13.700 1855.280 ;
        RECT 2906.300 1854.800 2914.100 1855.280 ;
        RECT 5.520 1849.360 13.700 1849.840 ;
        RECT 2906.300 1849.360 2914.100 1849.840 ;
        RECT 5.520 1843.920 13.700 1844.400 ;
        RECT 2906.300 1843.920 2914.100 1844.400 ;
        RECT 5.520 1838.480 13.700 1838.960 ;
        RECT 2906.300 1838.480 2914.100 1838.960 ;
        RECT 5.520 1833.040 13.700 1833.520 ;
        RECT 2906.300 1833.040 2914.100 1833.520 ;
        RECT 5.520 1827.600 13.700 1828.080 ;
        RECT 2906.300 1827.600 2914.100 1828.080 ;
        RECT 5.520 1822.160 13.700 1822.640 ;
        RECT 2906.300 1822.160 2914.100 1822.640 ;
        RECT 5.520 1816.720 13.700 1817.200 ;
        RECT 2906.300 1816.720 2914.100 1817.200 ;
        RECT 5.520 1811.280 13.700 1811.760 ;
        RECT 2906.300 1811.280 2914.100 1811.760 ;
        RECT 5.520 1805.840 13.700 1806.320 ;
        RECT 2906.300 1805.840 2914.100 1806.320 ;
        RECT 5.520 1800.400 13.700 1800.880 ;
        RECT 2906.300 1800.400 2914.100 1800.880 ;
        RECT 5.520 1794.960 13.700 1795.440 ;
        RECT 2906.300 1794.960 2914.100 1795.440 ;
        RECT 5.520 1789.520 13.700 1790.000 ;
        RECT 2906.300 1789.520 2914.100 1790.000 ;
        RECT 5.520 1784.080 13.700 1784.560 ;
        RECT 2906.300 1784.080 2914.100 1784.560 ;
        RECT 5.520 1778.640 13.700 1779.120 ;
        RECT 2906.300 1778.640 2914.100 1779.120 ;
        RECT 5.520 1773.200 13.700 1773.680 ;
        RECT 2906.300 1773.200 2914.100 1773.680 ;
        RECT 5.520 1767.760 13.700 1768.240 ;
        RECT 2906.300 1767.760 2914.100 1768.240 ;
        RECT 5.520 1762.320 13.700 1762.800 ;
        RECT 2906.300 1762.320 2914.100 1762.800 ;
        RECT 5.520 1756.880 13.700 1757.360 ;
        RECT 2906.300 1756.880 2914.100 1757.360 ;
        RECT 5.520 1751.440 13.700 1751.920 ;
        RECT 2906.300 1751.440 2914.100 1751.920 ;
        RECT 5.520 1746.000 13.700 1746.480 ;
        RECT 2906.300 1746.000 2914.100 1746.480 ;
        RECT 5.520 1740.560 13.700 1741.040 ;
        RECT 2906.300 1740.560 2914.100 1741.040 ;
        RECT 5.520 1735.120 13.700 1735.600 ;
        RECT 2906.300 1735.120 2914.100 1735.600 ;
        RECT 5.520 1729.680 13.700 1730.160 ;
        RECT 2906.300 1729.680 2914.100 1730.160 ;
        RECT 5.520 1724.240 13.700 1724.720 ;
        RECT 2906.300 1724.240 2914.100 1724.720 ;
        RECT 5.520 1718.800 13.700 1719.280 ;
        RECT 2906.300 1718.800 2914.100 1719.280 ;
        RECT 5.520 1713.360 13.700 1713.840 ;
        RECT 2906.300 1713.360 2914.100 1713.840 ;
        RECT 5.520 1707.920 13.700 1708.400 ;
        RECT 2906.300 1707.920 2914.100 1708.400 ;
        RECT 5.520 1702.480 13.700 1702.960 ;
        RECT 2906.300 1702.480 2914.100 1702.960 ;
        RECT 5.520 1697.040 13.700 1697.520 ;
        RECT 2906.300 1697.040 2914.100 1697.520 ;
        RECT 5.520 1691.600 13.700 1692.080 ;
        RECT 2906.300 1691.600 2914.100 1692.080 ;
        RECT 5.520 1686.160 13.700 1686.640 ;
        RECT 2906.300 1686.160 2914.100 1686.640 ;
        RECT 5.520 1680.720 13.700 1681.200 ;
        RECT 2906.300 1680.720 2914.100 1681.200 ;
        RECT 5.520 1675.280 13.700 1675.760 ;
        RECT 2906.300 1675.280 2914.100 1675.760 ;
        RECT 5.520 1669.840 13.700 1670.320 ;
        RECT 2906.300 1669.840 2914.100 1670.320 ;
        RECT 5.520 1664.400 13.700 1664.880 ;
        RECT 2906.300 1664.400 2914.100 1664.880 ;
        RECT 5.520 1658.960 13.700 1659.440 ;
        RECT 2906.300 1658.960 2914.100 1659.440 ;
        RECT 5.520 1653.520 13.700 1654.000 ;
        RECT 2906.300 1653.520 2914.100 1654.000 ;
        RECT 5.520 1648.080 13.700 1648.560 ;
        RECT 2906.300 1648.080 2914.100 1648.560 ;
        RECT 5.520 1642.640 13.700 1643.120 ;
        RECT 2906.300 1642.640 2914.100 1643.120 ;
        RECT 5.520 1637.200 13.700 1637.680 ;
        RECT 2906.300 1637.200 2914.100 1637.680 ;
        RECT 5.520 1631.760 13.700 1632.240 ;
        RECT 2906.300 1631.760 2914.100 1632.240 ;
        RECT 5.520 1626.320 13.700 1626.800 ;
        RECT 2906.300 1626.320 2914.100 1626.800 ;
        RECT 5.520 1620.880 13.700 1621.360 ;
        RECT 2906.300 1620.880 2914.100 1621.360 ;
        RECT 5.520 1615.440 13.700 1615.920 ;
        RECT 2906.300 1615.440 2914.100 1615.920 ;
        RECT 5.520 1610.000 13.700 1610.480 ;
        RECT 2906.300 1610.000 2914.100 1610.480 ;
        RECT 5.520 1604.560 13.700 1605.040 ;
        RECT 2906.300 1604.560 2914.100 1605.040 ;
        RECT 5.520 1599.120 13.700 1599.600 ;
        RECT 2906.300 1599.120 2914.100 1599.600 ;
        RECT 5.520 1593.680 13.700 1594.160 ;
        RECT 2906.300 1593.680 2914.100 1594.160 ;
        RECT 5.520 1588.240 13.700 1588.720 ;
        RECT 2906.300 1588.240 2914.100 1588.720 ;
        RECT 5.520 1582.800 13.700 1583.280 ;
        RECT 2906.300 1582.800 2914.100 1583.280 ;
        RECT 5.520 1577.360 13.700 1577.840 ;
        RECT 2906.300 1577.360 2914.100 1577.840 ;
        RECT 5.520 1571.920 13.700 1572.400 ;
        RECT 2906.300 1571.920 2914.100 1572.400 ;
        RECT 5.520 1566.480 13.700 1566.960 ;
        RECT 2906.300 1566.480 2914.100 1566.960 ;
        RECT 5.520 1561.040 13.700 1561.520 ;
        RECT 2906.300 1561.040 2914.100 1561.520 ;
        RECT 5.520 1555.600 13.700 1556.080 ;
        RECT 2906.300 1555.600 2914.100 1556.080 ;
        RECT 5.520 1550.160 13.700 1550.640 ;
        RECT 2906.300 1550.160 2914.100 1550.640 ;
        RECT 5.520 1544.720 13.700 1545.200 ;
        RECT 2906.300 1544.720 2914.100 1545.200 ;
        RECT 5.520 1539.280 13.700 1539.760 ;
        RECT 2906.300 1539.280 2914.100 1539.760 ;
        RECT 5.520 1533.840 13.700 1534.320 ;
        RECT 2906.300 1533.840 2914.100 1534.320 ;
        RECT 5.520 1528.400 13.700 1528.880 ;
        RECT 2906.300 1528.400 2914.100 1528.880 ;
        RECT 5.520 1522.960 13.700 1523.440 ;
        RECT 2906.300 1522.960 2914.100 1523.440 ;
        RECT 5.520 1517.520 13.700 1518.000 ;
        RECT 2906.300 1517.520 2914.100 1518.000 ;
        RECT 5.520 1512.080 13.700 1512.560 ;
        RECT 2906.300 1512.080 2914.100 1512.560 ;
        RECT 5.520 1506.640 13.700 1507.120 ;
        RECT 2906.300 1506.640 2914.100 1507.120 ;
        RECT 5.520 1501.200 13.700 1501.680 ;
        RECT 2906.300 1501.200 2914.100 1501.680 ;
        RECT 5.520 1495.760 13.700 1496.240 ;
        RECT 2906.300 1495.760 2914.100 1496.240 ;
        RECT 5.520 1490.320 13.700 1490.800 ;
        RECT 2906.300 1490.320 2914.100 1490.800 ;
        RECT 5.520 1484.880 13.700 1485.360 ;
        RECT 2906.300 1484.880 2914.100 1485.360 ;
        RECT 5.520 1479.440 13.700 1479.920 ;
        RECT 2906.300 1479.440 2914.100 1479.920 ;
        RECT 5.520 1474.000 13.700 1474.480 ;
        RECT 2906.300 1474.000 2914.100 1474.480 ;
        RECT 5.520 1468.560 13.700 1469.040 ;
        RECT 2906.300 1468.560 2914.100 1469.040 ;
        RECT 5.520 1463.120 13.700 1463.600 ;
        RECT 2906.300 1463.120 2914.100 1463.600 ;
        RECT 5.520 1457.680 13.700 1458.160 ;
        RECT 2906.300 1457.680 2914.100 1458.160 ;
        RECT 5.520 1452.240 13.700 1452.720 ;
        RECT 2906.300 1452.240 2914.100 1452.720 ;
        RECT 5.520 1446.800 13.700 1447.280 ;
        RECT 2906.300 1446.800 2914.100 1447.280 ;
        RECT 5.520 1441.360 13.700 1441.840 ;
        RECT 2906.300 1441.360 2914.100 1441.840 ;
        RECT 5.520 1435.920 13.700 1436.400 ;
        RECT 2906.300 1435.920 2914.100 1436.400 ;
        RECT 5.520 1430.480 13.700 1430.960 ;
        RECT 2906.300 1430.480 2914.100 1430.960 ;
        RECT 5.520 1425.040 13.700 1425.520 ;
        RECT 2906.300 1425.040 2914.100 1425.520 ;
        RECT 5.520 1419.600 13.700 1420.080 ;
        RECT 2906.300 1419.600 2914.100 1420.080 ;
        RECT 5.520 1414.160 13.700 1414.640 ;
        RECT 2906.300 1414.160 2914.100 1414.640 ;
        RECT 5.520 1408.720 13.700 1409.200 ;
        RECT 2906.300 1408.720 2914.100 1409.200 ;
        RECT 5.520 1403.280 13.700 1403.760 ;
        RECT 2906.300 1403.280 2914.100 1403.760 ;
        RECT 5.520 1397.840 13.700 1398.320 ;
        RECT 2906.300 1397.840 2914.100 1398.320 ;
        RECT 5.520 1392.400 13.700 1392.880 ;
        RECT 2906.300 1392.400 2914.100 1392.880 ;
        RECT 5.520 1386.960 13.700 1387.440 ;
        RECT 2906.300 1386.960 2914.100 1387.440 ;
        RECT 5.520 1381.520 13.700 1382.000 ;
        RECT 2906.300 1381.520 2914.100 1382.000 ;
        RECT 5.520 1376.080 13.700 1376.560 ;
        RECT 2906.300 1376.080 2914.100 1376.560 ;
        RECT 5.520 1370.640 13.700 1371.120 ;
        RECT 2906.300 1370.640 2914.100 1371.120 ;
        RECT 5.520 1365.200 13.700 1365.680 ;
        RECT 2906.300 1365.200 2914.100 1365.680 ;
        RECT 5.520 1359.760 13.700 1360.240 ;
        RECT 2906.300 1359.760 2914.100 1360.240 ;
        RECT 5.520 1354.320 13.700 1354.800 ;
        RECT 2906.300 1354.320 2914.100 1354.800 ;
        RECT 5.520 1348.880 13.700 1349.360 ;
        RECT 2906.300 1348.880 2914.100 1349.360 ;
        RECT 5.520 1343.440 13.700 1343.920 ;
        RECT 2906.300 1343.440 2914.100 1343.920 ;
        RECT 5.520 1338.000 13.700 1338.480 ;
        RECT 2906.300 1338.000 2914.100 1338.480 ;
        RECT 5.520 1332.560 13.700 1333.040 ;
        RECT 2906.300 1332.560 2914.100 1333.040 ;
        RECT 5.520 1327.120 13.700 1327.600 ;
        RECT 2906.300 1327.120 2914.100 1327.600 ;
        RECT 5.520 1321.680 13.700 1322.160 ;
        RECT 2906.300 1321.680 2914.100 1322.160 ;
        RECT 5.520 1316.240 13.700 1316.720 ;
        RECT 2906.300 1316.240 2914.100 1316.720 ;
        RECT 5.520 1310.800 13.700 1311.280 ;
        RECT 2906.300 1310.800 2914.100 1311.280 ;
        RECT 5.520 1305.360 13.700 1305.840 ;
        RECT 2906.300 1305.360 2914.100 1305.840 ;
        RECT 5.520 1299.920 13.700 1300.400 ;
        RECT 2906.300 1299.920 2914.100 1300.400 ;
        RECT 5.520 1294.480 13.700 1294.960 ;
        RECT 2906.300 1294.480 2914.100 1294.960 ;
        RECT 5.520 1289.040 13.700 1289.520 ;
        RECT 2906.300 1289.040 2914.100 1289.520 ;
        RECT 5.520 1283.600 13.700 1284.080 ;
        RECT 2906.300 1283.600 2914.100 1284.080 ;
        RECT 5.520 1278.160 13.700 1278.640 ;
        RECT 2906.300 1278.160 2914.100 1278.640 ;
        RECT 5.520 1272.720 13.700 1273.200 ;
        RECT 2906.300 1272.720 2914.100 1273.200 ;
        RECT 5.520 1267.280 13.700 1267.760 ;
        RECT 2906.300 1267.280 2914.100 1267.760 ;
        RECT 5.520 1261.840 13.700 1262.320 ;
        RECT 2906.300 1261.840 2914.100 1262.320 ;
        RECT 5.520 1256.400 13.700 1256.880 ;
        RECT 2906.300 1256.400 2914.100 1256.880 ;
        RECT 5.520 1250.960 13.700 1251.440 ;
        RECT 2906.300 1250.960 2914.100 1251.440 ;
        RECT 5.520 1245.520 13.700 1246.000 ;
        RECT 2906.300 1245.520 2914.100 1246.000 ;
        RECT 5.520 1240.080 13.700 1240.560 ;
        RECT 2906.300 1240.080 2914.100 1240.560 ;
        RECT 5.520 1234.640 13.700 1235.120 ;
        RECT 2906.300 1234.640 2914.100 1235.120 ;
        RECT 5.520 1229.200 13.700 1229.680 ;
        RECT 2906.300 1229.200 2914.100 1229.680 ;
        RECT 5.520 1223.760 13.700 1224.240 ;
        RECT 2906.300 1223.760 2914.100 1224.240 ;
        RECT 5.520 1218.320 13.700 1218.800 ;
        RECT 2906.300 1218.320 2914.100 1218.800 ;
        RECT 5.520 1212.880 13.700 1213.360 ;
        RECT 2906.300 1212.880 2914.100 1213.360 ;
        RECT 5.520 1207.440 13.700 1207.920 ;
        RECT 2906.300 1207.440 2914.100 1207.920 ;
        RECT 5.520 1202.000 13.700 1202.480 ;
        RECT 2906.300 1202.000 2914.100 1202.480 ;
        RECT 5.520 1196.560 13.700 1197.040 ;
        RECT 2906.300 1196.560 2914.100 1197.040 ;
        RECT 5.520 1191.120 13.700 1191.600 ;
        RECT 2906.300 1191.120 2914.100 1191.600 ;
        RECT 5.520 1185.680 13.700 1186.160 ;
        RECT 2906.300 1185.680 2914.100 1186.160 ;
        RECT 5.520 1180.240 13.700 1180.720 ;
        RECT 2906.300 1180.240 2914.100 1180.720 ;
        RECT 5.520 1174.800 13.700 1175.280 ;
        RECT 2906.300 1174.800 2914.100 1175.280 ;
        RECT 5.520 1169.360 13.700 1169.840 ;
        RECT 2906.300 1169.360 2914.100 1169.840 ;
        RECT 5.520 1163.920 13.700 1164.400 ;
        RECT 2906.300 1163.920 2914.100 1164.400 ;
        RECT 5.520 1158.480 13.700 1158.960 ;
        RECT 2906.300 1158.480 2914.100 1158.960 ;
        RECT 5.520 1153.040 13.700 1153.520 ;
        RECT 2906.300 1153.040 2914.100 1153.520 ;
        RECT 5.520 1147.600 13.700 1148.080 ;
        RECT 2906.300 1147.600 2914.100 1148.080 ;
        RECT 5.520 1142.160 13.700 1142.640 ;
        RECT 2906.300 1142.160 2914.100 1142.640 ;
        RECT 5.520 1136.720 13.700 1137.200 ;
        RECT 2906.300 1136.720 2914.100 1137.200 ;
        RECT 5.520 1131.280 13.700 1131.760 ;
        RECT 2906.300 1131.280 2914.100 1131.760 ;
        RECT 5.520 1125.840 13.700 1126.320 ;
        RECT 2906.300 1125.840 2914.100 1126.320 ;
        RECT 5.520 1120.400 13.700 1120.880 ;
        RECT 2906.300 1120.400 2914.100 1120.880 ;
        RECT 5.520 1114.960 13.700 1115.440 ;
        RECT 2906.300 1114.960 2914.100 1115.440 ;
        RECT 5.520 1109.520 13.700 1110.000 ;
        RECT 2906.300 1109.520 2914.100 1110.000 ;
        RECT 5.520 1104.080 13.700 1104.560 ;
        RECT 2906.300 1104.080 2914.100 1104.560 ;
        RECT 5.520 1098.640 13.700 1099.120 ;
        RECT 2906.300 1098.640 2914.100 1099.120 ;
        RECT 5.520 1093.200 13.700 1093.680 ;
        RECT 2906.300 1093.200 2914.100 1093.680 ;
        RECT 5.520 1087.760 13.700 1088.240 ;
        RECT 2906.300 1087.760 2914.100 1088.240 ;
        RECT 5.520 1082.320 13.700 1082.800 ;
        RECT 2906.300 1082.320 2914.100 1082.800 ;
        RECT 5.520 1076.880 13.700 1077.360 ;
        RECT 2906.300 1076.880 2914.100 1077.360 ;
        RECT 5.520 1071.440 13.700 1071.920 ;
        RECT 2906.300 1071.440 2914.100 1071.920 ;
        RECT 5.520 1066.000 13.700 1066.480 ;
        RECT 2906.300 1066.000 2914.100 1066.480 ;
        RECT 5.520 1060.560 13.700 1061.040 ;
        RECT 2906.300 1060.560 2914.100 1061.040 ;
        RECT 5.520 1055.120 13.700 1055.600 ;
        RECT 2906.300 1055.120 2914.100 1055.600 ;
        RECT 5.520 1049.680 13.700 1050.160 ;
        RECT 2906.300 1049.680 2914.100 1050.160 ;
        RECT 5.520 1044.240 13.700 1044.720 ;
        RECT 2906.300 1044.240 2914.100 1044.720 ;
        RECT 5.520 1038.800 13.700 1039.280 ;
        RECT 2906.300 1038.800 2914.100 1039.280 ;
        RECT 5.520 1033.360 13.700 1033.840 ;
        RECT 2906.300 1033.360 2914.100 1033.840 ;
        RECT 5.520 1027.920 13.700 1028.400 ;
        RECT 2906.300 1027.920 2914.100 1028.400 ;
        RECT 5.520 1022.480 13.700 1022.960 ;
        RECT 2906.300 1022.480 2914.100 1022.960 ;
        RECT 5.520 1017.040 13.700 1017.520 ;
        RECT 2906.300 1017.040 2914.100 1017.520 ;
        RECT 5.520 1011.600 13.700 1012.080 ;
        RECT 2906.300 1011.600 2914.100 1012.080 ;
        RECT 5.520 1006.160 13.700 1006.640 ;
        RECT 2906.300 1006.160 2914.100 1006.640 ;
        RECT 5.520 1000.720 13.700 1001.200 ;
        RECT 2906.300 1000.720 2914.100 1001.200 ;
        RECT 5.520 995.280 13.700 995.760 ;
        RECT 2906.300 995.280 2914.100 995.760 ;
        RECT 5.520 989.840 13.700 990.320 ;
        RECT 2906.300 989.840 2914.100 990.320 ;
        RECT 5.520 984.400 13.700 984.880 ;
        RECT 2906.300 984.400 2914.100 984.880 ;
        RECT 5.520 978.960 13.700 979.440 ;
        RECT 2906.300 978.960 2914.100 979.440 ;
        RECT 5.520 973.520 13.700 974.000 ;
        RECT 2906.300 973.520 2914.100 974.000 ;
        RECT 5.520 968.080 13.700 968.560 ;
        RECT 2906.300 968.080 2914.100 968.560 ;
        RECT 5.520 962.640 13.700 963.120 ;
        RECT 2906.300 962.640 2914.100 963.120 ;
        RECT 5.520 957.200 13.700 957.680 ;
        RECT 2906.300 957.200 2914.100 957.680 ;
        RECT 5.520 951.760 13.700 952.240 ;
        RECT 2906.300 951.760 2914.100 952.240 ;
        RECT 5.520 946.320 13.700 946.800 ;
        RECT 2906.300 946.320 2914.100 946.800 ;
        RECT 5.520 940.880 13.700 941.360 ;
        RECT 2906.300 940.880 2914.100 941.360 ;
        RECT 5.520 935.440 13.700 935.920 ;
        RECT 2906.300 935.440 2914.100 935.920 ;
        RECT 5.520 930.000 13.700 930.480 ;
        RECT 2906.300 930.000 2914.100 930.480 ;
        RECT 5.520 924.560 13.700 925.040 ;
        RECT 2906.300 924.560 2914.100 925.040 ;
        RECT 5.520 919.120 13.700 919.600 ;
        RECT 2906.300 919.120 2914.100 919.600 ;
        RECT 5.520 913.680 13.700 914.160 ;
        RECT 2906.300 913.680 2914.100 914.160 ;
        RECT 5.520 908.240 13.700 908.720 ;
        RECT 2906.300 908.240 2914.100 908.720 ;
        RECT 5.520 902.800 13.700 903.280 ;
        RECT 2906.300 902.800 2914.100 903.280 ;
        RECT 5.520 897.360 13.700 897.840 ;
        RECT 2906.300 897.360 2914.100 897.840 ;
        RECT 5.520 891.920 13.700 892.400 ;
        RECT 2906.300 891.920 2914.100 892.400 ;
        RECT 5.520 886.480 13.700 886.960 ;
        RECT 2906.300 886.480 2914.100 886.960 ;
        RECT 5.520 881.040 13.700 881.520 ;
        RECT 2906.300 881.040 2914.100 881.520 ;
        RECT 5.520 875.600 13.700 876.080 ;
        RECT 2906.300 875.600 2914.100 876.080 ;
        RECT 5.520 870.160 13.700 870.640 ;
        RECT 2906.300 870.160 2914.100 870.640 ;
        RECT 5.520 864.720 13.700 865.200 ;
        RECT 2906.300 864.720 2914.100 865.200 ;
        RECT 5.520 859.280 13.700 859.760 ;
        RECT 2906.300 859.280 2914.100 859.760 ;
        RECT 5.520 853.840 13.700 854.320 ;
        RECT 2906.300 853.840 2914.100 854.320 ;
        RECT 5.520 848.400 13.700 848.880 ;
        RECT 2906.300 848.400 2914.100 848.880 ;
        RECT 5.520 842.960 13.700 843.440 ;
        RECT 2906.300 842.960 2914.100 843.440 ;
        RECT 5.520 837.520 13.700 838.000 ;
        RECT 2906.300 837.520 2914.100 838.000 ;
        RECT 5.520 832.080 13.700 832.560 ;
        RECT 2906.300 832.080 2914.100 832.560 ;
        RECT 5.520 826.640 13.700 827.120 ;
        RECT 2906.300 826.640 2914.100 827.120 ;
        RECT 5.520 821.200 13.700 821.680 ;
        RECT 2906.300 821.200 2914.100 821.680 ;
        RECT 5.520 815.760 13.700 816.240 ;
        RECT 2906.300 815.760 2914.100 816.240 ;
        RECT 5.520 810.320 13.700 810.800 ;
        RECT 2906.300 810.320 2914.100 810.800 ;
        RECT 5.520 804.880 13.700 805.360 ;
        RECT 2906.300 804.880 2914.100 805.360 ;
        RECT 5.520 799.440 13.700 799.920 ;
        RECT 2906.300 799.440 2914.100 799.920 ;
        RECT 5.520 794.000 13.700 794.480 ;
        RECT 2906.300 794.000 2914.100 794.480 ;
        RECT 5.520 788.560 13.700 789.040 ;
        RECT 2906.300 788.560 2914.100 789.040 ;
        RECT 5.520 783.120 13.700 783.600 ;
        RECT 2906.300 783.120 2914.100 783.600 ;
        RECT 5.520 777.680 13.700 778.160 ;
        RECT 2906.300 777.680 2914.100 778.160 ;
        RECT 5.520 772.240 13.700 772.720 ;
        RECT 2906.300 772.240 2914.100 772.720 ;
        RECT 5.520 766.800 13.700 767.280 ;
        RECT 2906.300 766.800 2914.100 767.280 ;
        RECT 5.520 761.360 13.700 761.840 ;
        RECT 2906.300 761.360 2914.100 761.840 ;
        RECT 5.520 755.920 13.700 756.400 ;
        RECT 2906.300 755.920 2914.100 756.400 ;
        RECT 5.520 750.480 13.700 750.960 ;
        RECT 2906.300 750.480 2914.100 750.960 ;
        RECT 5.520 745.040 13.700 745.520 ;
        RECT 2906.300 745.040 2914.100 745.520 ;
        RECT 5.520 739.600 13.700 740.080 ;
        RECT 2906.300 739.600 2914.100 740.080 ;
        RECT 5.520 734.160 13.700 734.640 ;
        RECT 2906.300 734.160 2914.100 734.640 ;
        RECT 5.520 728.720 13.700 729.200 ;
        RECT 2906.300 728.720 2914.100 729.200 ;
        RECT 5.520 723.280 13.700 723.760 ;
        RECT 2906.300 723.280 2914.100 723.760 ;
        RECT 5.520 717.840 13.700 718.320 ;
        RECT 2906.300 717.840 2914.100 718.320 ;
        RECT 5.520 712.400 13.700 712.880 ;
        RECT 2906.300 712.400 2914.100 712.880 ;
        RECT 5.520 706.960 13.700 707.440 ;
        RECT 2906.300 706.960 2914.100 707.440 ;
        RECT 5.520 701.520 13.700 702.000 ;
        RECT 2906.300 701.520 2914.100 702.000 ;
        RECT 5.520 696.080 13.700 696.560 ;
        RECT 2906.300 696.080 2914.100 696.560 ;
        RECT 5.520 690.640 13.700 691.120 ;
        RECT 2906.300 690.640 2914.100 691.120 ;
        RECT 5.520 685.200 13.700 685.680 ;
        RECT 2906.300 685.200 2914.100 685.680 ;
        RECT 5.520 679.760 13.700 680.240 ;
        RECT 2906.300 679.760 2914.100 680.240 ;
        RECT 5.520 674.320 13.700 674.800 ;
        RECT 2906.300 674.320 2914.100 674.800 ;
        RECT 5.520 668.880 13.700 669.360 ;
        RECT 2906.300 668.880 2914.100 669.360 ;
        RECT 5.520 663.440 13.700 663.920 ;
        RECT 2906.300 663.440 2914.100 663.920 ;
        RECT 5.520 658.000 13.700 658.480 ;
        RECT 2906.300 658.000 2914.100 658.480 ;
        RECT 5.520 652.560 13.700 653.040 ;
        RECT 2906.300 652.560 2914.100 653.040 ;
        RECT 5.520 647.120 13.700 647.600 ;
        RECT 2906.300 647.120 2914.100 647.600 ;
        RECT 5.520 641.680 13.700 642.160 ;
        RECT 2906.300 641.680 2914.100 642.160 ;
        RECT 5.520 636.240 13.700 636.720 ;
        RECT 2906.300 636.240 2914.100 636.720 ;
        RECT 5.520 630.800 13.700 631.280 ;
        RECT 2906.300 630.800 2914.100 631.280 ;
        RECT 5.520 625.360 13.700 625.840 ;
        RECT 2906.300 625.360 2914.100 625.840 ;
        RECT 5.520 619.920 13.700 620.400 ;
        RECT 2906.300 619.920 2914.100 620.400 ;
        RECT 5.520 614.480 13.700 614.960 ;
        RECT 2906.300 614.480 2914.100 614.960 ;
        RECT 5.520 609.040 13.700 609.520 ;
        RECT 2906.300 609.040 2914.100 609.520 ;
        RECT 5.520 603.600 13.700 604.080 ;
        RECT 2906.300 603.600 2914.100 604.080 ;
        RECT 5.520 598.160 13.700 598.640 ;
        RECT 2906.300 598.160 2914.100 598.640 ;
        RECT 5.520 592.720 13.700 593.200 ;
        RECT 2906.300 592.720 2914.100 593.200 ;
        RECT 5.520 587.280 13.700 587.760 ;
        RECT 2906.300 587.280 2914.100 587.760 ;
        RECT 5.520 581.840 13.700 582.320 ;
        RECT 2906.300 581.840 2914.100 582.320 ;
        RECT 5.520 576.400 13.700 576.880 ;
        RECT 2906.300 576.400 2914.100 576.880 ;
        RECT 5.520 570.960 13.700 571.440 ;
        RECT 2906.300 570.960 2914.100 571.440 ;
        RECT 5.520 565.520 13.700 566.000 ;
        RECT 2906.300 565.520 2914.100 566.000 ;
        RECT 5.520 560.080 13.700 560.560 ;
        RECT 2906.300 560.080 2914.100 560.560 ;
        RECT 5.520 554.640 13.700 555.120 ;
        RECT 2906.300 554.640 2914.100 555.120 ;
        RECT 5.520 549.200 13.700 549.680 ;
        RECT 2906.300 549.200 2914.100 549.680 ;
        RECT 5.520 543.760 13.700 544.240 ;
        RECT 2906.300 543.760 2914.100 544.240 ;
        RECT 5.520 538.320 13.700 538.800 ;
        RECT 2906.300 538.320 2914.100 538.800 ;
        RECT 5.520 532.880 13.700 533.360 ;
        RECT 2906.300 532.880 2914.100 533.360 ;
        RECT 5.520 527.440 13.700 527.920 ;
        RECT 2906.300 527.440 2914.100 527.920 ;
        RECT 5.520 522.000 13.700 522.480 ;
        RECT 2906.300 522.000 2914.100 522.480 ;
        RECT 5.520 516.560 13.700 517.040 ;
        RECT 2906.300 516.560 2914.100 517.040 ;
        RECT 5.520 511.120 13.700 511.600 ;
        RECT 2906.300 511.120 2914.100 511.600 ;
        RECT 5.520 505.680 13.700 506.160 ;
        RECT 2906.300 505.680 2914.100 506.160 ;
        RECT 5.520 500.240 13.700 500.720 ;
        RECT 2906.300 500.240 2914.100 500.720 ;
        RECT 5.520 494.800 13.700 495.280 ;
        RECT 2906.300 494.800 2914.100 495.280 ;
        RECT 5.520 489.360 13.700 489.840 ;
        RECT 2906.300 489.360 2914.100 489.840 ;
        RECT 5.520 483.920 13.700 484.400 ;
        RECT 2906.300 483.920 2914.100 484.400 ;
        RECT 5.520 478.480 13.700 478.960 ;
        RECT 2906.300 478.480 2914.100 478.960 ;
        RECT 5.520 473.040 13.700 473.520 ;
        RECT 2906.300 473.040 2914.100 473.520 ;
        RECT 5.520 467.600 13.700 468.080 ;
        RECT 2906.300 467.600 2914.100 468.080 ;
        RECT 5.520 462.160 13.700 462.640 ;
        RECT 2906.300 462.160 2914.100 462.640 ;
        RECT 5.520 456.720 13.700 457.200 ;
        RECT 2906.300 456.720 2914.100 457.200 ;
        RECT 5.520 451.280 13.700 451.760 ;
        RECT 2906.300 451.280 2914.100 451.760 ;
        RECT 5.520 445.840 13.700 446.320 ;
        RECT 2906.300 445.840 2914.100 446.320 ;
        RECT 5.520 440.400 13.700 440.880 ;
        RECT 2906.300 440.400 2914.100 440.880 ;
        RECT 5.520 434.960 13.700 435.440 ;
        RECT 2906.300 434.960 2914.100 435.440 ;
        RECT 5.520 429.520 13.700 430.000 ;
        RECT 2906.300 429.520 2914.100 430.000 ;
        RECT 5.520 424.080 13.700 424.560 ;
        RECT 2906.300 424.080 2914.100 424.560 ;
        RECT 5.520 418.640 13.700 419.120 ;
        RECT 2906.300 418.640 2914.100 419.120 ;
        RECT 5.520 413.200 13.700 413.680 ;
        RECT 2906.300 413.200 2914.100 413.680 ;
        RECT 5.520 407.760 13.700 408.240 ;
        RECT 2906.300 407.760 2914.100 408.240 ;
        RECT 5.520 402.320 13.700 402.800 ;
        RECT 2906.300 402.320 2914.100 402.800 ;
        RECT 5.520 396.880 13.700 397.360 ;
        RECT 2906.300 396.880 2914.100 397.360 ;
        RECT 5.520 391.440 13.700 391.920 ;
        RECT 2906.300 391.440 2914.100 391.920 ;
        RECT 5.520 386.000 13.700 386.480 ;
        RECT 2906.300 386.000 2914.100 386.480 ;
        RECT 5.520 380.560 13.700 381.040 ;
        RECT 2906.300 380.560 2914.100 381.040 ;
        RECT 5.520 375.120 13.700 375.600 ;
        RECT 2906.300 375.120 2914.100 375.600 ;
        RECT 5.520 369.680 13.700 370.160 ;
        RECT 2906.300 369.680 2914.100 370.160 ;
        RECT 5.520 364.240 13.700 364.720 ;
        RECT 2906.300 364.240 2914.100 364.720 ;
        RECT 5.520 358.800 13.700 359.280 ;
        RECT 2906.300 358.800 2914.100 359.280 ;
        RECT 5.520 353.360 13.700 353.840 ;
        RECT 2906.300 353.360 2914.100 353.840 ;
        RECT 5.520 347.920 13.700 348.400 ;
        RECT 2906.300 347.920 2914.100 348.400 ;
        RECT 5.520 342.480 13.700 342.960 ;
        RECT 2906.300 342.480 2914.100 342.960 ;
        RECT 5.520 337.040 13.700 337.520 ;
        RECT 2906.300 337.040 2914.100 337.520 ;
        RECT 5.520 331.600 13.700 332.080 ;
        RECT 2906.300 331.600 2914.100 332.080 ;
        RECT 5.520 326.160 13.700 326.640 ;
        RECT 2906.300 326.160 2914.100 326.640 ;
        RECT 5.520 320.720 13.700 321.200 ;
        RECT 2906.300 320.720 2914.100 321.200 ;
        RECT 5.520 315.280 13.700 315.760 ;
        RECT 2906.300 315.280 2914.100 315.760 ;
        RECT 5.520 309.840 13.700 310.320 ;
        RECT 2906.300 309.840 2914.100 310.320 ;
        RECT 5.520 304.400 13.700 304.880 ;
        RECT 2906.300 304.400 2914.100 304.880 ;
        RECT 5.520 298.960 13.700 299.440 ;
        RECT 2906.300 298.960 2914.100 299.440 ;
        RECT 5.520 293.520 13.700 294.000 ;
        RECT 2906.300 293.520 2914.100 294.000 ;
        RECT 5.520 288.080 13.700 288.560 ;
        RECT 2906.300 288.080 2914.100 288.560 ;
        RECT 5.520 282.640 13.700 283.120 ;
        RECT 2906.300 282.640 2914.100 283.120 ;
        RECT 5.520 277.200 13.700 277.680 ;
        RECT 2906.300 277.200 2914.100 277.680 ;
        RECT 5.520 271.760 13.700 272.240 ;
        RECT 2906.300 271.760 2914.100 272.240 ;
        RECT 5.520 266.320 13.700 266.800 ;
        RECT 2906.300 266.320 2914.100 266.800 ;
        RECT 5.520 260.880 13.700 261.360 ;
        RECT 2906.300 260.880 2914.100 261.360 ;
        RECT 5.520 255.440 13.700 255.920 ;
        RECT 2906.300 255.440 2914.100 255.920 ;
        RECT 5.520 250.000 13.700 250.480 ;
        RECT 2906.300 250.000 2914.100 250.480 ;
        RECT 5.520 244.560 13.700 245.040 ;
        RECT 2906.300 244.560 2914.100 245.040 ;
        RECT 5.520 239.120 13.700 239.600 ;
        RECT 2906.300 239.120 2914.100 239.600 ;
        RECT 5.520 233.680 13.700 234.160 ;
        RECT 2906.300 233.680 2914.100 234.160 ;
        RECT 5.520 228.240 13.700 228.720 ;
        RECT 2906.300 228.240 2914.100 228.720 ;
        RECT 5.520 222.800 13.700 223.280 ;
        RECT 2906.300 222.800 2914.100 223.280 ;
        RECT 5.520 217.360 13.700 217.840 ;
        RECT 2906.300 217.360 2914.100 217.840 ;
        RECT 5.520 211.920 13.700 212.400 ;
        RECT 2906.300 211.920 2914.100 212.400 ;
        RECT 5.520 206.480 13.700 206.960 ;
        RECT 2906.300 206.480 2914.100 206.960 ;
        RECT 5.520 201.040 13.700 201.520 ;
        RECT 2906.300 201.040 2914.100 201.520 ;
        RECT 5.520 195.600 13.700 196.080 ;
        RECT 2906.300 195.600 2914.100 196.080 ;
        RECT 5.520 190.160 13.700 190.640 ;
        RECT 2906.300 190.160 2914.100 190.640 ;
        RECT 5.520 184.720 13.700 185.200 ;
        RECT 2906.300 184.720 2914.100 185.200 ;
        RECT 5.520 179.280 13.700 179.760 ;
        RECT 2906.300 179.280 2914.100 179.760 ;
        RECT 5.520 173.840 13.700 174.320 ;
        RECT 2906.300 173.840 2914.100 174.320 ;
        RECT 5.520 168.400 13.700 168.880 ;
        RECT 2906.300 168.400 2914.100 168.880 ;
        RECT 5.520 162.960 13.700 163.440 ;
        RECT 2906.300 162.960 2914.100 163.440 ;
        RECT 5.520 157.520 13.700 158.000 ;
        RECT 2906.300 157.520 2914.100 158.000 ;
        RECT 5.520 152.080 13.700 152.560 ;
        RECT 2906.300 152.080 2914.100 152.560 ;
        RECT 5.520 146.640 13.700 147.120 ;
        RECT 2906.300 146.640 2914.100 147.120 ;
        RECT 5.520 141.200 13.700 141.680 ;
        RECT 2906.300 141.200 2914.100 141.680 ;
        RECT 5.520 135.760 13.700 136.240 ;
        RECT 2906.300 135.760 2914.100 136.240 ;
        RECT 5.520 130.320 13.700 130.800 ;
        RECT 2906.300 130.320 2914.100 130.800 ;
        RECT 5.520 124.880 13.700 125.360 ;
        RECT 2906.300 124.880 2914.100 125.360 ;
        RECT 5.520 119.440 13.700 119.920 ;
        RECT 2906.300 119.440 2914.100 119.920 ;
        RECT 5.520 114.000 13.700 114.480 ;
        RECT 2906.300 114.000 2914.100 114.480 ;
        RECT 5.520 108.560 13.700 109.040 ;
        RECT 2906.300 108.560 2914.100 109.040 ;
        RECT 5.520 103.120 13.700 103.600 ;
        RECT 2906.300 103.120 2914.100 103.600 ;
        RECT 5.520 97.680 13.700 98.160 ;
        RECT 2906.300 97.680 2914.100 98.160 ;
        RECT 5.520 92.240 13.700 92.720 ;
        RECT 2906.300 92.240 2914.100 92.720 ;
        RECT 5.520 86.800 13.700 87.280 ;
        RECT 2906.300 86.800 2914.100 87.280 ;
        RECT 5.520 81.360 13.700 81.840 ;
        RECT 2906.300 81.360 2914.100 81.840 ;
        RECT 5.520 75.920 13.700 76.400 ;
        RECT 2906.300 75.920 2914.100 76.400 ;
        RECT 5.520 70.480 13.700 70.960 ;
        RECT 2906.300 70.480 2914.100 70.960 ;
        RECT 5.520 65.040 13.700 65.520 ;
        RECT 2906.300 65.040 2914.100 65.520 ;
        RECT 5.520 59.600 13.700 60.080 ;
        RECT 2906.300 59.600 2914.100 60.080 ;
        RECT 5.520 54.160 13.700 54.640 ;
        RECT 2906.300 54.160 2914.100 54.640 ;
        RECT 5.520 48.720 13.700 49.200 ;
        RECT 2906.300 48.720 2914.100 49.200 ;
        RECT 5.520 43.280 13.700 43.760 ;
        RECT 2906.300 43.280 2914.100 43.760 ;
        RECT 5.520 37.840 13.700 38.320 ;
        RECT 2906.300 37.840 2914.100 38.320 ;
        RECT 5.520 32.400 13.700 32.880 ;
        RECT 2906.300 32.400 2914.100 32.880 ;
        RECT 5.520 26.960 13.700 27.440 ;
        RECT 2906.300 26.960 2914.100 27.440 ;
        RECT 5.520 21.520 13.700 22.000 ;
        RECT 2906.300 21.520 2914.100 22.000 ;
        RECT 5.520 16.080 13.700 16.560 ;
        RECT 2906.300 16.080 2914.100 16.560 ;
        RECT 5.520 10.640 2914.100 11.120 ;
      LAYER via ;
        RECT 94.110 3508.670 94.370 3508.930 ;
        RECT 94.430 3508.670 94.690 3508.930 ;
        RECT 94.750 3508.670 95.010 3508.930 ;
        RECT 95.070 3508.670 95.330 3508.930 ;
        RECT 95.390 3508.670 95.650 3508.930 ;
        RECT 95.710 3508.670 95.970 3508.930 ;
        RECT 96.030 3508.670 96.290 3508.930 ;
        RECT 96.350 3508.670 96.610 3508.930 ;
        RECT 96.670 3508.670 96.930 3508.930 ;
        RECT 184.110 3508.670 184.370 3508.930 ;
        RECT 184.430 3508.670 184.690 3508.930 ;
        RECT 184.750 3508.670 185.010 3508.930 ;
        RECT 185.070 3508.670 185.330 3508.930 ;
        RECT 185.390 3508.670 185.650 3508.930 ;
        RECT 185.710 3508.670 185.970 3508.930 ;
        RECT 186.030 3508.670 186.290 3508.930 ;
        RECT 186.350 3508.670 186.610 3508.930 ;
        RECT 186.670 3508.670 186.930 3508.930 ;
        RECT 274.110 3508.670 274.370 3508.930 ;
        RECT 274.430 3508.670 274.690 3508.930 ;
        RECT 274.750 3508.670 275.010 3508.930 ;
        RECT 275.070 3508.670 275.330 3508.930 ;
        RECT 275.390 3508.670 275.650 3508.930 ;
        RECT 275.710 3508.670 275.970 3508.930 ;
        RECT 276.030 3508.670 276.290 3508.930 ;
        RECT 276.350 3508.670 276.610 3508.930 ;
        RECT 276.670 3508.670 276.930 3508.930 ;
        RECT 364.110 3508.670 364.370 3508.930 ;
        RECT 364.430 3508.670 364.690 3508.930 ;
        RECT 364.750 3508.670 365.010 3508.930 ;
        RECT 365.070 3508.670 365.330 3508.930 ;
        RECT 365.390 3508.670 365.650 3508.930 ;
        RECT 365.710 3508.670 365.970 3508.930 ;
        RECT 366.030 3508.670 366.290 3508.930 ;
        RECT 366.350 3508.670 366.610 3508.930 ;
        RECT 366.670 3508.670 366.930 3508.930 ;
        RECT 454.110 3508.670 454.370 3508.930 ;
        RECT 454.430 3508.670 454.690 3508.930 ;
        RECT 454.750 3508.670 455.010 3508.930 ;
        RECT 455.070 3508.670 455.330 3508.930 ;
        RECT 455.390 3508.670 455.650 3508.930 ;
        RECT 455.710 3508.670 455.970 3508.930 ;
        RECT 456.030 3508.670 456.290 3508.930 ;
        RECT 456.350 3508.670 456.610 3508.930 ;
        RECT 456.670 3508.670 456.930 3508.930 ;
        RECT 544.110 3508.670 544.370 3508.930 ;
        RECT 544.430 3508.670 544.690 3508.930 ;
        RECT 544.750 3508.670 545.010 3508.930 ;
        RECT 545.070 3508.670 545.330 3508.930 ;
        RECT 545.390 3508.670 545.650 3508.930 ;
        RECT 545.710 3508.670 545.970 3508.930 ;
        RECT 546.030 3508.670 546.290 3508.930 ;
        RECT 546.350 3508.670 546.610 3508.930 ;
        RECT 546.670 3508.670 546.930 3508.930 ;
        RECT 634.110 3508.670 634.370 3508.930 ;
        RECT 634.430 3508.670 634.690 3508.930 ;
        RECT 634.750 3508.670 635.010 3508.930 ;
        RECT 635.070 3508.670 635.330 3508.930 ;
        RECT 635.390 3508.670 635.650 3508.930 ;
        RECT 635.710 3508.670 635.970 3508.930 ;
        RECT 636.030 3508.670 636.290 3508.930 ;
        RECT 636.350 3508.670 636.610 3508.930 ;
        RECT 636.670 3508.670 636.930 3508.930 ;
        RECT 724.110 3508.670 724.370 3508.930 ;
        RECT 724.430 3508.670 724.690 3508.930 ;
        RECT 724.750 3508.670 725.010 3508.930 ;
        RECT 725.070 3508.670 725.330 3508.930 ;
        RECT 725.390 3508.670 725.650 3508.930 ;
        RECT 725.710 3508.670 725.970 3508.930 ;
        RECT 726.030 3508.670 726.290 3508.930 ;
        RECT 726.350 3508.670 726.610 3508.930 ;
        RECT 726.670 3508.670 726.930 3508.930 ;
        RECT 814.110 3508.670 814.370 3508.930 ;
        RECT 814.430 3508.670 814.690 3508.930 ;
        RECT 814.750 3508.670 815.010 3508.930 ;
        RECT 815.070 3508.670 815.330 3508.930 ;
        RECT 815.390 3508.670 815.650 3508.930 ;
        RECT 815.710 3508.670 815.970 3508.930 ;
        RECT 816.030 3508.670 816.290 3508.930 ;
        RECT 816.350 3508.670 816.610 3508.930 ;
        RECT 816.670 3508.670 816.930 3508.930 ;
        RECT 904.110 3508.670 904.370 3508.930 ;
        RECT 904.430 3508.670 904.690 3508.930 ;
        RECT 904.750 3508.670 905.010 3508.930 ;
        RECT 905.070 3508.670 905.330 3508.930 ;
        RECT 905.390 3508.670 905.650 3508.930 ;
        RECT 905.710 3508.670 905.970 3508.930 ;
        RECT 906.030 3508.670 906.290 3508.930 ;
        RECT 906.350 3508.670 906.610 3508.930 ;
        RECT 906.670 3508.670 906.930 3508.930 ;
        RECT 994.110 3508.670 994.370 3508.930 ;
        RECT 994.430 3508.670 994.690 3508.930 ;
        RECT 994.750 3508.670 995.010 3508.930 ;
        RECT 995.070 3508.670 995.330 3508.930 ;
        RECT 995.390 3508.670 995.650 3508.930 ;
        RECT 995.710 3508.670 995.970 3508.930 ;
        RECT 996.030 3508.670 996.290 3508.930 ;
        RECT 996.350 3508.670 996.610 3508.930 ;
        RECT 996.670 3508.670 996.930 3508.930 ;
        RECT 1084.110 3508.670 1084.370 3508.930 ;
        RECT 1084.430 3508.670 1084.690 3508.930 ;
        RECT 1084.750 3508.670 1085.010 3508.930 ;
        RECT 1085.070 3508.670 1085.330 3508.930 ;
        RECT 1085.390 3508.670 1085.650 3508.930 ;
        RECT 1085.710 3508.670 1085.970 3508.930 ;
        RECT 1086.030 3508.670 1086.290 3508.930 ;
        RECT 1086.350 3508.670 1086.610 3508.930 ;
        RECT 1086.670 3508.670 1086.930 3508.930 ;
        RECT 1174.110 3508.670 1174.370 3508.930 ;
        RECT 1174.430 3508.670 1174.690 3508.930 ;
        RECT 1174.750 3508.670 1175.010 3508.930 ;
        RECT 1175.070 3508.670 1175.330 3508.930 ;
        RECT 1175.390 3508.670 1175.650 3508.930 ;
        RECT 1175.710 3508.670 1175.970 3508.930 ;
        RECT 1176.030 3508.670 1176.290 3508.930 ;
        RECT 1176.350 3508.670 1176.610 3508.930 ;
        RECT 1176.670 3508.670 1176.930 3508.930 ;
        RECT 1264.110 3508.670 1264.370 3508.930 ;
        RECT 1264.430 3508.670 1264.690 3508.930 ;
        RECT 1264.750 3508.670 1265.010 3508.930 ;
        RECT 1265.070 3508.670 1265.330 3508.930 ;
        RECT 1265.390 3508.670 1265.650 3508.930 ;
        RECT 1265.710 3508.670 1265.970 3508.930 ;
        RECT 1266.030 3508.670 1266.290 3508.930 ;
        RECT 1266.350 3508.670 1266.610 3508.930 ;
        RECT 1266.670 3508.670 1266.930 3508.930 ;
        RECT 1354.110 3508.670 1354.370 3508.930 ;
        RECT 1354.430 3508.670 1354.690 3508.930 ;
        RECT 1354.750 3508.670 1355.010 3508.930 ;
        RECT 1355.070 3508.670 1355.330 3508.930 ;
        RECT 1355.390 3508.670 1355.650 3508.930 ;
        RECT 1355.710 3508.670 1355.970 3508.930 ;
        RECT 1356.030 3508.670 1356.290 3508.930 ;
        RECT 1356.350 3508.670 1356.610 3508.930 ;
        RECT 1356.670 3508.670 1356.930 3508.930 ;
        RECT 1444.110 3508.670 1444.370 3508.930 ;
        RECT 1444.430 3508.670 1444.690 3508.930 ;
        RECT 1444.750 3508.670 1445.010 3508.930 ;
        RECT 1445.070 3508.670 1445.330 3508.930 ;
        RECT 1445.390 3508.670 1445.650 3508.930 ;
        RECT 1445.710 3508.670 1445.970 3508.930 ;
        RECT 1446.030 3508.670 1446.290 3508.930 ;
        RECT 1446.350 3508.670 1446.610 3508.930 ;
        RECT 1446.670 3508.670 1446.930 3508.930 ;
        RECT 1534.110 3508.670 1534.370 3508.930 ;
        RECT 1534.430 3508.670 1534.690 3508.930 ;
        RECT 1534.750 3508.670 1535.010 3508.930 ;
        RECT 1535.070 3508.670 1535.330 3508.930 ;
        RECT 1535.390 3508.670 1535.650 3508.930 ;
        RECT 1535.710 3508.670 1535.970 3508.930 ;
        RECT 1536.030 3508.670 1536.290 3508.930 ;
        RECT 1536.350 3508.670 1536.610 3508.930 ;
        RECT 1536.670 3508.670 1536.930 3508.930 ;
        RECT 1624.110 3508.670 1624.370 3508.930 ;
        RECT 1624.430 3508.670 1624.690 3508.930 ;
        RECT 1624.750 3508.670 1625.010 3508.930 ;
        RECT 1625.070 3508.670 1625.330 3508.930 ;
        RECT 1625.390 3508.670 1625.650 3508.930 ;
        RECT 1625.710 3508.670 1625.970 3508.930 ;
        RECT 1626.030 3508.670 1626.290 3508.930 ;
        RECT 1626.350 3508.670 1626.610 3508.930 ;
        RECT 1626.670 3508.670 1626.930 3508.930 ;
        RECT 1714.110 3508.670 1714.370 3508.930 ;
        RECT 1714.430 3508.670 1714.690 3508.930 ;
        RECT 1714.750 3508.670 1715.010 3508.930 ;
        RECT 1715.070 3508.670 1715.330 3508.930 ;
        RECT 1715.390 3508.670 1715.650 3508.930 ;
        RECT 1715.710 3508.670 1715.970 3508.930 ;
        RECT 1716.030 3508.670 1716.290 3508.930 ;
        RECT 1716.350 3508.670 1716.610 3508.930 ;
        RECT 1716.670 3508.670 1716.930 3508.930 ;
        RECT 1804.110 3508.670 1804.370 3508.930 ;
        RECT 1804.430 3508.670 1804.690 3508.930 ;
        RECT 1804.750 3508.670 1805.010 3508.930 ;
        RECT 1805.070 3508.670 1805.330 3508.930 ;
        RECT 1805.390 3508.670 1805.650 3508.930 ;
        RECT 1805.710 3508.670 1805.970 3508.930 ;
        RECT 1806.030 3508.670 1806.290 3508.930 ;
        RECT 1806.350 3508.670 1806.610 3508.930 ;
        RECT 1806.670 3508.670 1806.930 3508.930 ;
        RECT 1894.110 3508.670 1894.370 3508.930 ;
        RECT 1894.430 3508.670 1894.690 3508.930 ;
        RECT 1894.750 3508.670 1895.010 3508.930 ;
        RECT 1895.070 3508.670 1895.330 3508.930 ;
        RECT 1895.390 3508.670 1895.650 3508.930 ;
        RECT 1895.710 3508.670 1895.970 3508.930 ;
        RECT 1896.030 3508.670 1896.290 3508.930 ;
        RECT 1896.350 3508.670 1896.610 3508.930 ;
        RECT 1896.670 3508.670 1896.930 3508.930 ;
        RECT 1984.110 3508.670 1984.370 3508.930 ;
        RECT 1984.430 3508.670 1984.690 3508.930 ;
        RECT 1984.750 3508.670 1985.010 3508.930 ;
        RECT 1985.070 3508.670 1985.330 3508.930 ;
        RECT 1985.390 3508.670 1985.650 3508.930 ;
        RECT 1985.710 3508.670 1985.970 3508.930 ;
        RECT 1986.030 3508.670 1986.290 3508.930 ;
        RECT 1986.350 3508.670 1986.610 3508.930 ;
        RECT 1986.670 3508.670 1986.930 3508.930 ;
        RECT 2074.110 3508.670 2074.370 3508.930 ;
        RECT 2074.430 3508.670 2074.690 3508.930 ;
        RECT 2074.750 3508.670 2075.010 3508.930 ;
        RECT 2075.070 3508.670 2075.330 3508.930 ;
        RECT 2075.390 3508.670 2075.650 3508.930 ;
        RECT 2075.710 3508.670 2075.970 3508.930 ;
        RECT 2076.030 3508.670 2076.290 3508.930 ;
        RECT 2076.350 3508.670 2076.610 3508.930 ;
        RECT 2076.670 3508.670 2076.930 3508.930 ;
        RECT 2164.110 3508.670 2164.370 3508.930 ;
        RECT 2164.430 3508.670 2164.690 3508.930 ;
        RECT 2164.750 3508.670 2165.010 3508.930 ;
        RECT 2165.070 3508.670 2165.330 3508.930 ;
        RECT 2165.390 3508.670 2165.650 3508.930 ;
        RECT 2165.710 3508.670 2165.970 3508.930 ;
        RECT 2166.030 3508.670 2166.290 3508.930 ;
        RECT 2166.350 3508.670 2166.610 3508.930 ;
        RECT 2166.670 3508.670 2166.930 3508.930 ;
        RECT 2254.110 3508.670 2254.370 3508.930 ;
        RECT 2254.430 3508.670 2254.690 3508.930 ;
        RECT 2254.750 3508.670 2255.010 3508.930 ;
        RECT 2255.070 3508.670 2255.330 3508.930 ;
        RECT 2255.390 3508.670 2255.650 3508.930 ;
        RECT 2255.710 3508.670 2255.970 3508.930 ;
        RECT 2256.030 3508.670 2256.290 3508.930 ;
        RECT 2256.350 3508.670 2256.610 3508.930 ;
        RECT 2256.670 3508.670 2256.930 3508.930 ;
        RECT 2344.110 3508.670 2344.370 3508.930 ;
        RECT 2344.430 3508.670 2344.690 3508.930 ;
        RECT 2344.750 3508.670 2345.010 3508.930 ;
        RECT 2345.070 3508.670 2345.330 3508.930 ;
        RECT 2345.390 3508.670 2345.650 3508.930 ;
        RECT 2345.710 3508.670 2345.970 3508.930 ;
        RECT 2346.030 3508.670 2346.290 3508.930 ;
        RECT 2346.350 3508.670 2346.610 3508.930 ;
        RECT 2346.670 3508.670 2346.930 3508.930 ;
        RECT 2434.110 3508.670 2434.370 3508.930 ;
        RECT 2434.430 3508.670 2434.690 3508.930 ;
        RECT 2434.750 3508.670 2435.010 3508.930 ;
        RECT 2435.070 3508.670 2435.330 3508.930 ;
        RECT 2435.390 3508.670 2435.650 3508.930 ;
        RECT 2435.710 3508.670 2435.970 3508.930 ;
        RECT 2436.030 3508.670 2436.290 3508.930 ;
        RECT 2436.350 3508.670 2436.610 3508.930 ;
        RECT 2436.670 3508.670 2436.930 3508.930 ;
        RECT 2524.110 3508.670 2524.370 3508.930 ;
        RECT 2524.430 3508.670 2524.690 3508.930 ;
        RECT 2524.750 3508.670 2525.010 3508.930 ;
        RECT 2525.070 3508.670 2525.330 3508.930 ;
        RECT 2525.390 3508.670 2525.650 3508.930 ;
        RECT 2525.710 3508.670 2525.970 3508.930 ;
        RECT 2526.030 3508.670 2526.290 3508.930 ;
        RECT 2526.350 3508.670 2526.610 3508.930 ;
        RECT 2526.670 3508.670 2526.930 3508.930 ;
        RECT 2614.110 3508.670 2614.370 3508.930 ;
        RECT 2614.430 3508.670 2614.690 3508.930 ;
        RECT 2614.750 3508.670 2615.010 3508.930 ;
        RECT 2615.070 3508.670 2615.330 3508.930 ;
        RECT 2615.390 3508.670 2615.650 3508.930 ;
        RECT 2615.710 3508.670 2615.970 3508.930 ;
        RECT 2616.030 3508.670 2616.290 3508.930 ;
        RECT 2616.350 3508.670 2616.610 3508.930 ;
        RECT 2616.670 3508.670 2616.930 3508.930 ;
        RECT 2704.110 3508.670 2704.370 3508.930 ;
        RECT 2704.430 3508.670 2704.690 3508.930 ;
        RECT 2704.750 3508.670 2705.010 3508.930 ;
        RECT 2705.070 3508.670 2705.330 3508.930 ;
        RECT 2705.390 3508.670 2705.650 3508.930 ;
        RECT 2705.710 3508.670 2705.970 3508.930 ;
        RECT 2706.030 3508.670 2706.290 3508.930 ;
        RECT 2706.350 3508.670 2706.610 3508.930 ;
        RECT 2706.670 3508.670 2706.930 3508.930 ;
        RECT 2794.110 3508.670 2794.370 3508.930 ;
        RECT 2794.430 3508.670 2794.690 3508.930 ;
        RECT 2794.750 3508.670 2795.010 3508.930 ;
        RECT 2795.070 3508.670 2795.330 3508.930 ;
        RECT 2795.390 3508.670 2795.650 3508.930 ;
        RECT 2795.710 3508.670 2795.970 3508.930 ;
        RECT 2796.030 3508.670 2796.290 3508.930 ;
        RECT 2796.350 3508.670 2796.610 3508.930 ;
        RECT 2796.670 3508.670 2796.930 3508.930 ;
        RECT 2884.110 3508.670 2884.370 3508.930 ;
        RECT 2884.430 3508.670 2884.690 3508.930 ;
        RECT 2884.750 3508.670 2885.010 3508.930 ;
        RECT 2885.070 3508.670 2885.330 3508.930 ;
        RECT 2885.390 3508.670 2885.650 3508.930 ;
        RECT 2885.710 3508.670 2885.970 3508.930 ;
        RECT 2886.030 3508.670 2886.290 3508.930 ;
        RECT 2886.350 3508.670 2886.610 3508.930 ;
        RECT 2886.670 3508.670 2886.930 3508.930 ;
        RECT 94.110 10.750 94.370 11.010 ;
        RECT 94.430 10.750 94.690 11.010 ;
        RECT 94.750 10.750 95.010 11.010 ;
        RECT 95.070 10.750 95.330 11.010 ;
        RECT 95.390 10.750 95.650 11.010 ;
        RECT 95.710 10.750 95.970 11.010 ;
        RECT 96.030 10.750 96.290 11.010 ;
        RECT 96.350 10.750 96.610 11.010 ;
        RECT 96.670 10.750 96.930 11.010 ;
        RECT 184.110 10.750 184.370 11.010 ;
        RECT 184.430 10.750 184.690 11.010 ;
        RECT 184.750 10.750 185.010 11.010 ;
        RECT 185.070 10.750 185.330 11.010 ;
        RECT 185.390 10.750 185.650 11.010 ;
        RECT 185.710 10.750 185.970 11.010 ;
        RECT 186.030 10.750 186.290 11.010 ;
        RECT 186.350 10.750 186.610 11.010 ;
        RECT 186.670 10.750 186.930 11.010 ;
        RECT 274.110 10.750 274.370 11.010 ;
        RECT 274.430 10.750 274.690 11.010 ;
        RECT 274.750 10.750 275.010 11.010 ;
        RECT 275.070 10.750 275.330 11.010 ;
        RECT 275.390 10.750 275.650 11.010 ;
        RECT 275.710 10.750 275.970 11.010 ;
        RECT 276.030 10.750 276.290 11.010 ;
        RECT 276.350 10.750 276.610 11.010 ;
        RECT 276.670 10.750 276.930 11.010 ;
        RECT 364.110 10.750 364.370 11.010 ;
        RECT 364.430 10.750 364.690 11.010 ;
        RECT 364.750 10.750 365.010 11.010 ;
        RECT 365.070 10.750 365.330 11.010 ;
        RECT 365.390 10.750 365.650 11.010 ;
        RECT 365.710 10.750 365.970 11.010 ;
        RECT 366.030 10.750 366.290 11.010 ;
        RECT 366.350 10.750 366.610 11.010 ;
        RECT 366.670 10.750 366.930 11.010 ;
        RECT 454.110 10.750 454.370 11.010 ;
        RECT 454.430 10.750 454.690 11.010 ;
        RECT 454.750 10.750 455.010 11.010 ;
        RECT 455.070 10.750 455.330 11.010 ;
        RECT 455.390 10.750 455.650 11.010 ;
        RECT 455.710 10.750 455.970 11.010 ;
        RECT 456.030 10.750 456.290 11.010 ;
        RECT 456.350 10.750 456.610 11.010 ;
        RECT 456.670 10.750 456.930 11.010 ;
        RECT 544.110 10.750 544.370 11.010 ;
        RECT 544.430 10.750 544.690 11.010 ;
        RECT 544.750 10.750 545.010 11.010 ;
        RECT 545.070 10.750 545.330 11.010 ;
        RECT 545.390 10.750 545.650 11.010 ;
        RECT 545.710 10.750 545.970 11.010 ;
        RECT 546.030 10.750 546.290 11.010 ;
        RECT 546.350 10.750 546.610 11.010 ;
        RECT 546.670 10.750 546.930 11.010 ;
        RECT 634.110 10.750 634.370 11.010 ;
        RECT 634.430 10.750 634.690 11.010 ;
        RECT 634.750 10.750 635.010 11.010 ;
        RECT 635.070 10.750 635.330 11.010 ;
        RECT 635.390 10.750 635.650 11.010 ;
        RECT 635.710 10.750 635.970 11.010 ;
        RECT 636.030 10.750 636.290 11.010 ;
        RECT 636.350 10.750 636.610 11.010 ;
        RECT 636.670 10.750 636.930 11.010 ;
        RECT 724.110 10.750 724.370 11.010 ;
        RECT 724.430 10.750 724.690 11.010 ;
        RECT 724.750 10.750 725.010 11.010 ;
        RECT 725.070 10.750 725.330 11.010 ;
        RECT 725.390 10.750 725.650 11.010 ;
        RECT 725.710 10.750 725.970 11.010 ;
        RECT 726.030 10.750 726.290 11.010 ;
        RECT 726.350 10.750 726.610 11.010 ;
        RECT 726.670 10.750 726.930 11.010 ;
        RECT 814.110 10.750 814.370 11.010 ;
        RECT 814.430 10.750 814.690 11.010 ;
        RECT 814.750 10.750 815.010 11.010 ;
        RECT 815.070 10.750 815.330 11.010 ;
        RECT 815.390 10.750 815.650 11.010 ;
        RECT 815.710 10.750 815.970 11.010 ;
        RECT 816.030 10.750 816.290 11.010 ;
        RECT 816.350 10.750 816.610 11.010 ;
        RECT 816.670 10.750 816.930 11.010 ;
        RECT 904.110 10.750 904.370 11.010 ;
        RECT 904.430 10.750 904.690 11.010 ;
        RECT 904.750 10.750 905.010 11.010 ;
        RECT 905.070 10.750 905.330 11.010 ;
        RECT 905.390 10.750 905.650 11.010 ;
        RECT 905.710 10.750 905.970 11.010 ;
        RECT 906.030 10.750 906.290 11.010 ;
        RECT 906.350 10.750 906.610 11.010 ;
        RECT 906.670 10.750 906.930 11.010 ;
        RECT 994.110 10.750 994.370 11.010 ;
        RECT 994.430 10.750 994.690 11.010 ;
        RECT 994.750 10.750 995.010 11.010 ;
        RECT 995.070 10.750 995.330 11.010 ;
        RECT 995.390 10.750 995.650 11.010 ;
        RECT 995.710 10.750 995.970 11.010 ;
        RECT 996.030 10.750 996.290 11.010 ;
        RECT 996.350 10.750 996.610 11.010 ;
        RECT 996.670 10.750 996.930 11.010 ;
        RECT 1084.110 10.750 1084.370 11.010 ;
        RECT 1084.430 10.750 1084.690 11.010 ;
        RECT 1084.750 10.750 1085.010 11.010 ;
        RECT 1085.070 10.750 1085.330 11.010 ;
        RECT 1085.390 10.750 1085.650 11.010 ;
        RECT 1085.710 10.750 1085.970 11.010 ;
        RECT 1086.030 10.750 1086.290 11.010 ;
        RECT 1086.350 10.750 1086.610 11.010 ;
        RECT 1086.670 10.750 1086.930 11.010 ;
        RECT 1174.110 10.750 1174.370 11.010 ;
        RECT 1174.430 10.750 1174.690 11.010 ;
        RECT 1174.750 10.750 1175.010 11.010 ;
        RECT 1175.070 10.750 1175.330 11.010 ;
        RECT 1175.390 10.750 1175.650 11.010 ;
        RECT 1175.710 10.750 1175.970 11.010 ;
        RECT 1176.030 10.750 1176.290 11.010 ;
        RECT 1176.350 10.750 1176.610 11.010 ;
        RECT 1176.670 10.750 1176.930 11.010 ;
        RECT 1264.110 10.750 1264.370 11.010 ;
        RECT 1264.430 10.750 1264.690 11.010 ;
        RECT 1264.750 10.750 1265.010 11.010 ;
        RECT 1265.070 10.750 1265.330 11.010 ;
        RECT 1265.390 10.750 1265.650 11.010 ;
        RECT 1265.710 10.750 1265.970 11.010 ;
        RECT 1266.030 10.750 1266.290 11.010 ;
        RECT 1266.350 10.750 1266.610 11.010 ;
        RECT 1266.670 10.750 1266.930 11.010 ;
        RECT 1354.110 10.750 1354.370 11.010 ;
        RECT 1354.430 10.750 1354.690 11.010 ;
        RECT 1354.750 10.750 1355.010 11.010 ;
        RECT 1355.070 10.750 1355.330 11.010 ;
        RECT 1355.390 10.750 1355.650 11.010 ;
        RECT 1355.710 10.750 1355.970 11.010 ;
        RECT 1356.030 10.750 1356.290 11.010 ;
        RECT 1356.350 10.750 1356.610 11.010 ;
        RECT 1356.670 10.750 1356.930 11.010 ;
        RECT 1444.110 10.750 1444.370 11.010 ;
        RECT 1444.430 10.750 1444.690 11.010 ;
        RECT 1444.750 10.750 1445.010 11.010 ;
        RECT 1445.070 10.750 1445.330 11.010 ;
        RECT 1445.390 10.750 1445.650 11.010 ;
        RECT 1445.710 10.750 1445.970 11.010 ;
        RECT 1446.030 10.750 1446.290 11.010 ;
        RECT 1446.350 10.750 1446.610 11.010 ;
        RECT 1446.670 10.750 1446.930 11.010 ;
        RECT 1534.110 10.750 1534.370 11.010 ;
        RECT 1534.430 10.750 1534.690 11.010 ;
        RECT 1534.750 10.750 1535.010 11.010 ;
        RECT 1535.070 10.750 1535.330 11.010 ;
        RECT 1535.390 10.750 1535.650 11.010 ;
        RECT 1535.710 10.750 1535.970 11.010 ;
        RECT 1536.030 10.750 1536.290 11.010 ;
        RECT 1536.350 10.750 1536.610 11.010 ;
        RECT 1536.670 10.750 1536.930 11.010 ;
        RECT 1624.110 10.750 1624.370 11.010 ;
        RECT 1624.430 10.750 1624.690 11.010 ;
        RECT 1624.750 10.750 1625.010 11.010 ;
        RECT 1625.070 10.750 1625.330 11.010 ;
        RECT 1625.390 10.750 1625.650 11.010 ;
        RECT 1625.710 10.750 1625.970 11.010 ;
        RECT 1626.030 10.750 1626.290 11.010 ;
        RECT 1626.350 10.750 1626.610 11.010 ;
        RECT 1626.670 10.750 1626.930 11.010 ;
        RECT 1714.110 10.750 1714.370 11.010 ;
        RECT 1714.430 10.750 1714.690 11.010 ;
        RECT 1714.750 10.750 1715.010 11.010 ;
        RECT 1715.070 10.750 1715.330 11.010 ;
        RECT 1715.390 10.750 1715.650 11.010 ;
        RECT 1715.710 10.750 1715.970 11.010 ;
        RECT 1716.030 10.750 1716.290 11.010 ;
        RECT 1716.350 10.750 1716.610 11.010 ;
        RECT 1716.670 10.750 1716.930 11.010 ;
        RECT 1804.110 10.750 1804.370 11.010 ;
        RECT 1804.430 10.750 1804.690 11.010 ;
        RECT 1804.750 10.750 1805.010 11.010 ;
        RECT 1805.070 10.750 1805.330 11.010 ;
        RECT 1805.390 10.750 1805.650 11.010 ;
        RECT 1805.710 10.750 1805.970 11.010 ;
        RECT 1806.030 10.750 1806.290 11.010 ;
        RECT 1806.350 10.750 1806.610 11.010 ;
        RECT 1806.670 10.750 1806.930 11.010 ;
        RECT 1894.110 10.750 1894.370 11.010 ;
        RECT 1894.430 10.750 1894.690 11.010 ;
        RECT 1894.750 10.750 1895.010 11.010 ;
        RECT 1895.070 10.750 1895.330 11.010 ;
        RECT 1895.390 10.750 1895.650 11.010 ;
        RECT 1895.710 10.750 1895.970 11.010 ;
        RECT 1896.030 10.750 1896.290 11.010 ;
        RECT 1896.350 10.750 1896.610 11.010 ;
        RECT 1896.670 10.750 1896.930 11.010 ;
        RECT 1984.110 10.750 1984.370 11.010 ;
        RECT 1984.430 10.750 1984.690 11.010 ;
        RECT 1984.750 10.750 1985.010 11.010 ;
        RECT 1985.070 10.750 1985.330 11.010 ;
        RECT 1985.390 10.750 1985.650 11.010 ;
        RECT 1985.710 10.750 1985.970 11.010 ;
        RECT 1986.030 10.750 1986.290 11.010 ;
        RECT 1986.350 10.750 1986.610 11.010 ;
        RECT 1986.670 10.750 1986.930 11.010 ;
        RECT 2074.110 10.750 2074.370 11.010 ;
        RECT 2074.430 10.750 2074.690 11.010 ;
        RECT 2074.750 10.750 2075.010 11.010 ;
        RECT 2075.070 10.750 2075.330 11.010 ;
        RECT 2075.390 10.750 2075.650 11.010 ;
        RECT 2075.710 10.750 2075.970 11.010 ;
        RECT 2076.030 10.750 2076.290 11.010 ;
        RECT 2076.350 10.750 2076.610 11.010 ;
        RECT 2076.670 10.750 2076.930 11.010 ;
        RECT 2164.110 10.750 2164.370 11.010 ;
        RECT 2164.430 10.750 2164.690 11.010 ;
        RECT 2164.750 10.750 2165.010 11.010 ;
        RECT 2165.070 10.750 2165.330 11.010 ;
        RECT 2165.390 10.750 2165.650 11.010 ;
        RECT 2165.710 10.750 2165.970 11.010 ;
        RECT 2166.030 10.750 2166.290 11.010 ;
        RECT 2166.350 10.750 2166.610 11.010 ;
        RECT 2166.670 10.750 2166.930 11.010 ;
        RECT 2254.110 10.750 2254.370 11.010 ;
        RECT 2254.430 10.750 2254.690 11.010 ;
        RECT 2254.750 10.750 2255.010 11.010 ;
        RECT 2255.070 10.750 2255.330 11.010 ;
        RECT 2255.390 10.750 2255.650 11.010 ;
        RECT 2255.710 10.750 2255.970 11.010 ;
        RECT 2256.030 10.750 2256.290 11.010 ;
        RECT 2256.350 10.750 2256.610 11.010 ;
        RECT 2256.670 10.750 2256.930 11.010 ;
        RECT 2344.110 10.750 2344.370 11.010 ;
        RECT 2344.430 10.750 2344.690 11.010 ;
        RECT 2344.750 10.750 2345.010 11.010 ;
        RECT 2345.070 10.750 2345.330 11.010 ;
        RECT 2345.390 10.750 2345.650 11.010 ;
        RECT 2345.710 10.750 2345.970 11.010 ;
        RECT 2346.030 10.750 2346.290 11.010 ;
        RECT 2346.350 10.750 2346.610 11.010 ;
        RECT 2346.670 10.750 2346.930 11.010 ;
        RECT 2434.110 10.750 2434.370 11.010 ;
        RECT 2434.430 10.750 2434.690 11.010 ;
        RECT 2434.750 10.750 2435.010 11.010 ;
        RECT 2435.070 10.750 2435.330 11.010 ;
        RECT 2435.390 10.750 2435.650 11.010 ;
        RECT 2435.710 10.750 2435.970 11.010 ;
        RECT 2436.030 10.750 2436.290 11.010 ;
        RECT 2436.350 10.750 2436.610 11.010 ;
        RECT 2436.670 10.750 2436.930 11.010 ;
        RECT 2524.110 10.750 2524.370 11.010 ;
        RECT 2524.430 10.750 2524.690 11.010 ;
        RECT 2524.750 10.750 2525.010 11.010 ;
        RECT 2525.070 10.750 2525.330 11.010 ;
        RECT 2525.390 10.750 2525.650 11.010 ;
        RECT 2525.710 10.750 2525.970 11.010 ;
        RECT 2526.030 10.750 2526.290 11.010 ;
        RECT 2526.350 10.750 2526.610 11.010 ;
        RECT 2526.670 10.750 2526.930 11.010 ;
        RECT 2614.110 10.750 2614.370 11.010 ;
        RECT 2614.430 10.750 2614.690 11.010 ;
        RECT 2614.750 10.750 2615.010 11.010 ;
        RECT 2615.070 10.750 2615.330 11.010 ;
        RECT 2615.390 10.750 2615.650 11.010 ;
        RECT 2615.710 10.750 2615.970 11.010 ;
        RECT 2616.030 10.750 2616.290 11.010 ;
        RECT 2616.350 10.750 2616.610 11.010 ;
        RECT 2616.670 10.750 2616.930 11.010 ;
        RECT 2704.110 10.750 2704.370 11.010 ;
        RECT 2704.430 10.750 2704.690 11.010 ;
        RECT 2704.750 10.750 2705.010 11.010 ;
        RECT 2705.070 10.750 2705.330 11.010 ;
        RECT 2705.390 10.750 2705.650 11.010 ;
        RECT 2705.710 10.750 2705.970 11.010 ;
        RECT 2706.030 10.750 2706.290 11.010 ;
        RECT 2706.350 10.750 2706.610 11.010 ;
        RECT 2706.670 10.750 2706.930 11.010 ;
        RECT 2794.110 10.750 2794.370 11.010 ;
        RECT 2794.430 10.750 2794.690 11.010 ;
        RECT 2794.750 10.750 2795.010 11.010 ;
        RECT 2795.070 10.750 2795.330 11.010 ;
        RECT 2795.390 10.750 2795.650 11.010 ;
        RECT 2795.710 10.750 2795.970 11.010 ;
        RECT 2796.030 10.750 2796.290 11.010 ;
        RECT 2796.350 10.750 2796.610 11.010 ;
        RECT 2796.670 10.750 2796.930 11.010 ;
        RECT 2884.110 10.750 2884.370 11.010 ;
        RECT 2884.430 10.750 2884.690 11.010 ;
        RECT 2884.750 10.750 2885.010 11.010 ;
        RECT 2885.070 10.750 2885.330 11.010 ;
        RECT 2885.390 10.750 2885.650 11.010 ;
        RECT 2885.710 10.750 2885.970 11.010 ;
        RECT 2886.030 10.750 2886.290 11.010 ;
        RECT 2886.350 10.750 2886.610 11.010 ;
        RECT 2886.670 10.750 2886.930 11.010 ;
      LAYER met2 ;
        RECT 94.110 3508.560 96.930 3509.040 ;
        RECT 184.110 3508.560 186.930 3509.040 ;
        RECT 274.110 3508.560 276.930 3509.040 ;
        RECT 364.110 3508.560 366.930 3509.040 ;
        RECT 454.110 3508.560 456.930 3509.040 ;
        RECT 544.110 3508.560 546.930 3509.040 ;
        RECT 634.110 3508.560 636.930 3509.040 ;
        RECT 724.110 3508.560 726.930 3509.040 ;
        RECT 814.110 3508.560 816.930 3509.040 ;
        RECT 904.110 3508.560 906.930 3509.040 ;
        RECT 994.110 3508.560 996.930 3509.040 ;
        RECT 1084.110 3508.560 1086.930 3509.040 ;
        RECT 1174.110 3508.560 1176.930 3509.040 ;
        RECT 1264.110 3508.560 1266.930 3509.040 ;
        RECT 1354.110 3508.560 1356.930 3509.040 ;
        RECT 1444.110 3508.560 1446.930 3509.040 ;
        RECT 1534.110 3508.560 1536.930 3509.040 ;
        RECT 1624.110 3508.560 1626.930 3509.040 ;
        RECT 1714.110 3508.560 1716.930 3509.040 ;
        RECT 1804.110 3508.560 1806.930 3509.040 ;
        RECT 1894.110 3508.560 1896.930 3509.040 ;
        RECT 1984.110 3508.560 1986.930 3509.040 ;
        RECT 2074.110 3508.560 2076.930 3509.040 ;
        RECT 2164.110 3508.560 2166.930 3509.040 ;
        RECT 2254.110 3508.560 2256.930 3509.040 ;
        RECT 2344.110 3508.560 2346.930 3509.040 ;
        RECT 2434.110 3508.560 2436.930 3509.040 ;
        RECT 2524.110 3508.560 2526.930 3509.040 ;
        RECT 2614.110 3508.560 2616.930 3509.040 ;
        RECT 2704.110 3508.560 2706.930 3509.040 ;
        RECT 2794.110 3508.560 2796.930 3509.040 ;
        RECT 2884.110 3508.560 2886.930 3509.040 ;
        RECT 94.110 10.640 96.930 11.120 ;
        RECT 184.110 10.640 186.930 11.120 ;
        RECT 274.110 10.640 276.930 11.120 ;
        RECT 364.110 10.640 366.930 11.120 ;
        RECT 454.110 10.640 456.930 11.120 ;
        RECT 544.110 10.640 546.930 11.120 ;
        RECT 634.110 10.640 636.930 11.120 ;
        RECT 724.110 10.640 726.930 11.120 ;
        RECT 814.110 10.640 816.930 11.120 ;
        RECT 904.110 10.640 906.930 11.120 ;
        RECT 994.110 10.640 996.930 11.120 ;
        RECT 1084.110 10.640 1086.930 11.120 ;
        RECT 1174.110 10.640 1176.930 11.120 ;
        RECT 1264.110 10.640 1266.930 11.120 ;
        RECT 1354.110 10.640 1356.930 11.120 ;
        RECT 1444.110 10.640 1446.930 11.120 ;
        RECT 1534.110 10.640 1536.930 11.120 ;
        RECT 1624.110 10.640 1626.930 11.120 ;
        RECT 1714.110 10.640 1716.930 11.120 ;
        RECT 1804.110 10.640 1806.930 11.120 ;
        RECT 1894.110 10.640 1896.930 11.120 ;
        RECT 1984.110 10.640 1986.930 11.120 ;
        RECT 2074.110 10.640 2076.930 11.120 ;
        RECT 2164.110 10.640 2166.930 11.120 ;
        RECT 2254.110 10.640 2256.930 11.120 ;
        RECT 2344.110 10.640 2346.930 11.120 ;
        RECT 2434.110 10.640 2436.930 11.120 ;
        RECT 2524.110 10.640 2526.930 11.120 ;
        RECT 2614.110 10.640 2616.930 11.120 ;
        RECT 2704.110 10.640 2706.930 11.120 ;
        RECT 2794.110 10.640 2796.930 11.120 ;
        RECT 2884.110 10.640 2886.930 11.120 ;
      LAYER via2 ;
        RECT 94.180 3508.660 94.460 3508.940 ;
        RECT 94.580 3508.660 94.860 3508.940 ;
        RECT 94.980 3508.660 95.260 3508.940 ;
        RECT 95.380 3508.660 95.660 3508.940 ;
        RECT 95.780 3508.660 96.060 3508.940 ;
        RECT 96.180 3508.660 96.460 3508.940 ;
        RECT 96.580 3508.660 96.860 3508.940 ;
        RECT 184.180 3508.660 184.460 3508.940 ;
        RECT 184.580 3508.660 184.860 3508.940 ;
        RECT 184.980 3508.660 185.260 3508.940 ;
        RECT 185.380 3508.660 185.660 3508.940 ;
        RECT 185.780 3508.660 186.060 3508.940 ;
        RECT 186.180 3508.660 186.460 3508.940 ;
        RECT 186.580 3508.660 186.860 3508.940 ;
        RECT 274.180 3508.660 274.460 3508.940 ;
        RECT 274.580 3508.660 274.860 3508.940 ;
        RECT 274.980 3508.660 275.260 3508.940 ;
        RECT 275.380 3508.660 275.660 3508.940 ;
        RECT 275.780 3508.660 276.060 3508.940 ;
        RECT 276.180 3508.660 276.460 3508.940 ;
        RECT 276.580 3508.660 276.860 3508.940 ;
        RECT 364.180 3508.660 364.460 3508.940 ;
        RECT 364.580 3508.660 364.860 3508.940 ;
        RECT 364.980 3508.660 365.260 3508.940 ;
        RECT 365.380 3508.660 365.660 3508.940 ;
        RECT 365.780 3508.660 366.060 3508.940 ;
        RECT 366.180 3508.660 366.460 3508.940 ;
        RECT 366.580 3508.660 366.860 3508.940 ;
        RECT 454.180 3508.660 454.460 3508.940 ;
        RECT 454.580 3508.660 454.860 3508.940 ;
        RECT 454.980 3508.660 455.260 3508.940 ;
        RECT 455.380 3508.660 455.660 3508.940 ;
        RECT 455.780 3508.660 456.060 3508.940 ;
        RECT 456.180 3508.660 456.460 3508.940 ;
        RECT 456.580 3508.660 456.860 3508.940 ;
        RECT 544.180 3508.660 544.460 3508.940 ;
        RECT 544.580 3508.660 544.860 3508.940 ;
        RECT 544.980 3508.660 545.260 3508.940 ;
        RECT 545.380 3508.660 545.660 3508.940 ;
        RECT 545.780 3508.660 546.060 3508.940 ;
        RECT 546.180 3508.660 546.460 3508.940 ;
        RECT 546.580 3508.660 546.860 3508.940 ;
        RECT 634.180 3508.660 634.460 3508.940 ;
        RECT 634.580 3508.660 634.860 3508.940 ;
        RECT 634.980 3508.660 635.260 3508.940 ;
        RECT 635.380 3508.660 635.660 3508.940 ;
        RECT 635.780 3508.660 636.060 3508.940 ;
        RECT 636.180 3508.660 636.460 3508.940 ;
        RECT 636.580 3508.660 636.860 3508.940 ;
        RECT 724.180 3508.660 724.460 3508.940 ;
        RECT 724.580 3508.660 724.860 3508.940 ;
        RECT 724.980 3508.660 725.260 3508.940 ;
        RECT 725.380 3508.660 725.660 3508.940 ;
        RECT 725.780 3508.660 726.060 3508.940 ;
        RECT 726.180 3508.660 726.460 3508.940 ;
        RECT 726.580 3508.660 726.860 3508.940 ;
        RECT 814.180 3508.660 814.460 3508.940 ;
        RECT 814.580 3508.660 814.860 3508.940 ;
        RECT 814.980 3508.660 815.260 3508.940 ;
        RECT 815.380 3508.660 815.660 3508.940 ;
        RECT 815.780 3508.660 816.060 3508.940 ;
        RECT 816.180 3508.660 816.460 3508.940 ;
        RECT 816.580 3508.660 816.860 3508.940 ;
        RECT 904.180 3508.660 904.460 3508.940 ;
        RECT 904.580 3508.660 904.860 3508.940 ;
        RECT 904.980 3508.660 905.260 3508.940 ;
        RECT 905.380 3508.660 905.660 3508.940 ;
        RECT 905.780 3508.660 906.060 3508.940 ;
        RECT 906.180 3508.660 906.460 3508.940 ;
        RECT 906.580 3508.660 906.860 3508.940 ;
        RECT 994.180 3508.660 994.460 3508.940 ;
        RECT 994.580 3508.660 994.860 3508.940 ;
        RECT 994.980 3508.660 995.260 3508.940 ;
        RECT 995.380 3508.660 995.660 3508.940 ;
        RECT 995.780 3508.660 996.060 3508.940 ;
        RECT 996.180 3508.660 996.460 3508.940 ;
        RECT 996.580 3508.660 996.860 3508.940 ;
        RECT 1084.180 3508.660 1084.460 3508.940 ;
        RECT 1084.580 3508.660 1084.860 3508.940 ;
        RECT 1084.980 3508.660 1085.260 3508.940 ;
        RECT 1085.380 3508.660 1085.660 3508.940 ;
        RECT 1085.780 3508.660 1086.060 3508.940 ;
        RECT 1086.180 3508.660 1086.460 3508.940 ;
        RECT 1086.580 3508.660 1086.860 3508.940 ;
        RECT 1174.180 3508.660 1174.460 3508.940 ;
        RECT 1174.580 3508.660 1174.860 3508.940 ;
        RECT 1174.980 3508.660 1175.260 3508.940 ;
        RECT 1175.380 3508.660 1175.660 3508.940 ;
        RECT 1175.780 3508.660 1176.060 3508.940 ;
        RECT 1176.180 3508.660 1176.460 3508.940 ;
        RECT 1176.580 3508.660 1176.860 3508.940 ;
        RECT 1264.180 3508.660 1264.460 3508.940 ;
        RECT 1264.580 3508.660 1264.860 3508.940 ;
        RECT 1264.980 3508.660 1265.260 3508.940 ;
        RECT 1265.380 3508.660 1265.660 3508.940 ;
        RECT 1265.780 3508.660 1266.060 3508.940 ;
        RECT 1266.180 3508.660 1266.460 3508.940 ;
        RECT 1266.580 3508.660 1266.860 3508.940 ;
        RECT 1354.180 3508.660 1354.460 3508.940 ;
        RECT 1354.580 3508.660 1354.860 3508.940 ;
        RECT 1354.980 3508.660 1355.260 3508.940 ;
        RECT 1355.380 3508.660 1355.660 3508.940 ;
        RECT 1355.780 3508.660 1356.060 3508.940 ;
        RECT 1356.180 3508.660 1356.460 3508.940 ;
        RECT 1356.580 3508.660 1356.860 3508.940 ;
        RECT 1444.180 3508.660 1444.460 3508.940 ;
        RECT 1444.580 3508.660 1444.860 3508.940 ;
        RECT 1444.980 3508.660 1445.260 3508.940 ;
        RECT 1445.380 3508.660 1445.660 3508.940 ;
        RECT 1445.780 3508.660 1446.060 3508.940 ;
        RECT 1446.180 3508.660 1446.460 3508.940 ;
        RECT 1446.580 3508.660 1446.860 3508.940 ;
        RECT 1534.180 3508.660 1534.460 3508.940 ;
        RECT 1534.580 3508.660 1534.860 3508.940 ;
        RECT 1534.980 3508.660 1535.260 3508.940 ;
        RECT 1535.380 3508.660 1535.660 3508.940 ;
        RECT 1535.780 3508.660 1536.060 3508.940 ;
        RECT 1536.180 3508.660 1536.460 3508.940 ;
        RECT 1536.580 3508.660 1536.860 3508.940 ;
        RECT 1624.180 3508.660 1624.460 3508.940 ;
        RECT 1624.580 3508.660 1624.860 3508.940 ;
        RECT 1624.980 3508.660 1625.260 3508.940 ;
        RECT 1625.380 3508.660 1625.660 3508.940 ;
        RECT 1625.780 3508.660 1626.060 3508.940 ;
        RECT 1626.180 3508.660 1626.460 3508.940 ;
        RECT 1626.580 3508.660 1626.860 3508.940 ;
        RECT 1714.180 3508.660 1714.460 3508.940 ;
        RECT 1714.580 3508.660 1714.860 3508.940 ;
        RECT 1714.980 3508.660 1715.260 3508.940 ;
        RECT 1715.380 3508.660 1715.660 3508.940 ;
        RECT 1715.780 3508.660 1716.060 3508.940 ;
        RECT 1716.180 3508.660 1716.460 3508.940 ;
        RECT 1716.580 3508.660 1716.860 3508.940 ;
        RECT 1804.180 3508.660 1804.460 3508.940 ;
        RECT 1804.580 3508.660 1804.860 3508.940 ;
        RECT 1804.980 3508.660 1805.260 3508.940 ;
        RECT 1805.380 3508.660 1805.660 3508.940 ;
        RECT 1805.780 3508.660 1806.060 3508.940 ;
        RECT 1806.180 3508.660 1806.460 3508.940 ;
        RECT 1806.580 3508.660 1806.860 3508.940 ;
        RECT 1894.180 3508.660 1894.460 3508.940 ;
        RECT 1894.580 3508.660 1894.860 3508.940 ;
        RECT 1894.980 3508.660 1895.260 3508.940 ;
        RECT 1895.380 3508.660 1895.660 3508.940 ;
        RECT 1895.780 3508.660 1896.060 3508.940 ;
        RECT 1896.180 3508.660 1896.460 3508.940 ;
        RECT 1896.580 3508.660 1896.860 3508.940 ;
        RECT 1984.180 3508.660 1984.460 3508.940 ;
        RECT 1984.580 3508.660 1984.860 3508.940 ;
        RECT 1984.980 3508.660 1985.260 3508.940 ;
        RECT 1985.380 3508.660 1985.660 3508.940 ;
        RECT 1985.780 3508.660 1986.060 3508.940 ;
        RECT 1986.180 3508.660 1986.460 3508.940 ;
        RECT 1986.580 3508.660 1986.860 3508.940 ;
        RECT 2074.180 3508.660 2074.460 3508.940 ;
        RECT 2074.580 3508.660 2074.860 3508.940 ;
        RECT 2074.980 3508.660 2075.260 3508.940 ;
        RECT 2075.380 3508.660 2075.660 3508.940 ;
        RECT 2075.780 3508.660 2076.060 3508.940 ;
        RECT 2076.180 3508.660 2076.460 3508.940 ;
        RECT 2076.580 3508.660 2076.860 3508.940 ;
        RECT 2164.180 3508.660 2164.460 3508.940 ;
        RECT 2164.580 3508.660 2164.860 3508.940 ;
        RECT 2164.980 3508.660 2165.260 3508.940 ;
        RECT 2165.380 3508.660 2165.660 3508.940 ;
        RECT 2165.780 3508.660 2166.060 3508.940 ;
        RECT 2166.180 3508.660 2166.460 3508.940 ;
        RECT 2166.580 3508.660 2166.860 3508.940 ;
        RECT 2254.180 3508.660 2254.460 3508.940 ;
        RECT 2254.580 3508.660 2254.860 3508.940 ;
        RECT 2254.980 3508.660 2255.260 3508.940 ;
        RECT 2255.380 3508.660 2255.660 3508.940 ;
        RECT 2255.780 3508.660 2256.060 3508.940 ;
        RECT 2256.180 3508.660 2256.460 3508.940 ;
        RECT 2256.580 3508.660 2256.860 3508.940 ;
        RECT 2344.180 3508.660 2344.460 3508.940 ;
        RECT 2344.580 3508.660 2344.860 3508.940 ;
        RECT 2344.980 3508.660 2345.260 3508.940 ;
        RECT 2345.380 3508.660 2345.660 3508.940 ;
        RECT 2345.780 3508.660 2346.060 3508.940 ;
        RECT 2346.180 3508.660 2346.460 3508.940 ;
        RECT 2346.580 3508.660 2346.860 3508.940 ;
        RECT 2434.180 3508.660 2434.460 3508.940 ;
        RECT 2434.580 3508.660 2434.860 3508.940 ;
        RECT 2434.980 3508.660 2435.260 3508.940 ;
        RECT 2435.380 3508.660 2435.660 3508.940 ;
        RECT 2435.780 3508.660 2436.060 3508.940 ;
        RECT 2436.180 3508.660 2436.460 3508.940 ;
        RECT 2436.580 3508.660 2436.860 3508.940 ;
        RECT 2524.180 3508.660 2524.460 3508.940 ;
        RECT 2524.580 3508.660 2524.860 3508.940 ;
        RECT 2524.980 3508.660 2525.260 3508.940 ;
        RECT 2525.380 3508.660 2525.660 3508.940 ;
        RECT 2525.780 3508.660 2526.060 3508.940 ;
        RECT 2526.180 3508.660 2526.460 3508.940 ;
        RECT 2526.580 3508.660 2526.860 3508.940 ;
        RECT 2614.180 3508.660 2614.460 3508.940 ;
        RECT 2614.580 3508.660 2614.860 3508.940 ;
        RECT 2614.980 3508.660 2615.260 3508.940 ;
        RECT 2615.380 3508.660 2615.660 3508.940 ;
        RECT 2615.780 3508.660 2616.060 3508.940 ;
        RECT 2616.180 3508.660 2616.460 3508.940 ;
        RECT 2616.580 3508.660 2616.860 3508.940 ;
        RECT 2704.180 3508.660 2704.460 3508.940 ;
        RECT 2704.580 3508.660 2704.860 3508.940 ;
        RECT 2704.980 3508.660 2705.260 3508.940 ;
        RECT 2705.380 3508.660 2705.660 3508.940 ;
        RECT 2705.780 3508.660 2706.060 3508.940 ;
        RECT 2706.180 3508.660 2706.460 3508.940 ;
        RECT 2706.580 3508.660 2706.860 3508.940 ;
        RECT 2794.180 3508.660 2794.460 3508.940 ;
        RECT 2794.580 3508.660 2794.860 3508.940 ;
        RECT 2794.980 3508.660 2795.260 3508.940 ;
        RECT 2795.380 3508.660 2795.660 3508.940 ;
        RECT 2795.780 3508.660 2796.060 3508.940 ;
        RECT 2796.180 3508.660 2796.460 3508.940 ;
        RECT 2796.580 3508.660 2796.860 3508.940 ;
        RECT 2884.180 3508.660 2884.460 3508.940 ;
        RECT 2884.580 3508.660 2884.860 3508.940 ;
        RECT 2884.980 3508.660 2885.260 3508.940 ;
        RECT 2885.380 3508.660 2885.660 3508.940 ;
        RECT 2885.780 3508.660 2886.060 3508.940 ;
        RECT 2886.180 3508.660 2886.460 3508.940 ;
        RECT 2886.580 3508.660 2886.860 3508.940 ;
        RECT 94.180 10.740 94.460 11.020 ;
        RECT 94.580 10.740 94.860 11.020 ;
        RECT 94.980 10.740 95.260 11.020 ;
        RECT 95.380 10.740 95.660 11.020 ;
        RECT 95.780 10.740 96.060 11.020 ;
        RECT 96.180 10.740 96.460 11.020 ;
        RECT 96.580 10.740 96.860 11.020 ;
        RECT 184.180 10.740 184.460 11.020 ;
        RECT 184.580 10.740 184.860 11.020 ;
        RECT 184.980 10.740 185.260 11.020 ;
        RECT 185.380 10.740 185.660 11.020 ;
        RECT 185.780 10.740 186.060 11.020 ;
        RECT 186.180 10.740 186.460 11.020 ;
        RECT 186.580 10.740 186.860 11.020 ;
        RECT 274.180 10.740 274.460 11.020 ;
        RECT 274.580 10.740 274.860 11.020 ;
        RECT 274.980 10.740 275.260 11.020 ;
        RECT 275.380 10.740 275.660 11.020 ;
        RECT 275.780 10.740 276.060 11.020 ;
        RECT 276.180 10.740 276.460 11.020 ;
        RECT 276.580 10.740 276.860 11.020 ;
        RECT 364.180 10.740 364.460 11.020 ;
        RECT 364.580 10.740 364.860 11.020 ;
        RECT 364.980 10.740 365.260 11.020 ;
        RECT 365.380 10.740 365.660 11.020 ;
        RECT 365.780 10.740 366.060 11.020 ;
        RECT 366.180 10.740 366.460 11.020 ;
        RECT 366.580 10.740 366.860 11.020 ;
        RECT 454.180 10.740 454.460 11.020 ;
        RECT 454.580 10.740 454.860 11.020 ;
        RECT 454.980 10.740 455.260 11.020 ;
        RECT 455.380 10.740 455.660 11.020 ;
        RECT 455.780 10.740 456.060 11.020 ;
        RECT 456.180 10.740 456.460 11.020 ;
        RECT 456.580 10.740 456.860 11.020 ;
        RECT 544.180 10.740 544.460 11.020 ;
        RECT 544.580 10.740 544.860 11.020 ;
        RECT 544.980 10.740 545.260 11.020 ;
        RECT 545.380 10.740 545.660 11.020 ;
        RECT 545.780 10.740 546.060 11.020 ;
        RECT 546.180 10.740 546.460 11.020 ;
        RECT 546.580 10.740 546.860 11.020 ;
        RECT 634.180 10.740 634.460 11.020 ;
        RECT 634.580 10.740 634.860 11.020 ;
        RECT 634.980 10.740 635.260 11.020 ;
        RECT 635.380 10.740 635.660 11.020 ;
        RECT 635.780 10.740 636.060 11.020 ;
        RECT 636.180 10.740 636.460 11.020 ;
        RECT 636.580 10.740 636.860 11.020 ;
        RECT 724.180 10.740 724.460 11.020 ;
        RECT 724.580 10.740 724.860 11.020 ;
        RECT 724.980 10.740 725.260 11.020 ;
        RECT 725.380 10.740 725.660 11.020 ;
        RECT 725.780 10.740 726.060 11.020 ;
        RECT 726.180 10.740 726.460 11.020 ;
        RECT 726.580 10.740 726.860 11.020 ;
        RECT 814.180 10.740 814.460 11.020 ;
        RECT 814.580 10.740 814.860 11.020 ;
        RECT 814.980 10.740 815.260 11.020 ;
        RECT 815.380 10.740 815.660 11.020 ;
        RECT 815.780 10.740 816.060 11.020 ;
        RECT 816.180 10.740 816.460 11.020 ;
        RECT 816.580 10.740 816.860 11.020 ;
        RECT 904.180 10.740 904.460 11.020 ;
        RECT 904.580 10.740 904.860 11.020 ;
        RECT 904.980 10.740 905.260 11.020 ;
        RECT 905.380 10.740 905.660 11.020 ;
        RECT 905.780 10.740 906.060 11.020 ;
        RECT 906.180 10.740 906.460 11.020 ;
        RECT 906.580 10.740 906.860 11.020 ;
        RECT 994.180 10.740 994.460 11.020 ;
        RECT 994.580 10.740 994.860 11.020 ;
        RECT 994.980 10.740 995.260 11.020 ;
        RECT 995.380 10.740 995.660 11.020 ;
        RECT 995.780 10.740 996.060 11.020 ;
        RECT 996.180 10.740 996.460 11.020 ;
        RECT 996.580 10.740 996.860 11.020 ;
        RECT 1084.180 10.740 1084.460 11.020 ;
        RECT 1084.580 10.740 1084.860 11.020 ;
        RECT 1084.980 10.740 1085.260 11.020 ;
        RECT 1085.380 10.740 1085.660 11.020 ;
        RECT 1085.780 10.740 1086.060 11.020 ;
        RECT 1086.180 10.740 1086.460 11.020 ;
        RECT 1086.580 10.740 1086.860 11.020 ;
        RECT 1174.180 10.740 1174.460 11.020 ;
        RECT 1174.580 10.740 1174.860 11.020 ;
        RECT 1174.980 10.740 1175.260 11.020 ;
        RECT 1175.380 10.740 1175.660 11.020 ;
        RECT 1175.780 10.740 1176.060 11.020 ;
        RECT 1176.180 10.740 1176.460 11.020 ;
        RECT 1176.580 10.740 1176.860 11.020 ;
        RECT 1264.180 10.740 1264.460 11.020 ;
        RECT 1264.580 10.740 1264.860 11.020 ;
        RECT 1264.980 10.740 1265.260 11.020 ;
        RECT 1265.380 10.740 1265.660 11.020 ;
        RECT 1265.780 10.740 1266.060 11.020 ;
        RECT 1266.180 10.740 1266.460 11.020 ;
        RECT 1266.580 10.740 1266.860 11.020 ;
        RECT 1354.180 10.740 1354.460 11.020 ;
        RECT 1354.580 10.740 1354.860 11.020 ;
        RECT 1354.980 10.740 1355.260 11.020 ;
        RECT 1355.380 10.740 1355.660 11.020 ;
        RECT 1355.780 10.740 1356.060 11.020 ;
        RECT 1356.180 10.740 1356.460 11.020 ;
        RECT 1356.580 10.740 1356.860 11.020 ;
        RECT 1444.180 10.740 1444.460 11.020 ;
        RECT 1444.580 10.740 1444.860 11.020 ;
        RECT 1444.980 10.740 1445.260 11.020 ;
        RECT 1445.380 10.740 1445.660 11.020 ;
        RECT 1445.780 10.740 1446.060 11.020 ;
        RECT 1446.180 10.740 1446.460 11.020 ;
        RECT 1446.580 10.740 1446.860 11.020 ;
        RECT 1534.180 10.740 1534.460 11.020 ;
        RECT 1534.580 10.740 1534.860 11.020 ;
        RECT 1534.980 10.740 1535.260 11.020 ;
        RECT 1535.380 10.740 1535.660 11.020 ;
        RECT 1535.780 10.740 1536.060 11.020 ;
        RECT 1536.180 10.740 1536.460 11.020 ;
        RECT 1536.580 10.740 1536.860 11.020 ;
        RECT 1624.180 10.740 1624.460 11.020 ;
        RECT 1624.580 10.740 1624.860 11.020 ;
        RECT 1624.980 10.740 1625.260 11.020 ;
        RECT 1625.380 10.740 1625.660 11.020 ;
        RECT 1625.780 10.740 1626.060 11.020 ;
        RECT 1626.180 10.740 1626.460 11.020 ;
        RECT 1626.580 10.740 1626.860 11.020 ;
        RECT 1714.180 10.740 1714.460 11.020 ;
        RECT 1714.580 10.740 1714.860 11.020 ;
        RECT 1714.980 10.740 1715.260 11.020 ;
        RECT 1715.380 10.740 1715.660 11.020 ;
        RECT 1715.780 10.740 1716.060 11.020 ;
        RECT 1716.180 10.740 1716.460 11.020 ;
        RECT 1716.580 10.740 1716.860 11.020 ;
        RECT 1804.180 10.740 1804.460 11.020 ;
        RECT 1804.580 10.740 1804.860 11.020 ;
        RECT 1804.980 10.740 1805.260 11.020 ;
        RECT 1805.380 10.740 1805.660 11.020 ;
        RECT 1805.780 10.740 1806.060 11.020 ;
        RECT 1806.180 10.740 1806.460 11.020 ;
        RECT 1806.580 10.740 1806.860 11.020 ;
        RECT 1894.180 10.740 1894.460 11.020 ;
        RECT 1894.580 10.740 1894.860 11.020 ;
        RECT 1894.980 10.740 1895.260 11.020 ;
        RECT 1895.380 10.740 1895.660 11.020 ;
        RECT 1895.780 10.740 1896.060 11.020 ;
        RECT 1896.180 10.740 1896.460 11.020 ;
        RECT 1896.580 10.740 1896.860 11.020 ;
        RECT 1984.180 10.740 1984.460 11.020 ;
        RECT 1984.580 10.740 1984.860 11.020 ;
        RECT 1984.980 10.740 1985.260 11.020 ;
        RECT 1985.380 10.740 1985.660 11.020 ;
        RECT 1985.780 10.740 1986.060 11.020 ;
        RECT 1986.180 10.740 1986.460 11.020 ;
        RECT 1986.580 10.740 1986.860 11.020 ;
        RECT 2074.180 10.740 2074.460 11.020 ;
        RECT 2074.580 10.740 2074.860 11.020 ;
        RECT 2074.980 10.740 2075.260 11.020 ;
        RECT 2075.380 10.740 2075.660 11.020 ;
        RECT 2075.780 10.740 2076.060 11.020 ;
        RECT 2076.180 10.740 2076.460 11.020 ;
        RECT 2076.580 10.740 2076.860 11.020 ;
        RECT 2164.180 10.740 2164.460 11.020 ;
        RECT 2164.580 10.740 2164.860 11.020 ;
        RECT 2164.980 10.740 2165.260 11.020 ;
        RECT 2165.380 10.740 2165.660 11.020 ;
        RECT 2165.780 10.740 2166.060 11.020 ;
        RECT 2166.180 10.740 2166.460 11.020 ;
        RECT 2166.580 10.740 2166.860 11.020 ;
        RECT 2254.180 10.740 2254.460 11.020 ;
        RECT 2254.580 10.740 2254.860 11.020 ;
        RECT 2254.980 10.740 2255.260 11.020 ;
        RECT 2255.380 10.740 2255.660 11.020 ;
        RECT 2255.780 10.740 2256.060 11.020 ;
        RECT 2256.180 10.740 2256.460 11.020 ;
        RECT 2256.580 10.740 2256.860 11.020 ;
        RECT 2344.180 10.740 2344.460 11.020 ;
        RECT 2344.580 10.740 2344.860 11.020 ;
        RECT 2344.980 10.740 2345.260 11.020 ;
        RECT 2345.380 10.740 2345.660 11.020 ;
        RECT 2345.780 10.740 2346.060 11.020 ;
        RECT 2346.180 10.740 2346.460 11.020 ;
        RECT 2346.580 10.740 2346.860 11.020 ;
        RECT 2434.180 10.740 2434.460 11.020 ;
        RECT 2434.580 10.740 2434.860 11.020 ;
        RECT 2434.980 10.740 2435.260 11.020 ;
        RECT 2435.380 10.740 2435.660 11.020 ;
        RECT 2435.780 10.740 2436.060 11.020 ;
        RECT 2436.180 10.740 2436.460 11.020 ;
        RECT 2436.580 10.740 2436.860 11.020 ;
        RECT 2524.180 10.740 2524.460 11.020 ;
        RECT 2524.580 10.740 2524.860 11.020 ;
        RECT 2524.980 10.740 2525.260 11.020 ;
        RECT 2525.380 10.740 2525.660 11.020 ;
        RECT 2525.780 10.740 2526.060 11.020 ;
        RECT 2526.180 10.740 2526.460 11.020 ;
        RECT 2526.580 10.740 2526.860 11.020 ;
        RECT 2614.180 10.740 2614.460 11.020 ;
        RECT 2614.580 10.740 2614.860 11.020 ;
        RECT 2614.980 10.740 2615.260 11.020 ;
        RECT 2615.380 10.740 2615.660 11.020 ;
        RECT 2615.780 10.740 2616.060 11.020 ;
        RECT 2616.180 10.740 2616.460 11.020 ;
        RECT 2616.580 10.740 2616.860 11.020 ;
        RECT 2704.180 10.740 2704.460 11.020 ;
        RECT 2704.580 10.740 2704.860 11.020 ;
        RECT 2704.980 10.740 2705.260 11.020 ;
        RECT 2705.380 10.740 2705.660 11.020 ;
        RECT 2705.780 10.740 2706.060 11.020 ;
        RECT 2706.180 10.740 2706.460 11.020 ;
        RECT 2706.580 10.740 2706.860 11.020 ;
        RECT 2794.180 10.740 2794.460 11.020 ;
        RECT 2794.580 10.740 2794.860 11.020 ;
        RECT 2794.980 10.740 2795.260 11.020 ;
        RECT 2795.380 10.740 2795.660 11.020 ;
        RECT 2795.780 10.740 2796.060 11.020 ;
        RECT 2796.180 10.740 2796.460 11.020 ;
        RECT 2796.580 10.740 2796.860 11.020 ;
        RECT 2884.180 10.740 2884.460 11.020 ;
        RECT 2884.580 10.740 2884.860 11.020 ;
        RECT 2884.980 10.740 2885.260 11.020 ;
        RECT 2885.380 10.740 2885.660 11.020 ;
        RECT 2885.780 10.740 2886.060 11.020 ;
        RECT 2886.180 10.740 2886.460 11.020 ;
        RECT 2886.580 10.740 2886.860 11.020 ;
      LAYER met3 ;
        RECT 94.020 3508.635 97.020 3508.965 ;
        RECT 184.020 3508.635 187.020 3508.965 ;
        RECT 274.020 3508.635 277.020 3508.965 ;
        RECT 364.020 3508.635 367.020 3508.965 ;
        RECT 454.020 3508.635 457.020 3508.965 ;
        RECT 544.020 3508.635 547.020 3508.965 ;
        RECT 634.020 3508.635 637.020 3508.965 ;
        RECT 724.020 3508.635 727.020 3508.965 ;
        RECT 814.020 3508.635 817.020 3508.965 ;
        RECT 904.020 3508.635 907.020 3508.965 ;
        RECT 994.020 3508.635 997.020 3508.965 ;
        RECT 1084.020 3508.635 1087.020 3508.965 ;
        RECT 1174.020 3508.635 1177.020 3508.965 ;
        RECT 1264.020 3508.635 1267.020 3508.965 ;
        RECT 1354.020 3508.635 1357.020 3508.965 ;
        RECT 1444.020 3508.635 1447.020 3508.965 ;
        RECT 1534.020 3508.635 1537.020 3508.965 ;
        RECT 1624.020 3508.635 1627.020 3508.965 ;
        RECT 1714.020 3508.635 1717.020 3508.965 ;
        RECT 1804.020 3508.635 1807.020 3508.965 ;
        RECT 1894.020 3508.635 1897.020 3508.965 ;
        RECT 1984.020 3508.635 1987.020 3508.965 ;
        RECT 2074.020 3508.635 2077.020 3508.965 ;
        RECT 2164.020 3508.635 2167.020 3508.965 ;
        RECT 2254.020 3508.635 2257.020 3508.965 ;
        RECT 2344.020 3508.635 2347.020 3508.965 ;
        RECT 2434.020 3508.635 2437.020 3508.965 ;
        RECT 2524.020 3508.635 2527.020 3508.965 ;
        RECT 2614.020 3508.635 2617.020 3508.965 ;
        RECT 2704.020 3508.635 2707.020 3508.965 ;
        RECT 2794.020 3508.635 2797.020 3508.965 ;
        RECT 2884.020 3508.635 2887.020 3508.965 ;
        RECT 94.020 10.715 97.020 11.045 ;
        RECT 184.020 10.715 187.020 11.045 ;
        RECT 274.020 10.715 277.020 11.045 ;
        RECT 364.020 10.715 367.020 11.045 ;
        RECT 454.020 10.715 457.020 11.045 ;
        RECT 544.020 10.715 547.020 11.045 ;
        RECT 634.020 10.715 637.020 11.045 ;
        RECT 724.020 10.715 727.020 11.045 ;
        RECT 814.020 10.715 817.020 11.045 ;
        RECT 904.020 10.715 907.020 11.045 ;
        RECT 994.020 10.715 997.020 11.045 ;
        RECT 1084.020 10.715 1087.020 11.045 ;
        RECT 1174.020 10.715 1177.020 11.045 ;
        RECT 1264.020 10.715 1267.020 11.045 ;
        RECT 1354.020 10.715 1357.020 11.045 ;
        RECT 1444.020 10.715 1447.020 11.045 ;
        RECT 1534.020 10.715 1537.020 11.045 ;
        RECT 1624.020 10.715 1627.020 11.045 ;
        RECT 1714.020 10.715 1717.020 11.045 ;
        RECT 1804.020 10.715 1807.020 11.045 ;
        RECT 1894.020 10.715 1897.020 11.045 ;
        RECT 1984.020 10.715 1987.020 11.045 ;
        RECT 2074.020 10.715 2077.020 11.045 ;
        RECT 2164.020 10.715 2167.020 11.045 ;
        RECT 2254.020 10.715 2257.020 11.045 ;
        RECT 2344.020 10.715 2347.020 11.045 ;
        RECT 2434.020 10.715 2437.020 11.045 ;
        RECT 2524.020 10.715 2527.020 11.045 ;
        RECT 2614.020 10.715 2617.020 11.045 ;
        RECT 2704.020 10.715 2707.020 11.045 ;
        RECT 2794.020 10.715 2797.020 11.045 ;
        RECT 2884.020 10.715 2887.020 11.045 ;
      LAYER via3 ;
        RECT 94.160 3508.640 94.480 3508.960 ;
        RECT 94.560 3508.640 94.880 3508.960 ;
        RECT 94.960 3508.640 95.280 3508.960 ;
        RECT 95.360 3508.640 95.680 3508.960 ;
        RECT 95.760 3508.640 96.080 3508.960 ;
        RECT 96.160 3508.640 96.480 3508.960 ;
        RECT 96.560 3508.640 96.880 3508.960 ;
        RECT 184.160 3508.640 184.480 3508.960 ;
        RECT 184.560 3508.640 184.880 3508.960 ;
        RECT 184.960 3508.640 185.280 3508.960 ;
        RECT 185.360 3508.640 185.680 3508.960 ;
        RECT 185.760 3508.640 186.080 3508.960 ;
        RECT 186.160 3508.640 186.480 3508.960 ;
        RECT 186.560 3508.640 186.880 3508.960 ;
        RECT 274.160 3508.640 274.480 3508.960 ;
        RECT 274.560 3508.640 274.880 3508.960 ;
        RECT 274.960 3508.640 275.280 3508.960 ;
        RECT 275.360 3508.640 275.680 3508.960 ;
        RECT 275.760 3508.640 276.080 3508.960 ;
        RECT 276.160 3508.640 276.480 3508.960 ;
        RECT 276.560 3508.640 276.880 3508.960 ;
        RECT 364.160 3508.640 364.480 3508.960 ;
        RECT 364.560 3508.640 364.880 3508.960 ;
        RECT 364.960 3508.640 365.280 3508.960 ;
        RECT 365.360 3508.640 365.680 3508.960 ;
        RECT 365.760 3508.640 366.080 3508.960 ;
        RECT 366.160 3508.640 366.480 3508.960 ;
        RECT 366.560 3508.640 366.880 3508.960 ;
        RECT 454.160 3508.640 454.480 3508.960 ;
        RECT 454.560 3508.640 454.880 3508.960 ;
        RECT 454.960 3508.640 455.280 3508.960 ;
        RECT 455.360 3508.640 455.680 3508.960 ;
        RECT 455.760 3508.640 456.080 3508.960 ;
        RECT 456.160 3508.640 456.480 3508.960 ;
        RECT 456.560 3508.640 456.880 3508.960 ;
        RECT 544.160 3508.640 544.480 3508.960 ;
        RECT 544.560 3508.640 544.880 3508.960 ;
        RECT 544.960 3508.640 545.280 3508.960 ;
        RECT 545.360 3508.640 545.680 3508.960 ;
        RECT 545.760 3508.640 546.080 3508.960 ;
        RECT 546.160 3508.640 546.480 3508.960 ;
        RECT 546.560 3508.640 546.880 3508.960 ;
        RECT 634.160 3508.640 634.480 3508.960 ;
        RECT 634.560 3508.640 634.880 3508.960 ;
        RECT 634.960 3508.640 635.280 3508.960 ;
        RECT 635.360 3508.640 635.680 3508.960 ;
        RECT 635.760 3508.640 636.080 3508.960 ;
        RECT 636.160 3508.640 636.480 3508.960 ;
        RECT 636.560 3508.640 636.880 3508.960 ;
        RECT 724.160 3508.640 724.480 3508.960 ;
        RECT 724.560 3508.640 724.880 3508.960 ;
        RECT 724.960 3508.640 725.280 3508.960 ;
        RECT 725.360 3508.640 725.680 3508.960 ;
        RECT 725.760 3508.640 726.080 3508.960 ;
        RECT 726.160 3508.640 726.480 3508.960 ;
        RECT 726.560 3508.640 726.880 3508.960 ;
        RECT 814.160 3508.640 814.480 3508.960 ;
        RECT 814.560 3508.640 814.880 3508.960 ;
        RECT 814.960 3508.640 815.280 3508.960 ;
        RECT 815.360 3508.640 815.680 3508.960 ;
        RECT 815.760 3508.640 816.080 3508.960 ;
        RECT 816.160 3508.640 816.480 3508.960 ;
        RECT 816.560 3508.640 816.880 3508.960 ;
        RECT 904.160 3508.640 904.480 3508.960 ;
        RECT 904.560 3508.640 904.880 3508.960 ;
        RECT 904.960 3508.640 905.280 3508.960 ;
        RECT 905.360 3508.640 905.680 3508.960 ;
        RECT 905.760 3508.640 906.080 3508.960 ;
        RECT 906.160 3508.640 906.480 3508.960 ;
        RECT 906.560 3508.640 906.880 3508.960 ;
        RECT 994.160 3508.640 994.480 3508.960 ;
        RECT 994.560 3508.640 994.880 3508.960 ;
        RECT 994.960 3508.640 995.280 3508.960 ;
        RECT 995.360 3508.640 995.680 3508.960 ;
        RECT 995.760 3508.640 996.080 3508.960 ;
        RECT 996.160 3508.640 996.480 3508.960 ;
        RECT 996.560 3508.640 996.880 3508.960 ;
        RECT 1084.160 3508.640 1084.480 3508.960 ;
        RECT 1084.560 3508.640 1084.880 3508.960 ;
        RECT 1084.960 3508.640 1085.280 3508.960 ;
        RECT 1085.360 3508.640 1085.680 3508.960 ;
        RECT 1085.760 3508.640 1086.080 3508.960 ;
        RECT 1086.160 3508.640 1086.480 3508.960 ;
        RECT 1086.560 3508.640 1086.880 3508.960 ;
        RECT 1174.160 3508.640 1174.480 3508.960 ;
        RECT 1174.560 3508.640 1174.880 3508.960 ;
        RECT 1174.960 3508.640 1175.280 3508.960 ;
        RECT 1175.360 3508.640 1175.680 3508.960 ;
        RECT 1175.760 3508.640 1176.080 3508.960 ;
        RECT 1176.160 3508.640 1176.480 3508.960 ;
        RECT 1176.560 3508.640 1176.880 3508.960 ;
        RECT 1264.160 3508.640 1264.480 3508.960 ;
        RECT 1264.560 3508.640 1264.880 3508.960 ;
        RECT 1264.960 3508.640 1265.280 3508.960 ;
        RECT 1265.360 3508.640 1265.680 3508.960 ;
        RECT 1265.760 3508.640 1266.080 3508.960 ;
        RECT 1266.160 3508.640 1266.480 3508.960 ;
        RECT 1266.560 3508.640 1266.880 3508.960 ;
        RECT 1354.160 3508.640 1354.480 3508.960 ;
        RECT 1354.560 3508.640 1354.880 3508.960 ;
        RECT 1354.960 3508.640 1355.280 3508.960 ;
        RECT 1355.360 3508.640 1355.680 3508.960 ;
        RECT 1355.760 3508.640 1356.080 3508.960 ;
        RECT 1356.160 3508.640 1356.480 3508.960 ;
        RECT 1356.560 3508.640 1356.880 3508.960 ;
        RECT 1444.160 3508.640 1444.480 3508.960 ;
        RECT 1444.560 3508.640 1444.880 3508.960 ;
        RECT 1444.960 3508.640 1445.280 3508.960 ;
        RECT 1445.360 3508.640 1445.680 3508.960 ;
        RECT 1445.760 3508.640 1446.080 3508.960 ;
        RECT 1446.160 3508.640 1446.480 3508.960 ;
        RECT 1446.560 3508.640 1446.880 3508.960 ;
        RECT 1534.160 3508.640 1534.480 3508.960 ;
        RECT 1534.560 3508.640 1534.880 3508.960 ;
        RECT 1534.960 3508.640 1535.280 3508.960 ;
        RECT 1535.360 3508.640 1535.680 3508.960 ;
        RECT 1535.760 3508.640 1536.080 3508.960 ;
        RECT 1536.160 3508.640 1536.480 3508.960 ;
        RECT 1536.560 3508.640 1536.880 3508.960 ;
        RECT 1624.160 3508.640 1624.480 3508.960 ;
        RECT 1624.560 3508.640 1624.880 3508.960 ;
        RECT 1624.960 3508.640 1625.280 3508.960 ;
        RECT 1625.360 3508.640 1625.680 3508.960 ;
        RECT 1625.760 3508.640 1626.080 3508.960 ;
        RECT 1626.160 3508.640 1626.480 3508.960 ;
        RECT 1626.560 3508.640 1626.880 3508.960 ;
        RECT 1714.160 3508.640 1714.480 3508.960 ;
        RECT 1714.560 3508.640 1714.880 3508.960 ;
        RECT 1714.960 3508.640 1715.280 3508.960 ;
        RECT 1715.360 3508.640 1715.680 3508.960 ;
        RECT 1715.760 3508.640 1716.080 3508.960 ;
        RECT 1716.160 3508.640 1716.480 3508.960 ;
        RECT 1716.560 3508.640 1716.880 3508.960 ;
        RECT 1804.160 3508.640 1804.480 3508.960 ;
        RECT 1804.560 3508.640 1804.880 3508.960 ;
        RECT 1804.960 3508.640 1805.280 3508.960 ;
        RECT 1805.360 3508.640 1805.680 3508.960 ;
        RECT 1805.760 3508.640 1806.080 3508.960 ;
        RECT 1806.160 3508.640 1806.480 3508.960 ;
        RECT 1806.560 3508.640 1806.880 3508.960 ;
        RECT 1894.160 3508.640 1894.480 3508.960 ;
        RECT 1894.560 3508.640 1894.880 3508.960 ;
        RECT 1894.960 3508.640 1895.280 3508.960 ;
        RECT 1895.360 3508.640 1895.680 3508.960 ;
        RECT 1895.760 3508.640 1896.080 3508.960 ;
        RECT 1896.160 3508.640 1896.480 3508.960 ;
        RECT 1896.560 3508.640 1896.880 3508.960 ;
        RECT 1984.160 3508.640 1984.480 3508.960 ;
        RECT 1984.560 3508.640 1984.880 3508.960 ;
        RECT 1984.960 3508.640 1985.280 3508.960 ;
        RECT 1985.360 3508.640 1985.680 3508.960 ;
        RECT 1985.760 3508.640 1986.080 3508.960 ;
        RECT 1986.160 3508.640 1986.480 3508.960 ;
        RECT 1986.560 3508.640 1986.880 3508.960 ;
        RECT 2074.160 3508.640 2074.480 3508.960 ;
        RECT 2074.560 3508.640 2074.880 3508.960 ;
        RECT 2074.960 3508.640 2075.280 3508.960 ;
        RECT 2075.360 3508.640 2075.680 3508.960 ;
        RECT 2075.760 3508.640 2076.080 3508.960 ;
        RECT 2076.160 3508.640 2076.480 3508.960 ;
        RECT 2076.560 3508.640 2076.880 3508.960 ;
        RECT 2164.160 3508.640 2164.480 3508.960 ;
        RECT 2164.560 3508.640 2164.880 3508.960 ;
        RECT 2164.960 3508.640 2165.280 3508.960 ;
        RECT 2165.360 3508.640 2165.680 3508.960 ;
        RECT 2165.760 3508.640 2166.080 3508.960 ;
        RECT 2166.160 3508.640 2166.480 3508.960 ;
        RECT 2166.560 3508.640 2166.880 3508.960 ;
        RECT 2254.160 3508.640 2254.480 3508.960 ;
        RECT 2254.560 3508.640 2254.880 3508.960 ;
        RECT 2254.960 3508.640 2255.280 3508.960 ;
        RECT 2255.360 3508.640 2255.680 3508.960 ;
        RECT 2255.760 3508.640 2256.080 3508.960 ;
        RECT 2256.160 3508.640 2256.480 3508.960 ;
        RECT 2256.560 3508.640 2256.880 3508.960 ;
        RECT 2344.160 3508.640 2344.480 3508.960 ;
        RECT 2344.560 3508.640 2344.880 3508.960 ;
        RECT 2344.960 3508.640 2345.280 3508.960 ;
        RECT 2345.360 3508.640 2345.680 3508.960 ;
        RECT 2345.760 3508.640 2346.080 3508.960 ;
        RECT 2346.160 3508.640 2346.480 3508.960 ;
        RECT 2346.560 3508.640 2346.880 3508.960 ;
        RECT 2434.160 3508.640 2434.480 3508.960 ;
        RECT 2434.560 3508.640 2434.880 3508.960 ;
        RECT 2434.960 3508.640 2435.280 3508.960 ;
        RECT 2435.360 3508.640 2435.680 3508.960 ;
        RECT 2435.760 3508.640 2436.080 3508.960 ;
        RECT 2436.160 3508.640 2436.480 3508.960 ;
        RECT 2436.560 3508.640 2436.880 3508.960 ;
        RECT 2524.160 3508.640 2524.480 3508.960 ;
        RECT 2524.560 3508.640 2524.880 3508.960 ;
        RECT 2524.960 3508.640 2525.280 3508.960 ;
        RECT 2525.360 3508.640 2525.680 3508.960 ;
        RECT 2525.760 3508.640 2526.080 3508.960 ;
        RECT 2526.160 3508.640 2526.480 3508.960 ;
        RECT 2526.560 3508.640 2526.880 3508.960 ;
        RECT 2614.160 3508.640 2614.480 3508.960 ;
        RECT 2614.560 3508.640 2614.880 3508.960 ;
        RECT 2614.960 3508.640 2615.280 3508.960 ;
        RECT 2615.360 3508.640 2615.680 3508.960 ;
        RECT 2615.760 3508.640 2616.080 3508.960 ;
        RECT 2616.160 3508.640 2616.480 3508.960 ;
        RECT 2616.560 3508.640 2616.880 3508.960 ;
        RECT 2704.160 3508.640 2704.480 3508.960 ;
        RECT 2704.560 3508.640 2704.880 3508.960 ;
        RECT 2704.960 3508.640 2705.280 3508.960 ;
        RECT 2705.360 3508.640 2705.680 3508.960 ;
        RECT 2705.760 3508.640 2706.080 3508.960 ;
        RECT 2706.160 3508.640 2706.480 3508.960 ;
        RECT 2706.560 3508.640 2706.880 3508.960 ;
        RECT 2794.160 3508.640 2794.480 3508.960 ;
        RECT 2794.560 3508.640 2794.880 3508.960 ;
        RECT 2794.960 3508.640 2795.280 3508.960 ;
        RECT 2795.360 3508.640 2795.680 3508.960 ;
        RECT 2795.760 3508.640 2796.080 3508.960 ;
        RECT 2796.160 3508.640 2796.480 3508.960 ;
        RECT 2796.560 3508.640 2796.880 3508.960 ;
        RECT 2884.160 3508.640 2884.480 3508.960 ;
        RECT 2884.560 3508.640 2884.880 3508.960 ;
        RECT 2884.960 3508.640 2885.280 3508.960 ;
        RECT 2885.360 3508.640 2885.680 3508.960 ;
        RECT 2885.760 3508.640 2886.080 3508.960 ;
        RECT 2886.160 3508.640 2886.480 3508.960 ;
        RECT 2886.560 3508.640 2886.880 3508.960 ;
        RECT 94.160 10.720 94.480 11.040 ;
        RECT 94.560 10.720 94.880 11.040 ;
        RECT 94.960 10.720 95.280 11.040 ;
        RECT 95.360 10.720 95.680 11.040 ;
        RECT 95.760 10.720 96.080 11.040 ;
        RECT 96.160 10.720 96.480 11.040 ;
        RECT 96.560 10.720 96.880 11.040 ;
        RECT 184.160 10.720 184.480 11.040 ;
        RECT 184.560 10.720 184.880 11.040 ;
        RECT 184.960 10.720 185.280 11.040 ;
        RECT 185.360 10.720 185.680 11.040 ;
        RECT 185.760 10.720 186.080 11.040 ;
        RECT 186.160 10.720 186.480 11.040 ;
        RECT 186.560 10.720 186.880 11.040 ;
        RECT 274.160 10.720 274.480 11.040 ;
        RECT 274.560 10.720 274.880 11.040 ;
        RECT 274.960 10.720 275.280 11.040 ;
        RECT 275.360 10.720 275.680 11.040 ;
        RECT 275.760 10.720 276.080 11.040 ;
        RECT 276.160 10.720 276.480 11.040 ;
        RECT 276.560 10.720 276.880 11.040 ;
        RECT 364.160 10.720 364.480 11.040 ;
        RECT 364.560 10.720 364.880 11.040 ;
        RECT 364.960 10.720 365.280 11.040 ;
        RECT 365.360 10.720 365.680 11.040 ;
        RECT 365.760 10.720 366.080 11.040 ;
        RECT 366.160 10.720 366.480 11.040 ;
        RECT 366.560 10.720 366.880 11.040 ;
        RECT 454.160 10.720 454.480 11.040 ;
        RECT 454.560 10.720 454.880 11.040 ;
        RECT 454.960 10.720 455.280 11.040 ;
        RECT 455.360 10.720 455.680 11.040 ;
        RECT 455.760 10.720 456.080 11.040 ;
        RECT 456.160 10.720 456.480 11.040 ;
        RECT 456.560 10.720 456.880 11.040 ;
        RECT 544.160 10.720 544.480 11.040 ;
        RECT 544.560 10.720 544.880 11.040 ;
        RECT 544.960 10.720 545.280 11.040 ;
        RECT 545.360 10.720 545.680 11.040 ;
        RECT 545.760 10.720 546.080 11.040 ;
        RECT 546.160 10.720 546.480 11.040 ;
        RECT 546.560 10.720 546.880 11.040 ;
        RECT 634.160 10.720 634.480 11.040 ;
        RECT 634.560 10.720 634.880 11.040 ;
        RECT 634.960 10.720 635.280 11.040 ;
        RECT 635.360 10.720 635.680 11.040 ;
        RECT 635.760 10.720 636.080 11.040 ;
        RECT 636.160 10.720 636.480 11.040 ;
        RECT 636.560 10.720 636.880 11.040 ;
        RECT 724.160 10.720 724.480 11.040 ;
        RECT 724.560 10.720 724.880 11.040 ;
        RECT 724.960 10.720 725.280 11.040 ;
        RECT 725.360 10.720 725.680 11.040 ;
        RECT 725.760 10.720 726.080 11.040 ;
        RECT 726.160 10.720 726.480 11.040 ;
        RECT 726.560 10.720 726.880 11.040 ;
        RECT 814.160 10.720 814.480 11.040 ;
        RECT 814.560 10.720 814.880 11.040 ;
        RECT 814.960 10.720 815.280 11.040 ;
        RECT 815.360 10.720 815.680 11.040 ;
        RECT 815.760 10.720 816.080 11.040 ;
        RECT 816.160 10.720 816.480 11.040 ;
        RECT 816.560 10.720 816.880 11.040 ;
        RECT 904.160 10.720 904.480 11.040 ;
        RECT 904.560 10.720 904.880 11.040 ;
        RECT 904.960 10.720 905.280 11.040 ;
        RECT 905.360 10.720 905.680 11.040 ;
        RECT 905.760 10.720 906.080 11.040 ;
        RECT 906.160 10.720 906.480 11.040 ;
        RECT 906.560 10.720 906.880 11.040 ;
        RECT 994.160 10.720 994.480 11.040 ;
        RECT 994.560 10.720 994.880 11.040 ;
        RECT 994.960 10.720 995.280 11.040 ;
        RECT 995.360 10.720 995.680 11.040 ;
        RECT 995.760 10.720 996.080 11.040 ;
        RECT 996.160 10.720 996.480 11.040 ;
        RECT 996.560 10.720 996.880 11.040 ;
        RECT 1084.160 10.720 1084.480 11.040 ;
        RECT 1084.560 10.720 1084.880 11.040 ;
        RECT 1084.960 10.720 1085.280 11.040 ;
        RECT 1085.360 10.720 1085.680 11.040 ;
        RECT 1085.760 10.720 1086.080 11.040 ;
        RECT 1086.160 10.720 1086.480 11.040 ;
        RECT 1086.560 10.720 1086.880 11.040 ;
        RECT 1174.160 10.720 1174.480 11.040 ;
        RECT 1174.560 10.720 1174.880 11.040 ;
        RECT 1174.960 10.720 1175.280 11.040 ;
        RECT 1175.360 10.720 1175.680 11.040 ;
        RECT 1175.760 10.720 1176.080 11.040 ;
        RECT 1176.160 10.720 1176.480 11.040 ;
        RECT 1176.560 10.720 1176.880 11.040 ;
        RECT 1264.160 10.720 1264.480 11.040 ;
        RECT 1264.560 10.720 1264.880 11.040 ;
        RECT 1264.960 10.720 1265.280 11.040 ;
        RECT 1265.360 10.720 1265.680 11.040 ;
        RECT 1265.760 10.720 1266.080 11.040 ;
        RECT 1266.160 10.720 1266.480 11.040 ;
        RECT 1266.560 10.720 1266.880 11.040 ;
        RECT 1354.160 10.720 1354.480 11.040 ;
        RECT 1354.560 10.720 1354.880 11.040 ;
        RECT 1354.960 10.720 1355.280 11.040 ;
        RECT 1355.360 10.720 1355.680 11.040 ;
        RECT 1355.760 10.720 1356.080 11.040 ;
        RECT 1356.160 10.720 1356.480 11.040 ;
        RECT 1356.560 10.720 1356.880 11.040 ;
        RECT 1444.160 10.720 1444.480 11.040 ;
        RECT 1444.560 10.720 1444.880 11.040 ;
        RECT 1444.960 10.720 1445.280 11.040 ;
        RECT 1445.360 10.720 1445.680 11.040 ;
        RECT 1445.760 10.720 1446.080 11.040 ;
        RECT 1446.160 10.720 1446.480 11.040 ;
        RECT 1446.560 10.720 1446.880 11.040 ;
        RECT 1534.160 10.720 1534.480 11.040 ;
        RECT 1534.560 10.720 1534.880 11.040 ;
        RECT 1534.960 10.720 1535.280 11.040 ;
        RECT 1535.360 10.720 1535.680 11.040 ;
        RECT 1535.760 10.720 1536.080 11.040 ;
        RECT 1536.160 10.720 1536.480 11.040 ;
        RECT 1536.560 10.720 1536.880 11.040 ;
        RECT 1624.160 10.720 1624.480 11.040 ;
        RECT 1624.560 10.720 1624.880 11.040 ;
        RECT 1624.960 10.720 1625.280 11.040 ;
        RECT 1625.360 10.720 1625.680 11.040 ;
        RECT 1625.760 10.720 1626.080 11.040 ;
        RECT 1626.160 10.720 1626.480 11.040 ;
        RECT 1626.560 10.720 1626.880 11.040 ;
        RECT 1714.160 10.720 1714.480 11.040 ;
        RECT 1714.560 10.720 1714.880 11.040 ;
        RECT 1714.960 10.720 1715.280 11.040 ;
        RECT 1715.360 10.720 1715.680 11.040 ;
        RECT 1715.760 10.720 1716.080 11.040 ;
        RECT 1716.160 10.720 1716.480 11.040 ;
        RECT 1716.560 10.720 1716.880 11.040 ;
        RECT 1804.160 10.720 1804.480 11.040 ;
        RECT 1804.560 10.720 1804.880 11.040 ;
        RECT 1804.960 10.720 1805.280 11.040 ;
        RECT 1805.360 10.720 1805.680 11.040 ;
        RECT 1805.760 10.720 1806.080 11.040 ;
        RECT 1806.160 10.720 1806.480 11.040 ;
        RECT 1806.560 10.720 1806.880 11.040 ;
        RECT 1894.160 10.720 1894.480 11.040 ;
        RECT 1894.560 10.720 1894.880 11.040 ;
        RECT 1894.960 10.720 1895.280 11.040 ;
        RECT 1895.360 10.720 1895.680 11.040 ;
        RECT 1895.760 10.720 1896.080 11.040 ;
        RECT 1896.160 10.720 1896.480 11.040 ;
        RECT 1896.560 10.720 1896.880 11.040 ;
        RECT 1984.160 10.720 1984.480 11.040 ;
        RECT 1984.560 10.720 1984.880 11.040 ;
        RECT 1984.960 10.720 1985.280 11.040 ;
        RECT 1985.360 10.720 1985.680 11.040 ;
        RECT 1985.760 10.720 1986.080 11.040 ;
        RECT 1986.160 10.720 1986.480 11.040 ;
        RECT 1986.560 10.720 1986.880 11.040 ;
        RECT 2074.160 10.720 2074.480 11.040 ;
        RECT 2074.560 10.720 2074.880 11.040 ;
        RECT 2074.960 10.720 2075.280 11.040 ;
        RECT 2075.360 10.720 2075.680 11.040 ;
        RECT 2075.760 10.720 2076.080 11.040 ;
        RECT 2076.160 10.720 2076.480 11.040 ;
        RECT 2076.560 10.720 2076.880 11.040 ;
        RECT 2164.160 10.720 2164.480 11.040 ;
        RECT 2164.560 10.720 2164.880 11.040 ;
        RECT 2164.960 10.720 2165.280 11.040 ;
        RECT 2165.360 10.720 2165.680 11.040 ;
        RECT 2165.760 10.720 2166.080 11.040 ;
        RECT 2166.160 10.720 2166.480 11.040 ;
        RECT 2166.560 10.720 2166.880 11.040 ;
        RECT 2254.160 10.720 2254.480 11.040 ;
        RECT 2254.560 10.720 2254.880 11.040 ;
        RECT 2254.960 10.720 2255.280 11.040 ;
        RECT 2255.360 10.720 2255.680 11.040 ;
        RECT 2255.760 10.720 2256.080 11.040 ;
        RECT 2256.160 10.720 2256.480 11.040 ;
        RECT 2256.560 10.720 2256.880 11.040 ;
        RECT 2344.160 10.720 2344.480 11.040 ;
        RECT 2344.560 10.720 2344.880 11.040 ;
        RECT 2344.960 10.720 2345.280 11.040 ;
        RECT 2345.360 10.720 2345.680 11.040 ;
        RECT 2345.760 10.720 2346.080 11.040 ;
        RECT 2346.160 10.720 2346.480 11.040 ;
        RECT 2346.560 10.720 2346.880 11.040 ;
        RECT 2434.160 10.720 2434.480 11.040 ;
        RECT 2434.560 10.720 2434.880 11.040 ;
        RECT 2434.960 10.720 2435.280 11.040 ;
        RECT 2435.360 10.720 2435.680 11.040 ;
        RECT 2435.760 10.720 2436.080 11.040 ;
        RECT 2436.160 10.720 2436.480 11.040 ;
        RECT 2436.560 10.720 2436.880 11.040 ;
        RECT 2524.160 10.720 2524.480 11.040 ;
        RECT 2524.560 10.720 2524.880 11.040 ;
        RECT 2524.960 10.720 2525.280 11.040 ;
        RECT 2525.360 10.720 2525.680 11.040 ;
        RECT 2525.760 10.720 2526.080 11.040 ;
        RECT 2526.160 10.720 2526.480 11.040 ;
        RECT 2526.560 10.720 2526.880 11.040 ;
        RECT 2614.160 10.720 2614.480 11.040 ;
        RECT 2614.560 10.720 2614.880 11.040 ;
        RECT 2614.960 10.720 2615.280 11.040 ;
        RECT 2615.360 10.720 2615.680 11.040 ;
        RECT 2615.760 10.720 2616.080 11.040 ;
        RECT 2616.160 10.720 2616.480 11.040 ;
        RECT 2616.560 10.720 2616.880 11.040 ;
        RECT 2704.160 10.720 2704.480 11.040 ;
        RECT 2704.560 10.720 2704.880 11.040 ;
        RECT 2704.960 10.720 2705.280 11.040 ;
        RECT 2705.360 10.720 2705.680 11.040 ;
        RECT 2705.760 10.720 2706.080 11.040 ;
        RECT 2706.160 10.720 2706.480 11.040 ;
        RECT 2706.560 10.720 2706.880 11.040 ;
        RECT 2794.160 10.720 2794.480 11.040 ;
        RECT 2794.560 10.720 2794.880 11.040 ;
        RECT 2794.960 10.720 2795.280 11.040 ;
        RECT 2795.360 10.720 2795.680 11.040 ;
        RECT 2795.760 10.720 2796.080 11.040 ;
        RECT 2796.160 10.720 2796.480 11.040 ;
        RECT 2796.560 10.720 2796.880 11.040 ;
        RECT 2884.160 10.720 2884.480 11.040 ;
        RECT 2884.560 10.720 2884.880 11.040 ;
        RECT 2884.960 10.720 2885.280 11.040 ;
        RECT 2885.360 10.720 2885.680 11.040 ;
        RECT 2885.760 10.720 2886.080 11.040 ;
        RECT 2886.160 10.720 2886.480 11.040 ;
        RECT 2886.560 10.720 2886.880 11.040 ;
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 94.020 3506.300 97.020 3529.000 ;
        RECT 184.020 3506.300 187.020 3529.000 ;
        RECT 274.020 3506.300 277.020 3529.000 ;
        RECT 364.020 3506.300 367.020 3529.000 ;
        RECT 454.020 3506.300 457.020 3529.000 ;
        RECT 544.020 3506.300 547.020 3529.000 ;
        RECT 634.020 3506.300 637.020 3529.000 ;
        RECT 724.020 3506.300 727.020 3529.000 ;
        RECT 814.020 3506.300 817.020 3529.000 ;
        RECT 904.020 3506.300 907.020 3529.000 ;
        RECT 994.020 3506.300 997.020 3529.000 ;
        RECT 1084.020 3506.300 1087.020 3529.000 ;
        RECT 1174.020 3506.300 1177.020 3529.000 ;
        RECT 1264.020 3506.300 1267.020 3529.000 ;
        RECT 1354.020 3506.300 1357.020 3529.000 ;
        RECT 1444.020 3506.300 1447.020 3529.000 ;
        RECT 1534.020 3506.300 1537.020 3529.000 ;
        RECT 1624.020 3506.300 1627.020 3529.000 ;
        RECT 1714.020 3506.300 1717.020 3529.000 ;
        RECT 1804.020 3506.300 1807.020 3529.000 ;
        RECT 1894.020 3506.300 1897.020 3529.000 ;
        RECT 1984.020 3506.300 1987.020 3529.000 ;
        RECT 2074.020 3506.300 2077.020 3529.000 ;
        RECT 2164.020 3506.300 2167.020 3529.000 ;
        RECT 2254.020 3506.300 2257.020 3529.000 ;
        RECT 2344.020 3506.300 2347.020 3529.000 ;
        RECT 2434.020 3506.300 2437.020 3529.000 ;
        RECT 2524.020 3506.300 2527.020 3529.000 ;
        RECT 2614.020 3506.300 2617.020 3529.000 ;
        RECT 2704.020 3506.300 2707.020 3529.000 ;
        RECT 2794.020 3506.300 2797.020 3529.000 ;
        RECT 2884.020 3506.300 2887.020 3529.000 ;
        RECT 94.020 -9.320 97.020 13.700 ;
        RECT 184.020 -9.320 187.020 13.700 ;
        RECT 274.020 -9.320 277.020 13.700 ;
        RECT 364.020 -9.320 367.020 13.700 ;
        RECT 454.020 -9.320 457.020 13.700 ;
        RECT 544.020 -9.320 547.020 13.700 ;
        RECT 634.020 -9.320 637.020 13.700 ;
        RECT 724.020 -9.320 727.020 13.700 ;
        RECT 814.020 -9.320 817.020 13.700 ;
        RECT 904.020 -9.320 907.020 13.700 ;
        RECT 994.020 -9.320 997.020 13.700 ;
        RECT 1084.020 -9.320 1087.020 13.700 ;
        RECT 1174.020 -9.320 1177.020 13.700 ;
        RECT 1264.020 -9.320 1267.020 13.700 ;
        RECT 1354.020 -9.320 1357.020 13.700 ;
        RECT 1444.020 -9.320 1447.020 13.700 ;
        RECT 1534.020 -9.320 1537.020 13.700 ;
        RECT 1624.020 -9.320 1627.020 13.700 ;
        RECT 1714.020 -9.320 1717.020 13.700 ;
        RECT 1804.020 -9.320 1807.020 13.700 ;
        RECT 1894.020 -9.320 1897.020 13.700 ;
        RECT 1984.020 -9.320 1987.020 13.700 ;
        RECT 2074.020 -9.320 2077.020 13.700 ;
        RECT 2164.020 -9.320 2167.020 13.700 ;
        RECT 2254.020 -9.320 2257.020 13.700 ;
        RECT 2344.020 -9.320 2347.020 13.700 ;
        RECT 2434.020 -9.320 2437.020 13.700 ;
        RECT 2524.020 -9.320 2527.020 13.700 ;
        RECT 2614.020 -9.320 2617.020 13.700 ;
        RECT 2704.020 -9.320 2707.020 13.700 ;
        RECT 2794.020 -9.320 2797.020 13.700 ;
        RECT 2884.020 -9.320 2887.020 13.700 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3430.850 -7.890 3432.030 ;
        RECT -9.070 3429.250 -7.890 3430.430 ;
        RECT -9.070 3340.850 -7.890 3342.030 ;
        RECT -9.070 3339.250 -7.890 3340.430 ;
        RECT -9.070 3250.850 -7.890 3252.030 ;
        RECT -9.070 3249.250 -7.890 3250.430 ;
        RECT -9.070 3160.850 -7.890 3162.030 ;
        RECT -9.070 3159.250 -7.890 3160.430 ;
        RECT -9.070 3070.850 -7.890 3072.030 ;
        RECT -9.070 3069.250 -7.890 3070.430 ;
        RECT -9.070 2980.850 -7.890 2982.030 ;
        RECT -9.070 2979.250 -7.890 2980.430 ;
        RECT -9.070 2890.850 -7.890 2892.030 ;
        RECT -9.070 2889.250 -7.890 2890.430 ;
        RECT -9.070 2800.850 -7.890 2802.030 ;
        RECT -9.070 2799.250 -7.890 2800.430 ;
        RECT -9.070 2710.850 -7.890 2712.030 ;
        RECT -9.070 2709.250 -7.890 2710.430 ;
        RECT -9.070 2620.850 -7.890 2622.030 ;
        RECT -9.070 2619.250 -7.890 2620.430 ;
        RECT -9.070 2530.850 -7.890 2532.030 ;
        RECT -9.070 2529.250 -7.890 2530.430 ;
        RECT -9.070 2440.850 -7.890 2442.030 ;
        RECT -9.070 2439.250 -7.890 2440.430 ;
        RECT -9.070 2350.850 -7.890 2352.030 ;
        RECT -9.070 2349.250 -7.890 2350.430 ;
        RECT -9.070 2260.850 -7.890 2262.030 ;
        RECT -9.070 2259.250 -7.890 2260.430 ;
        RECT -9.070 2170.850 -7.890 2172.030 ;
        RECT -9.070 2169.250 -7.890 2170.430 ;
        RECT -9.070 2080.850 -7.890 2082.030 ;
        RECT -9.070 2079.250 -7.890 2080.430 ;
        RECT -9.070 1990.850 -7.890 1992.030 ;
        RECT -9.070 1989.250 -7.890 1990.430 ;
        RECT -9.070 1900.850 -7.890 1902.030 ;
        RECT -9.070 1899.250 -7.890 1900.430 ;
        RECT -9.070 1810.850 -7.890 1812.030 ;
        RECT -9.070 1809.250 -7.890 1810.430 ;
        RECT -9.070 1720.850 -7.890 1722.030 ;
        RECT -9.070 1719.250 -7.890 1720.430 ;
        RECT -9.070 1630.850 -7.890 1632.030 ;
        RECT -9.070 1629.250 -7.890 1630.430 ;
        RECT -9.070 1540.850 -7.890 1542.030 ;
        RECT -9.070 1539.250 -7.890 1540.430 ;
        RECT -9.070 1450.850 -7.890 1452.030 ;
        RECT -9.070 1449.250 -7.890 1450.430 ;
        RECT -9.070 1360.850 -7.890 1362.030 ;
        RECT -9.070 1359.250 -7.890 1360.430 ;
        RECT -9.070 1270.850 -7.890 1272.030 ;
        RECT -9.070 1269.250 -7.890 1270.430 ;
        RECT -9.070 1180.850 -7.890 1182.030 ;
        RECT -9.070 1179.250 -7.890 1180.430 ;
        RECT -9.070 1090.850 -7.890 1092.030 ;
        RECT -9.070 1089.250 -7.890 1090.430 ;
        RECT -9.070 1000.850 -7.890 1002.030 ;
        RECT -9.070 999.250 -7.890 1000.430 ;
        RECT -9.070 910.850 -7.890 912.030 ;
        RECT -9.070 909.250 -7.890 910.430 ;
        RECT -9.070 820.850 -7.890 822.030 ;
        RECT -9.070 819.250 -7.890 820.430 ;
        RECT -9.070 730.850 -7.890 732.030 ;
        RECT -9.070 729.250 -7.890 730.430 ;
        RECT -9.070 640.850 -7.890 642.030 ;
        RECT -9.070 639.250 -7.890 640.430 ;
        RECT -9.070 550.850 -7.890 552.030 ;
        RECT -9.070 549.250 -7.890 550.430 ;
        RECT -9.070 460.850 -7.890 462.030 ;
        RECT -9.070 459.250 -7.890 460.430 ;
        RECT -9.070 370.850 -7.890 372.030 ;
        RECT -9.070 369.250 -7.890 370.430 ;
        RECT -9.070 280.850 -7.890 282.030 ;
        RECT -9.070 279.250 -7.890 280.430 ;
        RECT -9.070 190.850 -7.890 192.030 ;
        RECT -9.070 189.250 -7.890 190.430 ;
        RECT -9.070 100.850 -7.890 102.030 ;
        RECT -9.070 99.250 -7.890 100.430 ;
        RECT -9.070 10.850 -7.890 12.030 ;
        RECT -9.070 9.250 -7.890 10.430 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 94.930 3523.010 96.110 3524.190 ;
        RECT 94.930 3521.410 96.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 274.930 3523.010 276.110 3524.190 ;
        RECT 274.930 3521.410 276.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 454.930 3523.010 456.110 3524.190 ;
        RECT 454.930 3521.410 456.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 634.930 3523.010 636.110 3524.190 ;
        RECT 634.930 3521.410 636.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 814.930 3523.010 816.110 3524.190 ;
        RECT 814.930 3521.410 816.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 994.930 3523.010 996.110 3524.190 ;
        RECT 994.930 3521.410 996.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1174.930 3523.010 1176.110 3524.190 ;
        RECT 1174.930 3521.410 1176.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1354.930 3523.010 1356.110 3524.190 ;
        RECT 1354.930 3521.410 1356.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1534.930 3523.010 1536.110 3524.190 ;
        RECT 1534.930 3521.410 1536.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1714.930 3523.010 1716.110 3524.190 ;
        RECT 1714.930 3521.410 1716.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1894.930 3523.010 1896.110 3524.190 ;
        RECT 1894.930 3521.410 1896.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2074.930 3523.010 2076.110 3524.190 ;
        RECT 2074.930 3521.410 2076.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2254.930 3523.010 2256.110 3524.190 ;
        RECT 2254.930 3521.410 2256.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2434.930 3523.010 2436.110 3524.190 ;
        RECT 2434.930 3521.410 2436.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2614.930 3523.010 2616.110 3524.190 ;
        RECT 2614.930 3521.410 2616.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2794.930 3523.010 2796.110 3524.190 ;
        RECT 2794.930 3521.410 2796.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 4.930 3430.850 6.110 3432.030 ;
        RECT 4.930 3429.250 6.110 3430.430 ;
        RECT 4.930 3340.850 6.110 3342.030 ;
        RECT 4.930 3339.250 6.110 3340.430 ;
        RECT 4.930 3250.850 6.110 3252.030 ;
        RECT 4.930 3249.250 6.110 3250.430 ;
        RECT 4.930 3160.850 6.110 3162.030 ;
        RECT 4.930 3159.250 6.110 3160.430 ;
        RECT 4.930 3070.850 6.110 3072.030 ;
        RECT 4.930 3069.250 6.110 3070.430 ;
        RECT 4.930 2980.850 6.110 2982.030 ;
        RECT 4.930 2979.250 6.110 2980.430 ;
        RECT 4.930 2890.850 6.110 2892.030 ;
        RECT 4.930 2889.250 6.110 2890.430 ;
        RECT 4.930 2800.850 6.110 2802.030 ;
        RECT 4.930 2799.250 6.110 2800.430 ;
        RECT 4.930 2710.850 6.110 2712.030 ;
        RECT 4.930 2709.250 6.110 2710.430 ;
        RECT 4.930 2620.850 6.110 2622.030 ;
        RECT 4.930 2619.250 6.110 2620.430 ;
        RECT 4.930 2530.850 6.110 2532.030 ;
        RECT 4.930 2529.250 6.110 2530.430 ;
        RECT 4.930 2440.850 6.110 2442.030 ;
        RECT 4.930 2439.250 6.110 2440.430 ;
        RECT 4.930 2350.850 6.110 2352.030 ;
        RECT 4.930 2349.250 6.110 2350.430 ;
        RECT 4.930 2260.850 6.110 2262.030 ;
        RECT 4.930 2259.250 6.110 2260.430 ;
        RECT 4.930 2170.850 6.110 2172.030 ;
        RECT 4.930 2169.250 6.110 2170.430 ;
        RECT 4.930 2080.850 6.110 2082.030 ;
        RECT 4.930 2079.250 6.110 2080.430 ;
        RECT 4.930 1990.850 6.110 1992.030 ;
        RECT 4.930 1989.250 6.110 1990.430 ;
        RECT 4.930 1900.850 6.110 1902.030 ;
        RECT 4.930 1899.250 6.110 1900.430 ;
        RECT 4.930 1810.850 6.110 1812.030 ;
        RECT 4.930 1809.250 6.110 1810.430 ;
        RECT 4.930 1720.850 6.110 1722.030 ;
        RECT 4.930 1719.250 6.110 1720.430 ;
        RECT 4.930 1630.850 6.110 1632.030 ;
        RECT 4.930 1629.250 6.110 1630.430 ;
        RECT 4.930 1540.850 6.110 1542.030 ;
        RECT 4.930 1539.250 6.110 1540.430 ;
        RECT 4.930 1450.850 6.110 1452.030 ;
        RECT 4.930 1449.250 6.110 1450.430 ;
        RECT 4.930 1360.850 6.110 1362.030 ;
        RECT 4.930 1359.250 6.110 1360.430 ;
        RECT 4.930 1270.850 6.110 1272.030 ;
        RECT 4.930 1269.250 6.110 1270.430 ;
        RECT 4.930 1180.850 6.110 1182.030 ;
        RECT 4.930 1179.250 6.110 1180.430 ;
        RECT 4.930 1090.850 6.110 1092.030 ;
        RECT 4.930 1089.250 6.110 1090.430 ;
        RECT 4.930 1000.850 6.110 1002.030 ;
        RECT 4.930 999.250 6.110 1000.430 ;
        RECT 4.930 910.850 6.110 912.030 ;
        RECT 4.930 909.250 6.110 910.430 ;
        RECT 4.930 820.850 6.110 822.030 ;
        RECT 4.930 819.250 6.110 820.430 ;
        RECT 4.930 730.850 6.110 732.030 ;
        RECT 4.930 729.250 6.110 730.430 ;
        RECT 4.930 640.850 6.110 642.030 ;
        RECT 4.930 639.250 6.110 640.430 ;
        RECT 4.930 550.850 6.110 552.030 ;
        RECT 4.930 549.250 6.110 550.430 ;
        RECT 4.930 460.850 6.110 462.030 ;
        RECT 4.930 459.250 6.110 460.430 ;
        RECT 4.930 370.850 6.110 372.030 ;
        RECT 4.930 369.250 6.110 370.430 ;
        RECT 4.930 280.850 6.110 282.030 ;
        RECT 4.930 279.250 6.110 280.430 ;
        RECT 4.930 190.850 6.110 192.030 ;
        RECT 4.930 189.250 6.110 190.430 ;
        RECT 4.930 100.850 6.110 102.030 ;
        RECT 4.930 99.250 6.110 100.430 ;
        RECT 2927.510 3430.850 2928.690 3432.030 ;
        RECT 2927.510 3429.250 2928.690 3430.430 ;
        RECT 2927.510 3340.850 2928.690 3342.030 ;
        RECT 2927.510 3339.250 2928.690 3340.430 ;
        RECT 2927.510 3250.850 2928.690 3252.030 ;
        RECT 2927.510 3249.250 2928.690 3250.430 ;
        RECT 2927.510 3160.850 2928.690 3162.030 ;
        RECT 2927.510 3159.250 2928.690 3160.430 ;
        RECT 2927.510 3070.850 2928.690 3072.030 ;
        RECT 2927.510 3069.250 2928.690 3070.430 ;
        RECT 2927.510 2980.850 2928.690 2982.030 ;
        RECT 2927.510 2979.250 2928.690 2980.430 ;
        RECT 2927.510 2890.850 2928.690 2892.030 ;
        RECT 2927.510 2889.250 2928.690 2890.430 ;
        RECT 2927.510 2800.850 2928.690 2802.030 ;
        RECT 2927.510 2799.250 2928.690 2800.430 ;
        RECT 2927.510 2710.850 2928.690 2712.030 ;
        RECT 2927.510 2709.250 2928.690 2710.430 ;
        RECT 2927.510 2620.850 2928.690 2622.030 ;
        RECT 2927.510 2619.250 2928.690 2620.430 ;
        RECT 2927.510 2530.850 2928.690 2532.030 ;
        RECT 2927.510 2529.250 2928.690 2530.430 ;
        RECT 2927.510 2440.850 2928.690 2442.030 ;
        RECT 2927.510 2439.250 2928.690 2440.430 ;
        RECT 2927.510 2350.850 2928.690 2352.030 ;
        RECT 2927.510 2349.250 2928.690 2350.430 ;
        RECT 2927.510 2260.850 2928.690 2262.030 ;
        RECT 2927.510 2259.250 2928.690 2260.430 ;
        RECT 2927.510 2170.850 2928.690 2172.030 ;
        RECT 2927.510 2169.250 2928.690 2170.430 ;
        RECT 2927.510 2080.850 2928.690 2082.030 ;
        RECT 2927.510 2079.250 2928.690 2080.430 ;
        RECT 2927.510 1990.850 2928.690 1992.030 ;
        RECT 2927.510 1989.250 2928.690 1990.430 ;
        RECT 2927.510 1900.850 2928.690 1902.030 ;
        RECT 2927.510 1899.250 2928.690 1900.430 ;
        RECT 2927.510 1810.850 2928.690 1812.030 ;
        RECT 2927.510 1809.250 2928.690 1810.430 ;
        RECT 2927.510 1720.850 2928.690 1722.030 ;
        RECT 2927.510 1719.250 2928.690 1720.430 ;
        RECT 2927.510 1630.850 2928.690 1632.030 ;
        RECT 2927.510 1629.250 2928.690 1630.430 ;
        RECT 2927.510 1540.850 2928.690 1542.030 ;
        RECT 2927.510 1539.250 2928.690 1540.430 ;
        RECT 2927.510 1450.850 2928.690 1452.030 ;
        RECT 2927.510 1449.250 2928.690 1450.430 ;
        RECT 2927.510 1360.850 2928.690 1362.030 ;
        RECT 2927.510 1359.250 2928.690 1360.430 ;
        RECT 2927.510 1270.850 2928.690 1272.030 ;
        RECT 2927.510 1269.250 2928.690 1270.430 ;
        RECT 2927.510 1180.850 2928.690 1182.030 ;
        RECT 2927.510 1179.250 2928.690 1180.430 ;
        RECT 2927.510 1090.850 2928.690 1092.030 ;
        RECT 2927.510 1089.250 2928.690 1090.430 ;
        RECT 2927.510 1000.850 2928.690 1002.030 ;
        RECT 2927.510 999.250 2928.690 1000.430 ;
        RECT 2927.510 910.850 2928.690 912.030 ;
        RECT 2927.510 909.250 2928.690 910.430 ;
        RECT 2927.510 820.850 2928.690 822.030 ;
        RECT 2927.510 819.250 2928.690 820.430 ;
        RECT 2927.510 730.850 2928.690 732.030 ;
        RECT 2927.510 729.250 2928.690 730.430 ;
        RECT 2927.510 640.850 2928.690 642.030 ;
        RECT 2927.510 639.250 2928.690 640.430 ;
        RECT 2927.510 550.850 2928.690 552.030 ;
        RECT 2927.510 549.250 2928.690 550.430 ;
        RECT 2927.510 460.850 2928.690 462.030 ;
        RECT 2927.510 459.250 2928.690 460.430 ;
        RECT 2927.510 370.850 2928.690 372.030 ;
        RECT 2927.510 369.250 2928.690 370.430 ;
        RECT 2927.510 280.850 2928.690 282.030 ;
        RECT 2927.510 279.250 2928.690 280.430 ;
        RECT 2927.510 190.850 2928.690 192.030 ;
        RECT 2927.510 189.250 2928.690 190.430 ;
        RECT 2927.510 100.850 2928.690 102.030 ;
        RECT 2927.510 99.250 2928.690 100.430 ;
        RECT 4.930 10.850 6.110 12.030 ;
        RECT 4.930 9.250 6.110 10.430 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 94.930 10.850 96.110 12.030 ;
        RECT 94.930 9.250 96.110 10.430 ;
        RECT 94.930 -2.910 96.110 -1.730 ;
        RECT 94.930 -4.510 96.110 -3.330 ;
        RECT 184.930 10.850 186.110 12.030 ;
        RECT 184.930 9.250 186.110 10.430 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 274.930 10.850 276.110 12.030 ;
        RECT 274.930 9.250 276.110 10.430 ;
        RECT 274.930 -2.910 276.110 -1.730 ;
        RECT 274.930 -4.510 276.110 -3.330 ;
        RECT 364.930 10.850 366.110 12.030 ;
        RECT 364.930 9.250 366.110 10.430 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 454.930 10.850 456.110 12.030 ;
        RECT 454.930 9.250 456.110 10.430 ;
        RECT 454.930 -2.910 456.110 -1.730 ;
        RECT 454.930 -4.510 456.110 -3.330 ;
        RECT 544.930 10.850 546.110 12.030 ;
        RECT 544.930 9.250 546.110 10.430 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 634.930 10.850 636.110 12.030 ;
        RECT 634.930 9.250 636.110 10.430 ;
        RECT 634.930 -2.910 636.110 -1.730 ;
        RECT 634.930 -4.510 636.110 -3.330 ;
        RECT 724.930 10.850 726.110 12.030 ;
        RECT 724.930 9.250 726.110 10.430 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 814.930 10.850 816.110 12.030 ;
        RECT 814.930 9.250 816.110 10.430 ;
        RECT 814.930 -2.910 816.110 -1.730 ;
        RECT 814.930 -4.510 816.110 -3.330 ;
        RECT 904.930 10.850 906.110 12.030 ;
        RECT 904.930 9.250 906.110 10.430 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 994.930 10.850 996.110 12.030 ;
        RECT 994.930 9.250 996.110 10.430 ;
        RECT 994.930 -2.910 996.110 -1.730 ;
        RECT 994.930 -4.510 996.110 -3.330 ;
        RECT 1084.930 10.850 1086.110 12.030 ;
        RECT 1084.930 9.250 1086.110 10.430 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1174.930 10.850 1176.110 12.030 ;
        RECT 1174.930 9.250 1176.110 10.430 ;
        RECT 1174.930 -2.910 1176.110 -1.730 ;
        RECT 1174.930 -4.510 1176.110 -3.330 ;
        RECT 1264.930 10.850 1266.110 12.030 ;
        RECT 1264.930 9.250 1266.110 10.430 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1354.930 10.850 1356.110 12.030 ;
        RECT 1354.930 9.250 1356.110 10.430 ;
        RECT 1354.930 -2.910 1356.110 -1.730 ;
        RECT 1354.930 -4.510 1356.110 -3.330 ;
        RECT 1444.930 10.850 1446.110 12.030 ;
        RECT 1444.930 9.250 1446.110 10.430 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1534.930 10.850 1536.110 12.030 ;
        RECT 1534.930 9.250 1536.110 10.430 ;
        RECT 1534.930 -2.910 1536.110 -1.730 ;
        RECT 1534.930 -4.510 1536.110 -3.330 ;
        RECT 1624.930 10.850 1626.110 12.030 ;
        RECT 1624.930 9.250 1626.110 10.430 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1714.930 10.850 1716.110 12.030 ;
        RECT 1714.930 9.250 1716.110 10.430 ;
        RECT 1714.930 -2.910 1716.110 -1.730 ;
        RECT 1714.930 -4.510 1716.110 -3.330 ;
        RECT 1804.930 10.850 1806.110 12.030 ;
        RECT 1804.930 9.250 1806.110 10.430 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1894.930 10.850 1896.110 12.030 ;
        RECT 1894.930 9.250 1896.110 10.430 ;
        RECT 1894.930 -2.910 1896.110 -1.730 ;
        RECT 1894.930 -4.510 1896.110 -3.330 ;
        RECT 1984.930 10.850 1986.110 12.030 ;
        RECT 1984.930 9.250 1986.110 10.430 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2074.930 10.850 2076.110 12.030 ;
        RECT 2074.930 9.250 2076.110 10.430 ;
        RECT 2074.930 -2.910 2076.110 -1.730 ;
        RECT 2074.930 -4.510 2076.110 -3.330 ;
        RECT 2164.930 10.850 2166.110 12.030 ;
        RECT 2164.930 9.250 2166.110 10.430 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2254.930 10.850 2256.110 12.030 ;
        RECT 2254.930 9.250 2256.110 10.430 ;
        RECT 2254.930 -2.910 2256.110 -1.730 ;
        RECT 2254.930 -4.510 2256.110 -3.330 ;
        RECT 2344.930 10.850 2346.110 12.030 ;
        RECT 2344.930 9.250 2346.110 10.430 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2434.930 10.850 2436.110 12.030 ;
        RECT 2434.930 9.250 2436.110 10.430 ;
        RECT 2434.930 -2.910 2436.110 -1.730 ;
        RECT 2434.930 -4.510 2436.110 -3.330 ;
        RECT 2524.930 10.850 2526.110 12.030 ;
        RECT 2524.930 9.250 2526.110 10.430 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2614.930 10.850 2616.110 12.030 ;
        RECT 2614.930 9.250 2616.110 10.430 ;
        RECT 2614.930 -2.910 2616.110 -1.730 ;
        RECT 2614.930 -4.510 2616.110 -3.330 ;
        RECT 2704.930 10.850 2706.110 12.030 ;
        RECT 2704.930 9.250 2706.110 10.430 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2794.930 10.850 2796.110 12.030 ;
        RECT 2794.930 9.250 2796.110 10.430 ;
        RECT 2794.930 -2.910 2796.110 -1.730 ;
        RECT 2794.930 -4.510 2796.110 -3.330 ;
        RECT 2884.930 10.850 2886.110 12.030 ;
        RECT 2884.930 9.250 2886.110 10.430 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 10.850 2928.690 12.030 ;
        RECT 2927.510 9.250 2928.690 10.430 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 94.020 3524.300 97.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 274.020 3524.300 277.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 454.020 3524.300 457.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 634.020 3524.300 637.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 814.020 3524.300 817.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 994.020 3524.300 997.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1174.020 3524.300 1177.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1354.020 3524.300 1357.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1534.020 3524.300 1537.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1714.020 3524.300 1717.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1894.020 3524.300 1897.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2074.020 3524.300 2077.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2254.020 3524.300 2257.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2434.020 3524.300 2437.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2614.020 3524.300 2617.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2794.020 3524.300 2797.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 94.020 3521.290 97.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 274.020 3521.290 277.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 454.020 3521.290 457.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 634.020 3521.290 637.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 814.020 3521.290 817.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 994.020 3521.290 997.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1174.020 3521.290 1177.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1354.020 3521.290 1357.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1534.020 3521.290 1537.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1714.020 3521.290 1717.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1894.020 3521.290 1897.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2074.020 3521.290 2077.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2254.020 3521.290 2257.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2434.020 3521.290 2437.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2614.020 3521.290 2617.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2794.020 3521.290 2797.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.140 -6.980 3432.150 ;
        RECT 4.020 3432.140 7.020 3432.150 ;
        RECT 2926.600 3432.140 2929.600 3432.150 ;
        RECT -14.680 3429.140 13.700 3432.140 ;
        RECT 2906.300 3429.140 2934.300 3432.140 ;
        RECT -9.980 3429.130 -6.980 3429.140 ;
        RECT 4.020 3429.130 7.020 3429.140 ;
        RECT 2926.600 3429.130 2929.600 3429.140 ;
        RECT -9.980 3342.140 -6.980 3342.150 ;
        RECT 4.020 3342.140 7.020 3342.150 ;
        RECT 2926.600 3342.140 2929.600 3342.150 ;
        RECT -14.680 3339.140 13.700 3342.140 ;
        RECT 2906.300 3339.140 2934.300 3342.140 ;
        RECT -9.980 3339.130 -6.980 3339.140 ;
        RECT 4.020 3339.130 7.020 3339.140 ;
        RECT 2926.600 3339.130 2929.600 3339.140 ;
        RECT -9.980 3252.140 -6.980 3252.150 ;
        RECT 4.020 3252.140 7.020 3252.150 ;
        RECT 2926.600 3252.140 2929.600 3252.150 ;
        RECT -14.680 3249.140 13.700 3252.140 ;
        RECT 2906.300 3249.140 2934.300 3252.140 ;
        RECT -9.980 3249.130 -6.980 3249.140 ;
        RECT 4.020 3249.130 7.020 3249.140 ;
        RECT 2926.600 3249.130 2929.600 3249.140 ;
        RECT -9.980 3162.140 -6.980 3162.150 ;
        RECT 4.020 3162.140 7.020 3162.150 ;
        RECT 2926.600 3162.140 2929.600 3162.150 ;
        RECT -14.680 3159.140 13.700 3162.140 ;
        RECT 2906.300 3159.140 2934.300 3162.140 ;
        RECT -9.980 3159.130 -6.980 3159.140 ;
        RECT 4.020 3159.130 7.020 3159.140 ;
        RECT 2926.600 3159.130 2929.600 3159.140 ;
        RECT -9.980 3072.140 -6.980 3072.150 ;
        RECT 4.020 3072.140 7.020 3072.150 ;
        RECT 2926.600 3072.140 2929.600 3072.150 ;
        RECT -14.680 3069.140 13.700 3072.140 ;
        RECT 2906.300 3069.140 2934.300 3072.140 ;
        RECT -9.980 3069.130 -6.980 3069.140 ;
        RECT 4.020 3069.130 7.020 3069.140 ;
        RECT 2926.600 3069.130 2929.600 3069.140 ;
        RECT -9.980 2982.140 -6.980 2982.150 ;
        RECT 4.020 2982.140 7.020 2982.150 ;
        RECT 2926.600 2982.140 2929.600 2982.150 ;
        RECT -14.680 2979.140 13.700 2982.140 ;
        RECT 2906.300 2979.140 2934.300 2982.140 ;
        RECT -9.980 2979.130 -6.980 2979.140 ;
        RECT 4.020 2979.130 7.020 2979.140 ;
        RECT 2926.600 2979.130 2929.600 2979.140 ;
        RECT -9.980 2892.140 -6.980 2892.150 ;
        RECT 4.020 2892.140 7.020 2892.150 ;
        RECT 2926.600 2892.140 2929.600 2892.150 ;
        RECT -14.680 2889.140 13.700 2892.140 ;
        RECT 2906.300 2889.140 2934.300 2892.140 ;
        RECT -9.980 2889.130 -6.980 2889.140 ;
        RECT 4.020 2889.130 7.020 2889.140 ;
        RECT 2926.600 2889.130 2929.600 2889.140 ;
        RECT -9.980 2802.140 -6.980 2802.150 ;
        RECT 4.020 2802.140 7.020 2802.150 ;
        RECT 2926.600 2802.140 2929.600 2802.150 ;
        RECT -14.680 2799.140 13.700 2802.140 ;
        RECT 2906.300 2799.140 2934.300 2802.140 ;
        RECT -9.980 2799.130 -6.980 2799.140 ;
        RECT 4.020 2799.130 7.020 2799.140 ;
        RECT 2926.600 2799.130 2929.600 2799.140 ;
        RECT -9.980 2712.140 -6.980 2712.150 ;
        RECT 4.020 2712.140 7.020 2712.150 ;
        RECT 2926.600 2712.140 2929.600 2712.150 ;
        RECT -14.680 2709.140 13.700 2712.140 ;
        RECT 2906.300 2709.140 2934.300 2712.140 ;
        RECT -9.980 2709.130 -6.980 2709.140 ;
        RECT 4.020 2709.130 7.020 2709.140 ;
        RECT 2926.600 2709.130 2929.600 2709.140 ;
        RECT -9.980 2622.140 -6.980 2622.150 ;
        RECT 4.020 2622.140 7.020 2622.150 ;
        RECT 2926.600 2622.140 2929.600 2622.150 ;
        RECT -14.680 2619.140 13.700 2622.140 ;
        RECT 2906.300 2619.140 2934.300 2622.140 ;
        RECT -9.980 2619.130 -6.980 2619.140 ;
        RECT 4.020 2619.130 7.020 2619.140 ;
        RECT 2926.600 2619.130 2929.600 2619.140 ;
        RECT -9.980 2532.140 -6.980 2532.150 ;
        RECT 4.020 2532.140 7.020 2532.150 ;
        RECT 2926.600 2532.140 2929.600 2532.150 ;
        RECT -14.680 2529.140 13.700 2532.140 ;
        RECT 2906.300 2529.140 2934.300 2532.140 ;
        RECT -9.980 2529.130 -6.980 2529.140 ;
        RECT 4.020 2529.130 7.020 2529.140 ;
        RECT 2926.600 2529.130 2929.600 2529.140 ;
        RECT -9.980 2442.140 -6.980 2442.150 ;
        RECT 4.020 2442.140 7.020 2442.150 ;
        RECT 2926.600 2442.140 2929.600 2442.150 ;
        RECT -14.680 2439.140 13.700 2442.140 ;
        RECT 2906.300 2439.140 2934.300 2442.140 ;
        RECT -9.980 2439.130 -6.980 2439.140 ;
        RECT 4.020 2439.130 7.020 2439.140 ;
        RECT 2926.600 2439.130 2929.600 2439.140 ;
        RECT -9.980 2352.140 -6.980 2352.150 ;
        RECT 4.020 2352.140 7.020 2352.150 ;
        RECT 2926.600 2352.140 2929.600 2352.150 ;
        RECT -14.680 2349.140 13.700 2352.140 ;
        RECT 2906.300 2349.140 2934.300 2352.140 ;
        RECT -9.980 2349.130 -6.980 2349.140 ;
        RECT 4.020 2349.130 7.020 2349.140 ;
        RECT 2926.600 2349.130 2929.600 2349.140 ;
        RECT -9.980 2262.140 -6.980 2262.150 ;
        RECT 4.020 2262.140 7.020 2262.150 ;
        RECT 2926.600 2262.140 2929.600 2262.150 ;
        RECT -14.680 2259.140 13.700 2262.140 ;
        RECT 2906.300 2259.140 2934.300 2262.140 ;
        RECT -9.980 2259.130 -6.980 2259.140 ;
        RECT 4.020 2259.130 7.020 2259.140 ;
        RECT 2926.600 2259.130 2929.600 2259.140 ;
        RECT -9.980 2172.140 -6.980 2172.150 ;
        RECT 4.020 2172.140 7.020 2172.150 ;
        RECT 2926.600 2172.140 2929.600 2172.150 ;
        RECT -14.680 2169.140 13.700 2172.140 ;
        RECT 2906.300 2169.140 2934.300 2172.140 ;
        RECT -9.980 2169.130 -6.980 2169.140 ;
        RECT 4.020 2169.130 7.020 2169.140 ;
        RECT 2926.600 2169.130 2929.600 2169.140 ;
        RECT -9.980 2082.140 -6.980 2082.150 ;
        RECT 4.020 2082.140 7.020 2082.150 ;
        RECT 2926.600 2082.140 2929.600 2082.150 ;
        RECT -14.680 2079.140 13.700 2082.140 ;
        RECT 2906.300 2079.140 2934.300 2082.140 ;
        RECT -9.980 2079.130 -6.980 2079.140 ;
        RECT 4.020 2079.130 7.020 2079.140 ;
        RECT 2926.600 2079.130 2929.600 2079.140 ;
        RECT -9.980 1992.140 -6.980 1992.150 ;
        RECT 4.020 1992.140 7.020 1992.150 ;
        RECT 2926.600 1992.140 2929.600 1992.150 ;
        RECT -14.680 1989.140 13.700 1992.140 ;
        RECT 2906.300 1989.140 2934.300 1992.140 ;
        RECT -9.980 1989.130 -6.980 1989.140 ;
        RECT 4.020 1989.130 7.020 1989.140 ;
        RECT 2926.600 1989.130 2929.600 1989.140 ;
        RECT -9.980 1902.140 -6.980 1902.150 ;
        RECT 4.020 1902.140 7.020 1902.150 ;
        RECT 2926.600 1902.140 2929.600 1902.150 ;
        RECT -14.680 1899.140 13.700 1902.140 ;
        RECT 2906.300 1899.140 2934.300 1902.140 ;
        RECT -9.980 1899.130 -6.980 1899.140 ;
        RECT 4.020 1899.130 7.020 1899.140 ;
        RECT 2926.600 1899.130 2929.600 1899.140 ;
        RECT -9.980 1812.140 -6.980 1812.150 ;
        RECT 4.020 1812.140 7.020 1812.150 ;
        RECT 2926.600 1812.140 2929.600 1812.150 ;
        RECT -14.680 1809.140 13.700 1812.140 ;
        RECT 2906.300 1809.140 2934.300 1812.140 ;
        RECT -9.980 1809.130 -6.980 1809.140 ;
        RECT 4.020 1809.130 7.020 1809.140 ;
        RECT 2926.600 1809.130 2929.600 1809.140 ;
        RECT -9.980 1722.140 -6.980 1722.150 ;
        RECT 4.020 1722.140 7.020 1722.150 ;
        RECT 2926.600 1722.140 2929.600 1722.150 ;
        RECT -14.680 1719.140 13.700 1722.140 ;
        RECT 2906.300 1719.140 2934.300 1722.140 ;
        RECT -9.980 1719.130 -6.980 1719.140 ;
        RECT 4.020 1719.130 7.020 1719.140 ;
        RECT 2926.600 1719.130 2929.600 1719.140 ;
        RECT -9.980 1632.140 -6.980 1632.150 ;
        RECT 4.020 1632.140 7.020 1632.150 ;
        RECT 2926.600 1632.140 2929.600 1632.150 ;
        RECT -14.680 1629.140 13.700 1632.140 ;
        RECT 2906.300 1629.140 2934.300 1632.140 ;
        RECT -9.980 1629.130 -6.980 1629.140 ;
        RECT 4.020 1629.130 7.020 1629.140 ;
        RECT 2926.600 1629.130 2929.600 1629.140 ;
        RECT -9.980 1542.140 -6.980 1542.150 ;
        RECT 4.020 1542.140 7.020 1542.150 ;
        RECT 2926.600 1542.140 2929.600 1542.150 ;
        RECT -14.680 1539.140 13.700 1542.140 ;
        RECT 2906.300 1539.140 2934.300 1542.140 ;
        RECT -9.980 1539.130 -6.980 1539.140 ;
        RECT 4.020 1539.130 7.020 1539.140 ;
        RECT 2926.600 1539.130 2929.600 1539.140 ;
        RECT -9.980 1452.140 -6.980 1452.150 ;
        RECT 4.020 1452.140 7.020 1452.150 ;
        RECT 2926.600 1452.140 2929.600 1452.150 ;
        RECT -14.680 1449.140 13.700 1452.140 ;
        RECT 2906.300 1449.140 2934.300 1452.140 ;
        RECT -9.980 1449.130 -6.980 1449.140 ;
        RECT 4.020 1449.130 7.020 1449.140 ;
        RECT 2926.600 1449.130 2929.600 1449.140 ;
        RECT -9.980 1362.140 -6.980 1362.150 ;
        RECT 4.020 1362.140 7.020 1362.150 ;
        RECT 2926.600 1362.140 2929.600 1362.150 ;
        RECT -14.680 1359.140 13.700 1362.140 ;
        RECT 2906.300 1359.140 2934.300 1362.140 ;
        RECT -9.980 1359.130 -6.980 1359.140 ;
        RECT 4.020 1359.130 7.020 1359.140 ;
        RECT 2926.600 1359.130 2929.600 1359.140 ;
        RECT -9.980 1272.140 -6.980 1272.150 ;
        RECT 4.020 1272.140 7.020 1272.150 ;
        RECT 2926.600 1272.140 2929.600 1272.150 ;
        RECT -14.680 1269.140 13.700 1272.140 ;
        RECT 2906.300 1269.140 2934.300 1272.140 ;
        RECT -9.980 1269.130 -6.980 1269.140 ;
        RECT 4.020 1269.130 7.020 1269.140 ;
        RECT 2926.600 1269.130 2929.600 1269.140 ;
        RECT -9.980 1182.140 -6.980 1182.150 ;
        RECT 4.020 1182.140 7.020 1182.150 ;
        RECT 2926.600 1182.140 2929.600 1182.150 ;
        RECT -14.680 1179.140 13.700 1182.140 ;
        RECT 2906.300 1179.140 2934.300 1182.140 ;
        RECT -9.980 1179.130 -6.980 1179.140 ;
        RECT 4.020 1179.130 7.020 1179.140 ;
        RECT 2926.600 1179.130 2929.600 1179.140 ;
        RECT -9.980 1092.140 -6.980 1092.150 ;
        RECT 4.020 1092.140 7.020 1092.150 ;
        RECT 2926.600 1092.140 2929.600 1092.150 ;
        RECT -14.680 1089.140 13.700 1092.140 ;
        RECT 2906.300 1089.140 2934.300 1092.140 ;
        RECT -9.980 1089.130 -6.980 1089.140 ;
        RECT 4.020 1089.130 7.020 1089.140 ;
        RECT 2926.600 1089.130 2929.600 1089.140 ;
        RECT -9.980 1002.140 -6.980 1002.150 ;
        RECT 4.020 1002.140 7.020 1002.150 ;
        RECT 2926.600 1002.140 2929.600 1002.150 ;
        RECT -14.680 999.140 13.700 1002.140 ;
        RECT 2906.300 999.140 2934.300 1002.140 ;
        RECT -9.980 999.130 -6.980 999.140 ;
        RECT 4.020 999.130 7.020 999.140 ;
        RECT 2926.600 999.130 2929.600 999.140 ;
        RECT -9.980 912.140 -6.980 912.150 ;
        RECT 4.020 912.140 7.020 912.150 ;
        RECT 2926.600 912.140 2929.600 912.150 ;
        RECT -14.680 909.140 13.700 912.140 ;
        RECT 2906.300 909.140 2934.300 912.140 ;
        RECT -9.980 909.130 -6.980 909.140 ;
        RECT 4.020 909.130 7.020 909.140 ;
        RECT 2926.600 909.130 2929.600 909.140 ;
        RECT -9.980 822.140 -6.980 822.150 ;
        RECT 4.020 822.140 7.020 822.150 ;
        RECT 2926.600 822.140 2929.600 822.150 ;
        RECT -14.680 819.140 13.700 822.140 ;
        RECT 2906.300 819.140 2934.300 822.140 ;
        RECT -9.980 819.130 -6.980 819.140 ;
        RECT 4.020 819.130 7.020 819.140 ;
        RECT 2926.600 819.130 2929.600 819.140 ;
        RECT -9.980 732.140 -6.980 732.150 ;
        RECT 4.020 732.140 7.020 732.150 ;
        RECT 2926.600 732.140 2929.600 732.150 ;
        RECT -14.680 729.140 13.700 732.140 ;
        RECT 2906.300 729.140 2934.300 732.140 ;
        RECT -9.980 729.130 -6.980 729.140 ;
        RECT 4.020 729.130 7.020 729.140 ;
        RECT 2926.600 729.130 2929.600 729.140 ;
        RECT -9.980 642.140 -6.980 642.150 ;
        RECT 4.020 642.140 7.020 642.150 ;
        RECT 2926.600 642.140 2929.600 642.150 ;
        RECT -14.680 639.140 13.700 642.140 ;
        RECT 2906.300 639.140 2934.300 642.140 ;
        RECT -9.980 639.130 -6.980 639.140 ;
        RECT 4.020 639.130 7.020 639.140 ;
        RECT 2926.600 639.130 2929.600 639.140 ;
        RECT -9.980 552.140 -6.980 552.150 ;
        RECT 4.020 552.140 7.020 552.150 ;
        RECT 2926.600 552.140 2929.600 552.150 ;
        RECT -14.680 549.140 13.700 552.140 ;
        RECT 2906.300 549.140 2934.300 552.140 ;
        RECT -9.980 549.130 -6.980 549.140 ;
        RECT 4.020 549.130 7.020 549.140 ;
        RECT 2926.600 549.130 2929.600 549.140 ;
        RECT -9.980 462.140 -6.980 462.150 ;
        RECT 4.020 462.140 7.020 462.150 ;
        RECT 2926.600 462.140 2929.600 462.150 ;
        RECT -14.680 459.140 13.700 462.140 ;
        RECT 2906.300 459.140 2934.300 462.140 ;
        RECT -9.980 459.130 -6.980 459.140 ;
        RECT 4.020 459.130 7.020 459.140 ;
        RECT 2926.600 459.130 2929.600 459.140 ;
        RECT -9.980 372.140 -6.980 372.150 ;
        RECT 4.020 372.140 7.020 372.150 ;
        RECT 2926.600 372.140 2929.600 372.150 ;
        RECT -14.680 369.140 13.700 372.140 ;
        RECT 2906.300 369.140 2934.300 372.140 ;
        RECT -9.980 369.130 -6.980 369.140 ;
        RECT 4.020 369.130 7.020 369.140 ;
        RECT 2926.600 369.130 2929.600 369.140 ;
        RECT -9.980 282.140 -6.980 282.150 ;
        RECT 4.020 282.140 7.020 282.150 ;
        RECT 2926.600 282.140 2929.600 282.150 ;
        RECT -14.680 279.140 13.700 282.140 ;
        RECT 2906.300 279.140 2934.300 282.140 ;
        RECT -9.980 279.130 -6.980 279.140 ;
        RECT 4.020 279.130 7.020 279.140 ;
        RECT 2926.600 279.130 2929.600 279.140 ;
        RECT -9.980 192.140 -6.980 192.150 ;
        RECT 4.020 192.140 7.020 192.150 ;
        RECT 2926.600 192.140 2929.600 192.150 ;
        RECT -14.680 189.140 13.700 192.140 ;
        RECT 2906.300 189.140 2934.300 192.140 ;
        RECT -9.980 189.130 -6.980 189.140 ;
        RECT 4.020 189.130 7.020 189.140 ;
        RECT 2926.600 189.130 2929.600 189.140 ;
        RECT -9.980 102.140 -6.980 102.150 ;
        RECT 4.020 102.140 7.020 102.150 ;
        RECT 2926.600 102.140 2929.600 102.150 ;
        RECT -14.680 99.140 13.700 102.140 ;
        RECT 2906.300 99.140 2934.300 102.140 ;
        RECT -9.980 99.130 -6.980 99.140 ;
        RECT 4.020 99.130 7.020 99.140 ;
        RECT 2926.600 99.130 2929.600 99.140 ;
        RECT -9.980 12.140 -6.980 12.150 ;
        RECT 4.020 12.140 7.020 12.150 ;
        RECT 94.020 12.140 97.020 12.150 ;
        RECT 184.020 12.140 187.020 12.150 ;
        RECT 274.020 12.140 277.020 12.150 ;
        RECT 364.020 12.140 367.020 12.150 ;
        RECT 454.020 12.140 457.020 12.150 ;
        RECT 544.020 12.140 547.020 12.150 ;
        RECT 634.020 12.140 637.020 12.150 ;
        RECT 724.020 12.140 727.020 12.150 ;
        RECT 814.020 12.140 817.020 12.150 ;
        RECT 904.020 12.140 907.020 12.150 ;
        RECT 994.020 12.140 997.020 12.150 ;
        RECT 1084.020 12.140 1087.020 12.150 ;
        RECT 1174.020 12.140 1177.020 12.150 ;
        RECT 1264.020 12.140 1267.020 12.150 ;
        RECT 1354.020 12.140 1357.020 12.150 ;
        RECT 1444.020 12.140 1447.020 12.150 ;
        RECT 1534.020 12.140 1537.020 12.150 ;
        RECT 1624.020 12.140 1627.020 12.150 ;
        RECT 1714.020 12.140 1717.020 12.150 ;
        RECT 1804.020 12.140 1807.020 12.150 ;
        RECT 1894.020 12.140 1897.020 12.150 ;
        RECT 1984.020 12.140 1987.020 12.150 ;
        RECT 2074.020 12.140 2077.020 12.150 ;
        RECT 2164.020 12.140 2167.020 12.150 ;
        RECT 2254.020 12.140 2257.020 12.150 ;
        RECT 2344.020 12.140 2347.020 12.150 ;
        RECT 2434.020 12.140 2437.020 12.150 ;
        RECT 2524.020 12.140 2527.020 12.150 ;
        RECT 2614.020 12.140 2617.020 12.150 ;
        RECT 2704.020 12.140 2707.020 12.150 ;
        RECT 2794.020 12.140 2797.020 12.150 ;
        RECT 2884.020 12.140 2887.020 12.150 ;
        RECT 2926.600 12.140 2929.600 12.150 ;
        RECT -14.680 9.140 2934.300 12.140 ;
        RECT -9.980 9.130 -6.980 9.140 ;
        RECT 4.020 9.130 7.020 9.140 ;
        RECT 94.020 9.130 97.020 9.140 ;
        RECT 184.020 9.130 187.020 9.140 ;
        RECT 274.020 9.130 277.020 9.140 ;
        RECT 364.020 9.130 367.020 9.140 ;
        RECT 454.020 9.130 457.020 9.140 ;
        RECT 544.020 9.130 547.020 9.140 ;
        RECT 634.020 9.130 637.020 9.140 ;
        RECT 724.020 9.130 727.020 9.140 ;
        RECT 814.020 9.130 817.020 9.140 ;
        RECT 904.020 9.130 907.020 9.140 ;
        RECT 994.020 9.130 997.020 9.140 ;
        RECT 1084.020 9.130 1087.020 9.140 ;
        RECT 1174.020 9.130 1177.020 9.140 ;
        RECT 1264.020 9.130 1267.020 9.140 ;
        RECT 1354.020 9.130 1357.020 9.140 ;
        RECT 1444.020 9.130 1447.020 9.140 ;
        RECT 1534.020 9.130 1537.020 9.140 ;
        RECT 1624.020 9.130 1627.020 9.140 ;
        RECT 1714.020 9.130 1717.020 9.140 ;
        RECT 1804.020 9.130 1807.020 9.140 ;
        RECT 1894.020 9.130 1897.020 9.140 ;
        RECT 1984.020 9.130 1987.020 9.140 ;
        RECT 2074.020 9.130 2077.020 9.140 ;
        RECT 2164.020 9.130 2167.020 9.140 ;
        RECT 2254.020 9.130 2257.020 9.140 ;
        RECT 2344.020 9.130 2347.020 9.140 ;
        RECT 2434.020 9.130 2437.020 9.140 ;
        RECT 2524.020 9.130 2527.020 9.140 ;
        RECT 2614.020 9.130 2617.020 9.140 ;
        RECT 2704.020 9.130 2707.020 9.140 ;
        RECT 2794.020 9.130 2797.020 9.140 ;
        RECT 2884.020 9.130 2887.020 9.140 ;
        RECT 2926.600 9.130 2929.600 9.140 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 94.020 -1.620 97.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 274.020 -1.620 277.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 454.020 -1.620 457.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 634.020 -1.620 637.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 814.020 -1.620 817.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 994.020 -1.620 997.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1174.020 -1.620 1177.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1354.020 -1.620 1357.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1534.020 -1.620 1537.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1714.020 -1.620 1717.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1894.020 -1.620 1897.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2074.020 -1.620 2077.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2254.020 -1.620 2257.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2434.020 -1.620 2437.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2614.020 -1.620 2617.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2794.020 -1.620 2797.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 94.020 -4.630 97.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 274.020 -4.630 277.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 454.020 -4.630 457.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 634.020 -4.630 637.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 814.020 -4.630 817.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 994.020 -4.630 997.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1174.020 -4.630 1177.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1354.020 -4.630 1357.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1534.020 -4.630 1537.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1714.020 -4.630 1717.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1894.020 -4.630 1897.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2074.020 -4.630 2077.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2254.020 -4.630 2257.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2434.020 -4.630 2437.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2614.020 -4.630 2617.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2794.020 -4.630 2797.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    ANTENNAGATEAREA 1320.207520 ;
    ANTENNADIFFAREA 842.456604 ;
    PORT
      LAYER pwell ;
        RECT 19.925 3506.400 20.095 3506.925 ;
        RECT 34.185 3506.400 34.355 3506.925 ;
        RECT 48.445 3506.400 48.615 3506.925 ;
        RECT 62.705 3506.400 62.875 3506.925 ;
        RECT 76.965 3506.400 77.135 3506.925 ;
        RECT 91.225 3506.400 91.395 3506.925 ;
        RECT 105.485 3506.400 105.655 3506.925 ;
        RECT 119.745 3506.400 119.915 3506.925 ;
        RECT 134.005 3506.400 134.175 3506.925 ;
        RECT 148.265 3506.400 148.435 3506.925 ;
        RECT 162.525 3506.400 162.695 3506.925 ;
        RECT 176.785 3506.400 176.955 3506.925 ;
        RECT 191.045 3506.400 191.215 3506.925 ;
        RECT 205.305 3506.400 205.475 3506.925 ;
        RECT 219.565 3506.400 219.735 3506.925 ;
        RECT 233.825 3506.400 233.995 3506.925 ;
        RECT 248.085 3506.400 248.255 3506.925 ;
        RECT 262.345 3506.400 262.515 3506.925 ;
        RECT 276.605 3506.400 276.775 3506.925 ;
        RECT 290.865 3506.400 291.035 3506.925 ;
        RECT 305.125 3506.400 305.295 3506.925 ;
        RECT 319.385 3506.400 319.555 3506.925 ;
        RECT 333.645 3506.400 333.815 3506.925 ;
        RECT 347.905 3506.400 348.075 3506.925 ;
        RECT 362.165 3506.400 362.335 3506.925 ;
        RECT 376.425 3506.400 376.595 3506.925 ;
        RECT 390.685 3506.400 390.855 3506.925 ;
        RECT 404.945 3506.400 405.115 3506.925 ;
        RECT 419.205 3506.400 419.375 3506.925 ;
        RECT 433.465 3506.400 433.635 3506.925 ;
        RECT 447.725 3506.400 447.895 3506.925 ;
        RECT 461.985 3506.400 462.155 3506.925 ;
        RECT 476.245 3506.400 476.415 3506.925 ;
        RECT 490.505 3506.400 490.675 3506.925 ;
        RECT 504.765 3506.400 504.935 3506.925 ;
        RECT 519.025 3506.400 519.195 3506.925 ;
        RECT 533.285 3506.400 533.455 3506.925 ;
        RECT 547.545 3506.400 547.715 3506.925 ;
        RECT 561.805 3506.400 561.975 3506.925 ;
        RECT 576.065 3506.400 576.235 3506.925 ;
        RECT 590.325 3506.400 590.495 3506.925 ;
        RECT 604.585 3506.400 604.755 3506.925 ;
        RECT 618.845 3506.400 619.015 3506.925 ;
        RECT 633.105 3506.400 633.275 3506.925 ;
        RECT 647.365 3506.400 647.535 3506.925 ;
        RECT 661.625 3506.400 661.795 3506.925 ;
        RECT 675.885 3506.400 676.055 3506.925 ;
        RECT 690.145 3506.400 690.315 3506.925 ;
        RECT 704.405 3506.400 704.575 3506.925 ;
        RECT 718.665 3506.400 718.835 3506.925 ;
        RECT 732.925 3506.400 733.095 3506.925 ;
        RECT 747.185 3506.400 747.355 3506.925 ;
        RECT 761.445 3506.400 761.615 3506.925 ;
        RECT 775.705 3506.400 775.875 3506.925 ;
        RECT 789.965 3506.400 790.135 3506.925 ;
        RECT 804.225 3506.400 804.395 3506.925 ;
        RECT 818.485 3506.400 818.655 3506.925 ;
        RECT 832.745 3506.400 832.915 3506.925 ;
        RECT 847.005 3506.400 847.175 3506.925 ;
        RECT 861.265 3506.400 861.435 3506.925 ;
        RECT 875.525 3506.400 875.695 3506.925 ;
        RECT 889.785 3506.400 889.955 3506.925 ;
        RECT 904.045 3506.400 904.215 3506.925 ;
        RECT 918.305 3506.400 918.475 3506.925 ;
        RECT 932.565 3506.400 932.735 3506.925 ;
        RECT 946.825 3506.400 946.995 3506.925 ;
        RECT 961.085 3506.400 961.255 3506.925 ;
        RECT 975.345 3506.400 975.515 3506.925 ;
        RECT 989.605 3506.400 989.775 3506.925 ;
        RECT 1003.865 3506.400 1004.035 3506.925 ;
        RECT 1018.125 3506.400 1018.295 3506.925 ;
        RECT 1032.385 3506.400 1032.555 3506.925 ;
        RECT 1046.645 3506.400 1046.815 3506.925 ;
        RECT 1060.905 3506.400 1061.075 3506.925 ;
        RECT 1075.165 3506.400 1075.335 3506.925 ;
        RECT 1089.425 3506.400 1089.595 3506.925 ;
        RECT 1103.685 3506.400 1103.855 3506.925 ;
        RECT 1117.945 3506.400 1118.115 3506.925 ;
        RECT 1132.205 3506.400 1132.375 3506.925 ;
        RECT 1146.465 3506.400 1146.635 3506.925 ;
        RECT 1160.725 3506.400 1160.895 3506.925 ;
        RECT 1174.985 3506.400 1175.155 3506.925 ;
        RECT 1189.245 3506.400 1189.415 3506.925 ;
        RECT 1203.505 3506.400 1203.675 3506.925 ;
        RECT 1217.765 3506.400 1217.935 3506.925 ;
        RECT 1232.025 3506.400 1232.195 3506.925 ;
        RECT 1246.285 3506.400 1246.455 3506.925 ;
        RECT 1260.545 3506.400 1260.715 3506.925 ;
        RECT 1274.805 3506.400 1274.975 3506.925 ;
        RECT 1289.065 3506.400 1289.235 3506.925 ;
        RECT 1303.325 3506.400 1303.495 3506.925 ;
        RECT 1317.585 3506.400 1317.755 3506.925 ;
        RECT 1331.845 3506.400 1332.015 3506.925 ;
        RECT 1346.105 3506.400 1346.275 3506.925 ;
        RECT 1360.365 3506.400 1360.535 3506.925 ;
        RECT 1374.625 3506.400 1374.795 3506.925 ;
        RECT 1388.885 3506.400 1389.055 3506.925 ;
        RECT 1403.145 3506.400 1403.315 3506.925 ;
        RECT 1417.405 3506.400 1417.575 3506.925 ;
        RECT 1431.665 3506.400 1431.835 3506.925 ;
        RECT 1445.925 3506.400 1446.095 3506.925 ;
        RECT 1460.185 3506.400 1460.355 3506.925 ;
        RECT 1474.445 3506.400 1474.615 3506.925 ;
        RECT 1488.705 3506.400 1488.875 3506.925 ;
        RECT 1502.965 3506.400 1503.135 3506.925 ;
        RECT 1517.225 3506.400 1517.395 3506.925 ;
        RECT 1531.485 3506.400 1531.655 3506.925 ;
        RECT 1545.745 3506.400 1545.915 3506.925 ;
        RECT 1560.005 3506.400 1560.175 3506.925 ;
        RECT 1574.265 3506.400 1574.435 3506.925 ;
        RECT 1588.525 3506.400 1588.695 3506.925 ;
        RECT 1602.785 3506.400 1602.955 3506.925 ;
        RECT 1617.045 3506.400 1617.215 3506.925 ;
        RECT 1631.305 3506.400 1631.475 3506.925 ;
        RECT 1645.565 3506.400 1645.735 3506.925 ;
        RECT 1659.825 3506.400 1659.995 3506.925 ;
        RECT 1674.085 3506.400 1674.255 3506.925 ;
        RECT 1688.345 3506.400 1688.515 3506.925 ;
        RECT 1702.605 3506.400 1702.775 3506.925 ;
        RECT 1716.865 3506.400 1717.035 3506.925 ;
        RECT 1731.125 3506.400 1731.295 3506.925 ;
        RECT 1745.385 3506.400 1745.555 3506.925 ;
        RECT 1759.645 3506.400 1759.815 3506.925 ;
        RECT 1773.905 3506.400 1774.075 3506.925 ;
        RECT 1788.165 3506.400 1788.335 3506.925 ;
        RECT 1802.425 3506.400 1802.595 3506.925 ;
        RECT 1816.685 3506.400 1816.855 3506.925 ;
        RECT 1830.945 3506.400 1831.115 3506.925 ;
        RECT 1845.205 3506.400 1845.375 3506.925 ;
        RECT 1859.465 3506.400 1859.635 3506.925 ;
        RECT 1873.725 3506.400 1873.895 3506.925 ;
        RECT 1887.985 3506.400 1888.155 3506.925 ;
        RECT 1902.245 3506.400 1902.415 3506.925 ;
        RECT 1916.505 3506.400 1916.675 3506.925 ;
        RECT 1930.765 3506.400 1930.935 3506.925 ;
        RECT 1945.025 3506.400 1945.195 3506.925 ;
        RECT 1959.285 3506.400 1959.455 3506.925 ;
        RECT 1973.545 3506.400 1973.715 3506.925 ;
        RECT 1987.805 3506.400 1987.975 3506.925 ;
        RECT 2002.065 3506.400 2002.235 3506.925 ;
        RECT 2016.325 3506.400 2016.495 3506.925 ;
        RECT 2030.585 3506.400 2030.755 3506.925 ;
        RECT 2044.845 3506.400 2045.015 3506.925 ;
        RECT 2059.105 3506.400 2059.275 3506.925 ;
        RECT 2073.365 3506.400 2073.535 3506.925 ;
        RECT 2087.625 3506.400 2087.795 3506.925 ;
        RECT 2101.885 3506.400 2102.055 3506.925 ;
        RECT 2116.145 3506.400 2116.315 3506.925 ;
        RECT 2130.405 3506.400 2130.575 3506.925 ;
        RECT 2144.665 3506.400 2144.835 3506.925 ;
        RECT 2158.925 3506.400 2159.095 3506.925 ;
        RECT 2173.185 3506.400 2173.355 3506.925 ;
        RECT 2187.445 3506.400 2187.615 3506.925 ;
        RECT 2201.705 3506.400 2201.875 3506.925 ;
        RECT 2215.965 3506.400 2216.135 3506.925 ;
        RECT 2230.225 3506.400 2230.395 3506.925 ;
        RECT 2244.485 3506.400 2244.655 3506.925 ;
        RECT 2258.745 3506.400 2258.915 3506.925 ;
        RECT 2273.005 3506.400 2273.175 3506.925 ;
        RECT 2287.265 3506.400 2287.435 3506.925 ;
        RECT 2301.525 3506.400 2301.695 3506.925 ;
        RECT 2315.785 3506.400 2315.955 3506.925 ;
        RECT 2330.045 3506.400 2330.215 3506.925 ;
        RECT 2344.305 3506.400 2344.475 3506.925 ;
        RECT 2358.565 3506.400 2358.735 3506.925 ;
        RECT 2372.825 3506.400 2372.995 3506.925 ;
        RECT 2387.085 3506.400 2387.255 3506.925 ;
        RECT 2401.345 3506.400 2401.515 3506.925 ;
        RECT 2415.605 3506.400 2415.775 3506.925 ;
        RECT 2429.865 3506.400 2430.035 3506.925 ;
        RECT 2444.125 3506.400 2444.295 3506.925 ;
        RECT 2458.385 3506.400 2458.555 3506.925 ;
        RECT 2472.645 3506.400 2472.815 3506.925 ;
        RECT 2486.905 3506.400 2487.075 3506.925 ;
        RECT 2501.165 3506.400 2501.335 3506.925 ;
        RECT 2515.425 3506.400 2515.595 3506.925 ;
        RECT 2529.685 3506.400 2529.855 3506.925 ;
        RECT 2543.945 3506.400 2544.115 3506.925 ;
        RECT 2558.205 3506.400 2558.375 3506.925 ;
        RECT 2572.465 3506.400 2572.635 3506.925 ;
        RECT 2586.725 3506.400 2586.895 3506.925 ;
        RECT 2600.985 3506.400 2601.155 3506.925 ;
        RECT 2615.245 3506.400 2615.415 3506.925 ;
        RECT 2629.505 3506.400 2629.675 3506.925 ;
        RECT 2643.765 3506.400 2643.935 3506.925 ;
        RECT 2658.025 3506.400 2658.195 3506.925 ;
        RECT 2672.285 3506.400 2672.455 3506.925 ;
        RECT 2686.545 3506.400 2686.715 3506.925 ;
        RECT 2700.805 3506.400 2700.975 3506.925 ;
        RECT 2715.065 3506.400 2715.235 3506.925 ;
        RECT 2729.325 3506.400 2729.495 3506.925 ;
        RECT 2743.585 3506.400 2743.755 3506.925 ;
        RECT 2757.845 3506.400 2758.015 3506.925 ;
        RECT 2772.105 3506.400 2772.275 3506.925 ;
        RECT 2786.365 3506.400 2786.535 3506.925 ;
        RECT 2800.625 3506.400 2800.795 3506.925 ;
        RECT 2814.885 3506.400 2815.055 3506.925 ;
        RECT 2829.145 3506.400 2829.315 3506.925 ;
        RECT 2843.405 3506.400 2843.575 3506.925 ;
        RECT 2857.665 3506.400 2857.835 3506.925 ;
        RECT 2871.925 3506.400 2872.095 3506.925 ;
        RECT 2886.185 3506.400 2886.355 3506.925 ;
        RECT 2900.445 3506.400 2900.615 3506.925 ;
        RECT 2910.105 3500.960 2910.275 3501.485 ;
        RECT 2910.105 3495.520 2910.275 3496.045 ;
        RECT 2910.105 3490.080 2910.275 3490.605 ;
        RECT 2910.105 3484.640 2910.275 3485.165 ;
        RECT 2910.105 3479.200 2910.275 3479.725 ;
        RECT 2910.105 3473.760 2910.275 3474.285 ;
        RECT 2910.105 3468.320 2910.275 3468.845 ;
        RECT 2910.105 3462.880 2910.275 3463.405 ;
        RECT 2910.105 3457.440 2910.275 3457.965 ;
        RECT 2910.105 3452.000 2910.275 3452.525 ;
        RECT 2910.105 3446.560 2910.275 3447.085 ;
        RECT 2910.105 3441.120 2910.275 3441.645 ;
        RECT 2910.105 3435.680 2910.275 3436.205 ;
        RECT 2910.105 3430.240 2910.275 3430.765 ;
        RECT 2910.105 3424.800 2910.275 3425.325 ;
        RECT 2910.105 3419.360 2910.275 3419.885 ;
        RECT 2910.105 3413.920 2910.275 3414.445 ;
        RECT 2910.105 3408.480 2910.275 3409.005 ;
        RECT 2910.105 3403.040 2910.275 3403.565 ;
        RECT 2910.105 3397.600 2910.275 3398.125 ;
        RECT 2910.105 3392.160 2910.275 3392.685 ;
        RECT 2910.105 3386.720 2910.275 3387.245 ;
        RECT 2910.105 3381.280 2910.275 3381.805 ;
        RECT 2910.105 3375.840 2910.275 3376.365 ;
        RECT 2910.105 3370.400 2910.275 3370.925 ;
        RECT 2910.105 3364.960 2910.275 3365.485 ;
        RECT 2910.105 3359.520 2910.275 3360.045 ;
        RECT 2910.105 3354.080 2910.275 3354.605 ;
        RECT 2910.105 3348.640 2910.275 3349.165 ;
        RECT 2910.105 3343.200 2910.275 3343.725 ;
        RECT 2910.105 3337.760 2910.275 3338.285 ;
        RECT 2910.105 3332.320 2910.275 3332.845 ;
        RECT 2910.105 3326.880 2910.275 3327.405 ;
        RECT 2910.105 3321.440 2910.275 3321.965 ;
        RECT 2910.105 3316.000 2910.275 3316.525 ;
        RECT 2910.105 3310.560 2910.275 3311.085 ;
        RECT 2910.105 3305.120 2910.275 3305.645 ;
        RECT 2910.105 3299.680 2910.275 3300.205 ;
        RECT 2910.105 3294.240 2910.275 3294.765 ;
        RECT 2910.105 3288.800 2910.275 3289.325 ;
        RECT 2910.105 3283.360 2910.275 3283.885 ;
        RECT 2910.105 3277.920 2910.275 3278.445 ;
        RECT 2910.105 3272.480 2910.275 3273.005 ;
        RECT 2910.105 3267.040 2910.275 3267.565 ;
        RECT 2910.105 3261.600 2910.275 3262.125 ;
        RECT 2910.105 3256.160 2910.275 3256.685 ;
        RECT 2910.105 3250.720 2910.275 3251.245 ;
        RECT 2910.105 3245.280 2910.275 3245.805 ;
        RECT 2910.105 3239.840 2910.275 3240.365 ;
        RECT 2910.105 3234.400 2910.275 3234.925 ;
        RECT 2910.105 3228.960 2910.275 3229.485 ;
        RECT 2910.105 3223.520 2910.275 3224.045 ;
        RECT 2910.105 3218.080 2910.275 3218.605 ;
        RECT 2910.105 3212.640 2910.275 3213.165 ;
        RECT 2910.105 3207.200 2910.275 3207.725 ;
        RECT 2910.105 3201.760 2910.275 3202.285 ;
        RECT 2910.105 3196.320 2910.275 3196.845 ;
        RECT 2910.105 3190.880 2910.275 3191.405 ;
        RECT 2910.105 3185.440 2910.275 3185.965 ;
        RECT 2910.105 3180.000 2910.275 3180.525 ;
        RECT 2910.105 3174.560 2910.275 3175.085 ;
        RECT 2910.105 3169.120 2910.275 3169.645 ;
        RECT 2910.105 3163.680 2910.275 3164.205 ;
        RECT 2910.105 3158.240 2910.275 3158.765 ;
        RECT 2910.105 3152.800 2910.275 3153.325 ;
        RECT 2910.105 3147.360 2910.275 3147.885 ;
        RECT 2910.105 3141.920 2910.275 3142.445 ;
        RECT 2910.105 3136.480 2910.275 3137.005 ;
        RECT 2910.105 3131.040 2910.275 3131.565 ;
        RECT 2910.105 3125.600 2910.275 3126.125 ;
        RECT 2910.105 3120.160 2910.275 3120.685 ;
        RECT 2910.105 3114.720 2910.275 3115.245 ;
        RECT 2910.105 3109.280 2910.275 3109.805 ;
        RECT 2910.105 3103.840 2910.275 3104.365 ;
        RECT 2910.105 3098.400 2910.275 3098.925 ;
        RECT 2910.105 3092.960 2910.275 3093.485 ;
        RECT 2910.105 3087.520 2910.275 3088.045 ;
        RECT 2910.105 3082.080 2910.275 3082.605 ;
        RECT 2910.105 3076.640 2910.275 3077.165 ;
        RECT 2910.105 3071.200 2910.275 3071.725 ;
        RECT 2910.105 3065.760 2910.275 3066.285 ;
        RECT 2910.105 3060.320 2910.275 3060.845 ;
        RECT 2910.105 3054.880 2910.275 3055.405 ;
        RECT 2910.105 3049.440 2910.275 3049.965 ;
        RECT 2910.105 3044.000 2910.275 3044.525 ;
        RECT 2910.105 3038.560 2910.275 3039.085 ;
        RECT 2910.105 3033.120 2910.275 3033.645 ;
        RECT 2910.105 3027.680 2910.275 3028.205 ;
        RECT 2910.105 3022.240 2910.275 3022.765 ;
        RECT 2910.105 3016.800 2910.275 3017.325 ;
        RECT 2910.105 3011.360 2910.275 3011.885 ;
        RECT 2910.105 3005.920 2910.275 3006.445 ;
        RECT 2910.105 3000.480 2910.275 3001.005 ;
        RECT 2910.105 2995.040 2910.275 2995.565 ;
        RECT 2910.105 2989.600 2910.275 2990.125 ;
        RECT 2910.105 2984.160 2910.275 2984.685 ;
        RECT 2910.105 2978.720 2910.275 2979.245 ;
        RECT 2910.105 2973.280 2910.275 2973.805 ;
        RECT 2910.105 2967.840 2910.275 2968.365 ;
        RECT 2910.105 2962.400 2910.275 2962.925 ;
        RECT 2910.105 2956.960 2910.275 2957.485 ;
        RECT 2910.105 2951.520 2910.275 2952.045 ;
        RECT 2910.105 2946.080 2910.275 2946.605 ;
        RECT 2910.105 2940.640 2910.275 2941.165 ;
        RECT 2910.105 2935.200 2910.275 2935.725 ;
        RECT 2910.105 2929.760 2910.275 2930.285 ;
        RECT 2910.105 2924.320 2910.275 2924.845 ;
        RECT 2910.105 2918.880 2910.275 2919.405 ;
        RECT 2910.105 2913.440 2910.275 2913.965 ;
        RECT 2910.105 2908.000 2910.275 2908.525 ;
        RECT 2910.105 2902.560 2910.275 2903.085 ;
        RECT 2910.105 2897.120 2910.275 2897.645 ;
        RECT 2910.105 2891.680 2910.275 2892.205 ;
        RECT 2910.105 2886.240 2910.275 2886.765 ;
        RECT 2910.105 2880.800 2910.275 2881.325 ;
        RECT 2910.105 2875.360 2910.275 2875.885 ;
        RECT 2910.105 2869.920 2910.275 2870.445 ;
        RECT 2910.105 2864.480 2910.275 2865.005 ;
        RECT 2910.105 2859.040 2910.275 2859.565 ;
        RECT 2910.105 2853.600 2910.275 2854.125 ;
        RECT 2910.105 2848.160 2910.275 2848.685 ;
        RECT 2910.105 2842.720 2910.275 2843.245 ;
        RECT 2910.105 2837.280 2910.275 2837.805 ;
        RECT 2910.105 2831.840 2910.275 2832.365 ;
        RECT 2910.105 2826.400 2910.275 2826.925 ;
        RECT 2910.105 2820.960 2910.275 2821.485 ;
        RECT 2910.105 2815.520 2910.275 2816.045 ;
        RECT 2910.105 2810.080 2910.275 2810.605 ;
        RECT 2910.105 2804.640 2910.275 2805.165 ;
        RECT 2910.105 2799.200 2910.275 2799.725 ;
        RECT 2910.105 2793.760 2910.275 2794.285 ;
        RECT 2910.105 2788.320 2910.275 2788.845 ;
        RECT 2910.105 2782.880 2910.275 2783.405 ;
        RECT 2910.105 2777.440 2910.275 2777.965 ;
        RECT 2910.105 2772.000 2910.275 2772.525 ;
        RECT 2910.105 2766.560 2910.275 2767.085 ;
        RECT 2910.105 2761.120 2910.275 2761.645 ;
        RECT 2910.105 2755.680 2910.275 2756.205 ;
        RECT 2910.105 2750.240 2910.275 2750.765 ;
        RECT 2910.105 2744.800 2910.275 2745.325 ;
        RECT 2910.105 2739.360 2910.275 2739.885 ;
        RECT 2910.105 2733.920 2910.275 2734.445 ;
        RECT 2910.105 2728.480 2910.275 2729.005 ;
        RECT 2910.105 2723.040 2910.275 2723.565 ;
        RECT 2910.105 2717.600 2910.275 2718.125 ;
        RECT 2910.105 2712.160 2910.275 2712.685 ;
        RECT 2910.105 2706.720 2910.275 2707.245 ;
        RECT 2910.105 2701.280 2910.275 2701.805 ;
        RECT 2910.105 2695.840 2910.275 2696.365 ;
        RECT 2906.425 2689.235 2906.595 2689.760 ;
        RECT 2906.425 2683.795 2906.595 2684.320 ;
        RECT 2906.425 2678.355 2906.595 2678.880 ;
        RECT 2906.425 2672.915 2906.595 2673.440 ;
        RECT 2906.425 2667.475 2906.595 2668.000 ;
        RECT 2906.425 2662.035 2906.595 2662.560 ;
        RECT 2906.425 2656.595 2906.595 2657.120 ;
        RECT 2906.425 2651.155 2906.595 2651.680 ;
        RECT 2906.425 2645.715 2906.595 2646.240 ;
        RECT 2906.425 2640.275 2906.595 2640.800 ;
        RECT 2906.425 2634.835 2906.595 2635.360 ;
        RECT 2906.425 2629.395 2906.595 2629.920 ;
        RECT 2906.425 2623.955 2906.595 2624.480 ;
        RECT 2906.425 2618.515 2906.595 2619.040 ;
        RECT 2906.425 2613.075 2906.595 2613.600 ;
        RECT 2906.425 2607.635 2906.595 2608.160 ;
        RECT 2906.425 2602.195 2906.595 2602.720 ;
        RECT 2906.425 2596.755 2906.595 2597.280 ;
        RECT 2906.425 2591.315 2906.595 2591.840 ;
        RECT 2906.425 2585.875 2906.595 2586.400 ;
        RECT 2906.425 2580.435 2906.595 2580.960 ;
        RECT 2906.425 2574.995 2906.595 2575.520 ;
        RECT 2906.425 2569.555 2906.595 2570.080 ;
        RECT 2906.425 2564.115 2906.595 2564.640 ;
        RECT 2906.425 2558.675 2906.595 2559.200 ;
        RECT 2906.425 2553.235 2906.595 2553.760 ;
        RECT 2906.425 2547.795 2906.595 2548.320 ;
        RECT 2906.425 2542.355 2906.595 2542.880 ;
        RECT 2906.425 2536.915 2906.595 2537.440 ;
        RECT 2906.425 2531.475 2906.595 2532.000 ;
        RECT 2906.425 2526.035 2906.595 2526.560 ;
        RECT 2906.425 2520.595 2906.595 2521.120 ;
        RECT 2906.425 2515.155 2906.595 2515.680 ;
        RECT 2906.425 2509.715 2906.595 2510.240 ;
        RECT 2906.425 2504.275 2906.595 2504.800 ;
        RECT 2906.425 2498.835 2906.595 2499.360 ;
        RECT 2906.425 2493.395 2906.595 2493.920 ;
        RECT 2906.425 2487.955 2906.595 2488.480 ;
        RECT 2906.425 2482.515 2906.595 2483.040 ;
        RECT 2906.425 2477.075 2906.595 2477.600 ;
        RECT 2906.425 2471.635 2906.595 2472.160 ;
        RECT 2906.425 2466.195 2906.595 2466.720 ;
        RECT 2906.425 2460.755 2906.595 2461.280 ;
        RECT 2906.425 2455.315 2906.595 2455.840 ;
        RECT 2906.425 2449.875 2906.595 2450.400 ;
        RECT 2906.425 2444.435 2906.595 2444.960 ;
        RECT 2906.425 2438.995 2906.595 2439.520 ;
        RECT 2906.425 2433.555 2906.595 2434.080 ;
        RECT 2906.425 2428.115 2906.595 2428.640 ;
        RECT 2906.425 2422.675 2906.595 2423.200 ;
        RECT 2906.425 2417.235 2906.595 2417.760 ;
        RECT 2906.425 2411.795 2906.595 2412.320 ;
        RECT 2906.425 2406.355 2906.595 2406.880 ;
        RECT 2906.425 2400.915 2906.595 2401.440 ;
        RECT 2906.425 2395.475 2906.595 2396.000 ;
        RECT 2906.425 2390.035 2906.595 2390.560 ;
        RECT 2906.425 2384.595 2906.595 2385.120 ;
        RECT 2906.425 2379.155 2906.595 2379.680 ;
        RECT 2906.425 2373.715 2906.595 2374.240 ;
        RECT 2906.425 2368.275 2906.595 2368.800 ;
        RECT 2906.425 2362.835 2906.595 2363.360 ;
        RECT 2906.425 2357.395 2906.595 2357.920 ;
        RECT 2906.425 2351.955 2906.595 2352.480 ;
        RECT 2906.425 2346.515 2906.595 2347.040 ;
        RECT 2906.425 2341.075 2906.595 2341.600 ;
        RECT 2906.425 2335.635 2906.595 2336.160 ;
        RECT 2906.425 2330.195 2906.595 2330.720 ;
        RECT 2906.425 2324.755 2906.595 2325.280 ;
        RECT 2906.425 2319.315 2906.595 2319.840 ;
        RECT 2906.425 2313.875 2906.595 2314.400 ;
        RECT 2906.425 2308.435 2906.595 2308.960 ;
        RECT 2906.425 2302.995 2906.595 2303.520 ;
        RECT 2906.425 2297.555 2906.595 2298.080 ;
        RECT 2906.425 2292.115 2906.595 2292.640 ;
        RECT 2906.425 2286.675 2906.595 2287.200 ;
        RECT 2906.425 2281.235 2906.595 2281.760 ;
        RECT 2906.425 2275.795 2906.595 2276.320 ;
        RECT 2906.425 2270.355 2906.595 2270.880 ;
        RECT 2906.425 2264.915 2906.595 2265.440 ;
        RECT 2906.425 2259.475 2906.595 2260.000 ;
        RECT 2906.425 2254.035 2906.595 2254.560 ;
        RECT 2906.425 2248.595 2906.595 2249.120 ;
        RECT 2906.425 2243.155 2906.595 2243.680 ;
        RECT 2906.425 2237.715 2906.595 2238.240 ;
        RECT 2906.425 2232.275 2906.595 2232.800 ;
        RECT 2906.425 2226.835 2906.595 2227.360 ;
        RECT 2906.425 2221.395 2906.595 2221.920 ;
        RECT 2906.425 2215.955 2906.595 2216.480 ;
        RECT 2906.425 2210.515 2906.595 2211.040 ;
        RECT 2906.425 2205.075 2906.595 2205.600 ;
        RECT 2906.425 2199.635 2906.595 2200.160 ;
        RECT 2906.425 2194.195 2906.595 2194.720 ;
        RECT 2906.425 2188.755 2906.595 2189.280 ;
        RECT 2906.425 2183.315 2906.595 2183.840 ;
        RECT 2906.425 2177.875 2906.595 2178.400 ;
        RECT 2906.425 2172.435 2906.595 2172.960 ;
        RECT 2906.425 2166.995 2906.595 2167.520 ;
        RECT 2906.425 2161.555 2906.595 2162.080 ;
        RECT 2906.425 2156.115 2906.595 2156.640 ;
        RECT 2906.425 2150.675 2906.595 2151.200 ;
        RECT 2906.425 2145.235 2906.595 2145.760 ;
        RECT 2906.425 2139.795 2906.595 2140.320 ;
        RECT 2906.425 2134.355 2906.595 2134.880 ;
        RECT 2906.425 2128.915 2906.595 2129.440 ;
        RECT 2906.425 2123.475 2906.595 2124.000 ;
        RECT 2906.425 2118.035 2906.595 2118.560 ;
        RECT 2906.425 2112.595 2906.595 2113.120 ;
        RECT 2906.425 2107.155 2906.595 2107.680 ;
        RECT 2906.425 2101.715 2906.595 2102.240 ;
        RECT 2906.425 2096.275 2906.595 2096.800 ;
        RECT 2906.425 2090.835 2906.595 2091.360 ;
        RECT 2906.425 2085.395 2906.595 2085.920 ;
        RECT 2906.425 2079.955 2906.595 2080.480 ;
        RECT 2906.425 2074.515 2906.595 2075.040 ;
        RECT 2906.425 2069.075 2906.595 2069.600 ;
        RECT 2906.425 2063.635 2906.595 2064.160 ;
        RECT 2906.425 2058.195 2906.595 2058.720 ;
        RECT 2906.425 2052.755 2906.595 2053.280 ;
        RECT 2906.425 2047.315 2906.595 2047.840 ;
        RECT 2906.425 2041.875 2906.595 2042.400 ;
        RECT 2906.425 2036.435 2906.595 2036.960 ;
        RECT 2906.425 2030.995 2906.595 2031.520 ;
        RECT 2906.425 2025.555 2906.595 2026.080 ;
        RECT 2906.425 2020.115 2906.595 2020.640 ;
        RECT 2906.425 2014.675 2906.595 2015.200 ;
        RECT 2906.425 2009.235 2906.595 2009.760 ;
        RECT 2906.425 2003.795 2906.595 2004.320 ;
        RECT 2906.425 1998.355 2906.595 1998.880 ;
        RECT 2906.425 1992.915 2906.595 1993.440 ;
        RECT 2906.425 1987.475 2906.595 1988.000 ;
        RECT 2906.425 1982.035 2906.595 1982.560 ;
        RECT 2906.425 1976.595 2906.595 1977.120 ;
        RECT 2906.425 1971.155 2906.595 1971.680 ;
        RECT 2906.425 1965.715 2906.595 1966.240 ;
        RECT 2906.425 1960.275 2906.595 1960.800 ;
        RECT 2906.425 1954.835 2906.595 1955.360 ;
        RECT 2906.425 1949.395 2906.595 1949.920 ;
        RECT 2906.425 1943.955 2906.595 1944.480 ;
        RECT 2906.425 1938.515 2906.595 1939.040 ;
        RECT 2906.425 1933.075 2906.595 1933.600 ;
        RECT 2906.425 1927.635 2906.595 1928.160 ;
        RECT 2906.425 1922.195 2906.595 1922.720 ;
        RECT 2906.425 1916.755 2906.595 1917.280 ;
        RECT 2906.425 1911.315 2906.595 1911.840 ;
        RECT 2906.425 1905.875 2906.595 1906.400 ;
        RECT 2906.425 1900.435 2906.595 1900.960 ;
        RECT 2906.425 1894.995 2906.595 1895.520 ;
        RECT 2906.425 1889.555 2906.595 1890.080 ;
        RECT 2906.425 1884.115 2906.595 1884.640 ;
        RECT 2906.425 1878.675 2906.595 1879.200 ;
        RECT 2906.425 1873.235 2906.595 1873.760 ;
        RECT 2906.425 1867.795 2906.595 1868.320 ;
        RECT 2906.425 1862.355 2906.595 1862.880 ;
        RECT 2906.425 1856.915 2906.595 1857.440 ;
        RECT 2906.425 1851.475 2906.595 1852.000 ;
        RECT 2906.425 1846.035 2906.595 1846.560 ;
        RECT 2906.425 1840.595 2906.595 1841.120 ;
        RECT 2906.425 1835.155 2906.595 1835.680 ;
        RECT 2906.425 1829.715 2906.595 1830.240 ;
        RECT 2906.425 1824.275 2906.595 1824.800 ;
        RECT 2906.425 1818.835 2906.595 1819.360 ;
        RECT 2906.425 1813.395 2906.595 1813.920 ;
        RECT 2906.425 1807.955 2906.595 1808.480 ;
        RECT 2906.425 1802.515 2906.595 1803.040 ;
        RECT 2906.425 1797.075 2906.595 1797.600 ;
        RECT 2906.425 1791.635 2906.595 1792.160 ;
        RECT 2906.425 1786.195 2906.595 1786.720 ;
        RECT 2906.425 1780.755 2906.595 1781.280 ;
        RECT 2906.425 1775.315 2906.595 1775.840 ;
        RECT 2906.425 1769.875 2906.595 1770.400 ;
        RECT 2906.425 1764.435 2906.595 1764.960 ;
        RECT 2906.425 1758.995 2906.595 1759.520 ;
        RECT 2906.425 1753.555 2906.595 1754.080 ;
        RECT 2906.425 1748.115 2906.595 1748.640 ;
        RECT 2906.425 1742.675 2906.595 1743.200 ;
        RECT 2906.425 1737.235 2906.595 1737.760 ;
        RECT 2906.425 1731.795 2906.595 1732.320 ;
        RECT 2906.425 1726.355 2906.595 1726.880 ;
        RECT 2906.425 1720.915 2906.595 1721.440 ;
        RECT 2906.425 1715.475 2906.595 1716.000 ;
        RECT 2906.425 1710.035 2906.595 1710.560 ;
        RECT 2906.425 1704.595 2906.595 1705.120 ;
        RECT 2906.425 1699.155 2906.595 1699.680 ;
        RECT 2906.425 1693.715 2906.595 1694.240 ;
        RECT 2906.425 1688.275 2906.595 1688.800 ;
        RECT 2906.425 1682.835 2906.595 1683.360 ;
        RECT 2906.425 1677.395 2906.595 1677.920 ;
        RECT 2906.425 1671.955 2906.595 1672.480 ;
        RECT 2906.425 1666.515 2906.595 1667.040 ;
        RECT 2906.425 1661.075 2906.595 1661.600 ;
        RECT 2906.425 1655.635 2906.595 1656.160 ;
        RECT 2906.425 1650.195 2906.595 1650.720 ;
        RECT 2906.425 1644.755 2906.595 1645.280 ;
        RECT 2906.425 1639.315 2906.595 1639.840 ;
        RECT 2906.425 1633.875 2906.595 1634.400 ;
        RECT 2906.425 1628.435 2906.595 1628.960 ;
        RECT 2906.425 1622.995 2906.595 1623.520 ;
        RECT 2906.425 1617.555 2906.595 1618.080 ;
        RECT 2906.425 1612.115 2906.595 1612.640 ;
        RECT 2906.425 1606.675 2906.595 1607.200 ;
        RECT 2906.425 1601.235 2906.595 1601.760 ;
        RECT 2906.425 1595.795 2906.595 1596.320 ;
        RECT 2906.425 1590.355 2906.595 1590.880 ;
        RECT 2906.425 1584.915 2906.595 1585.440 ;
        RECT 2906.425 1579.475 2906.595 1580.000 ;
        RECT 2906.425 1574.035 2906.595 1574.560 ;
        RECT 2906.425 1568.595 2906.595 1569.120 ;
        RECT 2906.425 1563.155 2906.595 1563.680 ;
        RECT 2906.425 1557.715 2906.595 1558.240 ;
        RECT 2906.425 1552.275 2906.595 1552.800 ;
        RECT 2906.425 1546.835 2906.595 1547.360 ;
        RECT 2906.425 1541.395 2906.595 1541.920 ;
        RECT 2906.425 1535.955 2906.595 1536.480 ;
        RECT 2906.425 1530.515 2906.595 1531.040 ;
        RECT 2906.425 1525.075 2906.595 1525.600 ;
        RECT 2906.425 1519.635 2906.595 1520.160 ;
        RECT 2906.425 1514.195 2906.595 1514.720 ;
        RECT 2906.425 1508.755 2906.595 1509.280 ;
        RECT 2906.425 1503.315 2906.595 1503.840 ;
        RECT 2906.425 1497.875 2906.595 1498.400 ;
        RECT 2906.425 1492.435 2906.595 1492.960 ;
        RECT 2906.425 1486.995 2906.595 1487.520 ;
        RECT 2906.425 1481.555 2906.595 1482.080 ;
        RECT 2906.425 1476.115 2906.595 1476.640 ;
        RECT 2906.425 1470.675 2906.595 1471.200 ;
        RECT 2906.425 1465.235 2906.595 1465.760 ;
        RECT 2906.425 1459.795 2906.595 1460.320 ;
        RECT 2906.425 1454.355 2906.595 1454.880 ;
        RECT 2906.425 1448.915 2906.595 1449.440 ;
        RECT 2906.425 1443.475 2906.595 1444.000 ;
        RECT 2906.425 1438.035 2906.595 1438.560 ;
        RECT 2906.425 1432.595 2906.595 1433.120 ;
        RECT 2906.425 1427.155 2906.595 1427.680 ;
        RECT 2906.425 1421.715 2906.595 1422.240 ;
        RECT 2906.425 1416.275 2906.595 1416.800 ;
        RECT 2906.425 1410.835 2906.595 1411.360 ;
        RECT 2906.425 1405.395 2906.595 1405.920 ;
        RECT 2906.425 1399.955 2906.595 1400.480 ;
        RECT 2906.425 1394.515 2906.595 1395.040 ;
        RECT 2906.425 1389.075 2906.595 1389.600 ;
        RECT 2906.425 1383.635 2906.595 1384.160 ;
        RECT 2906.425 1378.195 2906.595 1378.720 ;
        RECT 2906.425 1372.755 2906.595 1373.280 ;
        RECT 2906.425 1367.315 2906.595 1367.840 ;
        RECT 2906.425 1361.875 2906.595 1362.400 ;
        RECT 2906.425 1356.435 2906.595 1356.960 ;
        RECT 2906.425 1350.995 2906.595 1351.520 ;
        RECT 2906.425 1345.555 2906.595 1346.080 ;
        RECT 2906.425 1340.115 2906.595 1340.640 ;
        RECT 2906.425 1334.675 2906.595 1335.200 ;
        RECT 2906.425 1329.235 2906.595 1329.760 ;
        RECT 2906.425 1323.795 2906.595 1324.320 ;
        RECT 2906.425 1318.355 2906.595 1318.880 ;
        RECT 2906.425 1312.915 2906.595 1313.440 ;
        RECT 2906.425 1307.475 2906.595 1308.000 ;
        RECT 2906.425 1302.035 2906.595 1302.560 ;
        RECT 2906.425 1296.595 2906.595 1297.120 ;
        RECT 2906.425 1291.155 2906.595 1291.680 ;
        RECT 2906.425 1285.715 2906.595 1286.240 ;
        RECT 2906.425 1280.275 2906.595 1280.800 ;
        RECT 2906.425 1274.835 2906.595 1275.360 ;
        RECT 2906.425 1269.395 2906.595 1269.920 ;
        RECT 2906.425 1263.955 2906.595 1264.480 ;
        RECT 2906.425 1258.515 2906.595 1259.040 ;
        RECT 2906.425 1253.075 2906.595 1253.600 ;
        RECT 2906.425 1247.635 2906.595 1248.160 ;
        RECT 2910.105 1237.920 2910.275 1238.445 ;
        RECT 2910.105 1232.480 2910.275 1233.005 ;
        RECT 2910.105 1227.040 2910.275 1227.565 ;
        RECT 2910.105 1221.600 2910.275 1222.125 ;
        RECT 2910.105 1216.160 2910.275 1216.685 ;
        RECT 2910.105 1210.720 2910.275 1211.245 ;
        RECT 2910.105 1205.280 2910.275 1205.805 ;
        RECT 2910.105 1199.840 2910.275 1200.365 ;
        RECT 2910.105 1194.400 2910.275 1194.925 ;
        RECT 2910.105 1188.960 2910.275 1189.485 ;
        RECT 2910.105 1183.520 2910.275 1184.045 ;
        RECT 2910.105 1178.080 2910.275 1178.605 ;
        RECT 2910.105 1172.640 2910.275 1173.165 ;
        RECT 2910.105 1167.200 2910.275 1167.725 ;
        RECT 2910.105 1161.760 2910.275 1162.285 ;
        RECT 2910.105 1156.320 2910.275 1156.845 ;
        RECT 2910.105 1150.880 2910.275 1151.405 ;
        RECT 2910.105 1145.440 2910.275 1145.965 ;
        RECT 2910.105 1140.000 2910.275 1140.525 ;
        RECT 2910.105 1134.560 2910.275 1135.085 ;
        RECT 2910.105 1129.120 2910.275 1129.645 ;
        RECT 2910.105 1123.680 2910.275 1124.205 ;
        RECT 2910.105 1118.240 2910.275 1118.765 ;
        RECT 2910.105 1112.800 2910.275 1113.325 ;
        RECT 2910.105 1107.360 2910.275 1107.885 ;
        RECT 2910.105 1101.920 2910.275 1102.445 ;
        RECT 2910.105 1096.480 2910.275 1097.005 ;
        RECT 2910.105 1091.040 2910.275 1091.565 ;
        RECT 2910.105 1085.600 2910.275 1086.125 ;
        RECT 2910.105 1080.160 2910.275 1080.685 ;
        RECT 2910.105 1074.720 2910.275 1075.245 ;
        RECT 2910.105 1069.280 2910.275 1069.805 ;
        RECT 2910.105 1063.840 2910.275 1064.365 ;
        RECT 2910.105 1058.400 2910.275 1058.925 ;
        RECT 2910.105 1052.960 2910.275 1053.485 ;
        RECT 2910.105 1047.520 2910.275 1048.045 ;
        RECT 2910.105 1042.080 2910.275 1042.605 ;
        RECT 2910.105 1036.640 2910.275 1037.165 ;
        RECT 2910.105 1031.200 2910.275 1031.725 ;
        RECT 2910.105 1025.760 2910.275 1026.285 ;
        RECT 2910.105 1020.320 2910.275 1020.845 ;
        RECT 2910.105 1014.880 2910.275 1015.405 ;
        RECT 2910.105 1009.440 2910.275 1009.965 ;
        RECT 2910.105 1004.000 2910.275 1004.525 ;
        RECT 2910.105 998.560 2910.275 999.085 ;
        RECT 2910.105 993.120 2910.275 993.645 ;
        RECT 2910.105 987.680 2910.275 988.205 ;
        RECT 2910.105 982.240 2910.275 982.765 ;
        RECT 2910.105 976.800 2910.275 977.325 ;
        RECT 2910.105 971.360 2910.275 971.885 ;
        RECT 2910.105 965.920 2910.275 966.445 ;
        RECT 2910.105 960.480 2910.275 961.005 ;
        RECT 2910.105 955.040 2910.275 955.565 ;
        RECT 2910.105 949.600 2910.275 950.125 ;
        RECT 2910.105 944.160 2910.275 944.685 ;
        RECT 2910.105 938.720 2910.275 939.245 ;
        RECT 2910.105 933.280 2910.275 933.805 ;
        RECT 2910.105 927.840 2910.275 928.365 ;
        RECT 2910.105 922.400 2910.275 922.925 ;
        RECT 2910.105 916.960 2910.275 917.485 ;
        RECT 2910.105 911.520 2910.275 912.045 ;
        RECT 2910.105 906.080 2910.275 906.605 ;
        RECT 2910.105 900.640 2910.275 901.165 ;
        RECT 2910.105 895.200 2910.275 895.725 ;
        RECT 2910.105 889.760 2910.275 890.285 ;
        RECT 2910.105 884.320 2910.275 884.845 ;
        RECT 2910.105 878.880 2910.275 879.405 ;
        RECT 2910.105 873.440 2910.275 873.965 ;
        RECT 2910.105 868.000 2910.275 868.525 ;
        RECT 2910.105 862.560 2910.275 863.085 ;
        RECT 2910.105 857.120 2910.275 857.645 ;
        RECT 2910.105 851.680 2910.275 852.205 ;
        RECT 2910.105 846.240 2910.275 846.765 ;
        RECT 2910.105 840.800 2910.275 841.325 ;
        RECT 2910.105 835.360 2910.275 835.885 ;
        RECT 2910.105 829.920 2910.275 830.445 ;
        RECT 2910.105 824.480 2910.275 825.005 ;
        RECT 2910.105 819.040 2910.275 819.565 ;
        RECT 2910.105 813.600 2910.275 814.125 ;
        RECT 2910.105 808.160 2910.275 808.685 ;
        RECT 2910.105 802.720 2910.275 803.245 ;
        RECT 2910.105 797.280 2910.275 797.805 ;
        RECT 2910.105 791.840 2910.275 792.365 ;
        RECT 2910.105 786.400 2910.275 786.925 ;
        RECT 2910.105 780.960 2910.275 781.485 ;
        RECT 2910.105 775.520 2910.275 776.045 ;
        RECT 2910.105 770.080 2910.275 770.605 ;
        RECT 2910.105 764.640 2910.275 765.165 ;
        RECT 2910.105 759.200 2910.275 759.725 ;
        RECT 2910.105 753.760 2910.275 754.285 ;
        RECT 2910.105 748.320 2910.275 748.845 ;
        RECT 2910.105 742.880 2910.275 743.405 ;
        RECT 2910.105 737.440 2910.275 737.965 ;
        RECT 2910.105 732.000 2910.275 732.525 ;
        RECT 2910.105 726.560 2910.275 727.085 ;
        RECT 2910.105 721.120 2910.275 721.645 ;
        RECT 2910.105 715.680 2910.275 716.205 ;
        RECT 2910.105 710.240 2910.275 710.765 ;
        RECT 2910.105 704.800 2910.275 705.325 ;
        RECT 2910.105 699.360 2910.275 699.885 ;
        RECT 2910.105 693.920 2910.275 694.445 ;
        RECT 2910.105 688.480 2910.275 689.005 ;
        RECT 2910.105 683.040 2910.275 683.565 ;
        RECT 2910.105 677.600 2910.275 678.125 ;
        RECT 2910.105 672.160 2910.275 672.685 ;
        RECT 2910.105 666.720 2910.275 667.245 ;
        RECT 2910.105 661.280 2910.275 661.805 ;
        RECT 2910.105 655.840 2910.275 656.365 ;
        RECT 2910.105 650.400 2910.275 650.925 ;
        RECT 2910.105 644.960 2910.275 645.485 ;
        RECT 2910.105 639.520 2910.275 640.045 ;
        RECT 2910.105 634.080 2910.275 634.605 ;
        RECT 2910.105 628.640 2910.275 629.165 ;
        RECT 2910.105 623.200 2910.275 623.725 ;
        RECT 2910.105 617.760 2910.275 618.285 ;
        RECT 2910.105 612.320 2910.275 612.845 ;
        RECT 2910.105 606.880 2910.275 607.405 ;
        RECT 2910.105 601.440 2910.275 601.965 ;
        RECT 2910.105 596.000 2910.275 596.525 ;
        RECT 2910.105 590.560 2910.275 591.085 ;
        RECT 2910.105 585.120 2910.275 585.645 ;
        RECT 2910.105 579.680 2910.275 580.205 ;
        RECT 2910.105 574.240 2910.275 574.765 ;
        RECT 2910.105 568.800 2910.275 569.325 ;
        RECT 2910.105 563.360 2910.275 563.885 ;
        RECT 2910.105 557.920 2910.275 558.445 ;
        RECT 2910.105 552.480 2910.275 553.005 ;
        RECT 2910.105 547.040 2910.275 547.565 ;
        RECT 2910.105 541.600 2910.275 542.125 ;
        RECT 2910.105 536.160 2910.275 536.685 ;
        RECT 2910.105 530.720 2910.275 531.245 ;
        RECT 2910.105 525.280 2910.275 525.805 ;
        RECT 2910.105 519.840 2910.275 520.365 ;
        RECT 2910.105 514.400 2910.275 514.925 ;
        RECT 2910.105 508.960 2910.275 509.485 ;
        RECT 2910.105 503.520 2910.275 504.045 ;
        RECT 2910.105 498.080 2910.275 498.605 ;
        RECT 2910.105 492.640 2910.275 493.165 ;
        RECT 2910.105 487.200 2910.275 487.725 ;
        RECT 2910.105 481.760 2910.275 482.285 ;
        RECT 2910.105 476.320 2910.275 476.845 ;
        RECT 2910.105 470.880 2910.275 471.405 ;
        RECT 2910.105 465.440 2910.275 465.965 ;
        RECT 2910.105 460.000 2910.275 460.525 ;
        RECT 2910.105 454.560 2910.275 455.085 ;
        RECT 2910.105 449.120 2910.275 449.645 ;
        RECT 2910.105 443.680 2910.275 444.205 ;
        RECT 2910.105 438.240 2910.275 438.765 ;
        RECT 2910.105 432.800 2910.275 433.325 ;
        RECT 2910.105 427.360 2910.275 427.885 ;
        RECT 2910.105 421.920 2910.275 422.445 ;
        RECT 2910.105 416.480 2910.275 417.005 ;
        RECT 2910.105 411.040 2910.275 411.565 ;
        RECT 2910.105 405.600 2910.275 406.125 ;
        RECT 2910.105 400.160 2910.275 400.685 ;
        RECT 2910.105 394.720 2910.275 395.245 ;
        RECT 2910.105 389.280 2910.275 389.805 ;
        RECT 2910.105 383.840 2910.275 384.365 ;
        RECT 2910.105 378.400 2910.275 378.925 ;
        RECT 2910.105 372.960 2910.275 373.485 ;
        RECT 2910.105 367.520 2910.275 368.045 ;
        RECT 2910.105 362.080 2910.275 362.605 ;
        RECT 2910.105 356.640 2910.275 357.165 ;
        RECT 2910.105 351.200 2910.275 351.725 ;
        RECT 2910.105 345.760 2910.275 346.285 ;
        RECT 2910.105 340.320 2910.275 340.845 ;
        RECT 2910.105 334.880 2910.275 335.405 ;
        RECT 2910.105 329.440 2910.275 329.965 ;
        RECT 2910.105 324.000 2910.275 324.525 ;
        RECT 2910.105 318.560 2910.275 319.085 ;
        RECT 2910.105 313.120 2910.275 313.645 ;
        RECT 2910.105 307.680 2910.275 308.205 ;
        RECT 2910.105 302.240 2910.275 302.765 ;
        RECT 2910.105 296.800 2910.275 297.325 ;
        RECT 2910.105 291.360 2910.275 291.885 ;
        RECT 2910.105 285.920 2910.275 286.445 ;
        RECT 2910.105 280.480 2910.275 281.005 ;
        RECT 2910.105 275.040 2910.275 275.565 ;
        RECT 2910.105 269.600 2910.275 270.125 ;
        RECT 2910.105 264.160 2910.275 264.685 ;
        RECT 2910.105 258.720 2910.275 259.245 ;
        RECT 2910.105 253.280 2910.275 253.805 ;
        RECT 2910.105 247.840 2910.275 248.365 ;
        RECT 2910.105 242.400 2910.275 242.925 ;
        RECT 2910.105 236.960 2910.275 237.485 ;
        RECT 2910.105 231.520 2910.275 232.045 ;
        RECT 2910.105 226.080 2910.275 226.605 ;
        RECT 2910.105 220.640 2910.275 221.165 ;
        RECT 2910.105 215.200 2910.275 215.725 ;
        RECT 2910.105 209.760 2910.275 210.285 ;
        RECT 2910.105 204.320 2910.275 204.845 ;
        RECT 2910.105 198.880 2910.275 199.405 ;
        RECT 2910.105 193.440 2910.275 193.965 ;
        RECT 2910.105 188.000 2910.275 188.525 ;
        RECT 2910.105 182.560 2910.275 183.085 ;
        RECT 2910.105 177.120 2910.275 177.645 ;
        RECT 2910.105 171.680 2910.275 172.205 ;
        RECT 2910.105 166.240 2910.275 166.765 ;
        RECT 2910.105 160.800 2910.275 161.325 ;
        RECT 2910.105 155.360 2910.275 155.885 ;
        RECT 2910.105 149.920 2910.275 150.445 ;
        RECT 2910.105 144.480 2910.275 145.005 ;
        RECT 2910.105 139.040 2910.275 139.565 ;
        RECT 2910.105 133.600 2910.275 134.125 ;
        RECT 2910.105 128.160 2910.275 128.685 ;
        RECT 2910.105 122.720 2910.275 123.245 ;
        RECT 2910.105 117.280 2910.275 117.805 ;
        RECT 2910.105 111.840 2910.275 112.365 ;
        RECT 2910.105 106.400 2910.275 106.925 ;
        RECT 2910.105 100.960 2910.275 101.485 ;
        RECT 2910.105 95.520 2910.275 96.045 ;
        RECT 2910.105 90.080 2910.275 90.605 ;
        RECT 2910.105 84.640 2910.275 85.165 ;
        RECT 2910.105 79.200 2910.275 79.725 ;
        RECT 2910.105 73.760 2910.275 74.285 ;
        RECT 2910.105 68.320 2910.275 68.845 ;
        RECT 2910.105 62.880 2910.275 63.405 ;
        RECT 2910.105 57.440 2910.275 57.965 ;
        RECT 2910.105 52.000 2910.275 52.525 ;
        RECT 2910.105 46.560 2910.275 47.085 ;
        RECT 2910.105 41.120 2910.275 41.645 ;
        RECT 2910.105 35.680 2910.275 36.205 ;
        RECT 2910.105 30.240 2910.275 30.765 ;
        RECT 2910.105 24.800 2910.275 25.325 ;
        RECT 2910.105 19.360 2910.275 19.885 ;
        RECT 2910.105 13.920 2910.275 14.445 ;
        RECT 19.925 12.755 20.095 13.280 ;
        RECT 34.185 12.755 34.355 13.280 ;
        RECT 48.445 12.755 48.615 13.280 ;
        RECT 62.705 12.755 62.875 13.280 ;
        RECT 76.965 12.755 77.135 13.280 ;
        RECT 91.225 12.755 91.395 13.280 ;
        RECT 105.485 12.755 105.655 13.280 ;
        RECT 119.745 12.755 119.915 13.280 ;
        RECT 134.005 12.755 134.175 13.280 ;
        RECT 148.265 12.755 148.435 13.280 ;
        RECT 162.525 12.755 162.695 13.280 ;
        RECT 176.785 12.755 176.955 13.280 ;
        RECT 191.045 12.755 191.215 13.280 ;
        RECT 205.305 12.755 205.475 13.280 ;
        RECT 219.565 12.755 219.735 13.280 ;
        RECT 233.825 12.755 233.995 13.280 ;
        RECT 248.085 12.755 248.255 13.280 ;
        RECT 262.345 12.755 262.515 13.280 ;
        RECT 276.605 12.755 276.775 13.280 ;
        RECT 290.865 12.755 291.035 13.280 ;
        RECT 305.125 12.755 305.295 13.280 ;
        RECT 319.385 12.755 319.555 13.280 ;
        RECT 333.645 12.755 333.815 13.280 ;
        RECT 347.905 12.755 348.075 13.280 ;
        RECT 362.165 12.755 362.335 13.280 ;
        RECT 376.425 12.755 376.595 13.280 ;
        RECT 390.685 12.755 390.855 13.280 ;
        RECT 404.945 12.755 405.115 13.280 ;
        RECT 419.205 12.755 419.375 13.280 ;
        RECT 433.465 12.755 433.635 13.280 ;
        RECT 447.725 12.755 447.895 13.280 ;
        RECT 461.985 12.755 462.155 13.280 ;
        RECT 476.245 12.755 476.415 13.280 ;
        RECT 490.505 12.755 490.675 13.280 ;
        RECT 504.765 12.755 504.935 13.280 ;
        RECT 519.025 12.755 519.195 13.280 ;
        RECT 533.285 12.755 533.455 13.280 ;
        RECT 547.545 12.755 547.715 13.280 ;
        RECT 561.805 12.755 561.975 13.280 ;
        RECT 576.065 12.755 576.235 13.280 ;
        RECT 590.325 12.755 590.495 13.280 ;
        RECT 604.585 12.755 604.755 13.280 ;
        RECT 618.845 12.755 619.015 13.280 ;
        RECT 633.105 12.755 633.275 13.280 ;
        RECT 647.365 12.755 647.535 13.280 ;
        RECT 661.625 12.755 661.795 13.280 ;
        RECT 675.885 12.755 676.055 13.280 ;
        RECT 690.145 12.755 690.315 13.280 ;
        RECT 704.405 12.755 704.575 13.280 ;
        RECT 718.665 12.755 718.835 13.280 ;
        RECT 732.925 12.755 733.095 13.280 ;
        RECT 747.185 12.755 747.355 13.280 ;
        RECT 761.445 12.755 761.615 13.280 ;
        RECT 775.705 12.755 775.875 13.280 ;
        RECT 789.965 12.755 790.135 13.280 ;
        RECT 804.225 12.755 804.395 13.280 ;
        RECT 818.485 12.755 818.655 13.280 ;
        RECT 832.745 12.755 832.915 13.280 ;
        RECT 847.005 12.755 847.175 13.280 ;
        RECT 861.265 12.755 861.435 13.280 ;
        RECT 875.525 12.755 875.695 13.280 ;
        RECT 889.785 12.755 889.955 13.280 ;
        RECT 904.045 12.755 904.215 13.280 ;
        RECT 918.305 12.755 918.475 13.280 ;
        RECT 932.565 12.755 932.735 13.280 ;
        RECT 946.825 12.755 946.995 13.280 ;
        RECT 961.085 12.755 961.255 13.280 ;
        RECT 975.345 12.755 975.515 13.280 ;
        RECT 989.605 12.755 989.775 13.280 ;
        RECT 1003.865 12.755 1004.035 13.280 ;
        RECT 1018.125 12.755 1018.295 13.280 ;
        RECT 1032.385 12.755 1032.555 13.280 ;
        RECT 1046.645 12.755 1046.815 13.280 ;
        RECT 1060.905 12.755 1061.075 13.280 ;
        RECT 1075.165 12.755 1075.335 13.280 ;
        RECT 1089.425 12.755 1089.595 13.280 ;
        RECT 1103.685 12.755 1103.855 13.280 ;
        RECT 1117.945 12.755 1118.115 13.280 ;
        RECT 1132.205 12.755 1132.375 13.280 ;
        RECT 1146.465 12.755 1146.635 13.280 ;
        RECT 1160.725 12.755 1160.895 13.280 ;
        RECT 1174.985 12.755 1175.155 13.280 ;
        RECT 1189.245 12.755 1189.415 13.280 ;
        RECT 1203.505 12.755 1203.675 13.280 ;
        RECT 1217.765 12.755 1217.935 13.280 ;
        RECT 1232.025 12.755 1232.195 13.280 ;
        RECT 1246.285 12.755 1246.455 13.280 ;
        RECT 1260.545 12.755 1260.715 13.280 ;
        RECT 1274.805 12.755 1274.975 13.280 ;
        RECT 1289.065 12.755 1289.235 13.280 ;
        RECT 1303.325 12.755 1303.495 13.280 ;
        RECT 1317.585 12.755 1317.755 13.280 ;
        RECT 1331.845 12.755 1332.015 13.280 ;
        RECT 1346.105 12.755 1346.275 13.280 ;
        RECT 1360.365 12.755 1360.535 13.280 ;
        RECT 1374.625 12.755 1374.795 13.280 ;
        RECT 1388.885 12.755 1389.055 13.280 ;
        RECT 1403.145 12.755 1403.315 13.280 ;
        RECT 1417.405 12.755 1417.575 13.280 ;
        RECT 1431.665 12.755 1431.835 13.280 ;
        RECT 1445.925 12.755 1446.095 13.280 ;
        RECT 1460.185 12.755 1460.355 13.280 ;
        RECT 1474.445 12.755 1474.615 13.280 ;
        RECT 1488.705 12.755 1488.875 13.280 ;
        RECT 1502.965 12.755 1503.135 13.280 ;
        RECT 1517.225 12.755 1517.395 13.280 ;
        RECT 1531.485 12.755 1531.655 13.280 ;
        RECT 1545.745 12.755 1545.915 13.280 ;
        RECT 1560.005 12.755 1560.175 13.280 ;
        RECT 1574.265 12.755 1574.435 13.280 ;
        RECT 1588.525 12.755 1588.695 13.280 ;
        RECT 1602.785 12.755 1602.955 13.280 ;
        RECT 1617.045 12.755 1617.215 13.280 ;
        RECT 1631.305 12.755 1631.475 13.280 ;
        RECT 1645.565 12.755 1645.735 13.280 ;
        RECT 1659.825 12.755 1659.995 13.280 ;
        RECT 1674.085 12.755 1674.255 13.280 ;
        RECT 1688.345 12.755 1688.515 13.280 ;
        RECT 1702.605 12.755 1702.775 13.280 ;
        RECT 1716.865 12.755 1717.035 13.280 ;
        RECT 1731.125 12.755 1731.295 13.280 ;
        RECT 1745.385 12.755 1745.555 13.280 ;
        RECT 1759.645 12.755 1759.815 13.280 ;
        RECT 1773.905 12.755 1774.075 13.280 ;
        RECT 1788.165 12.755 1788.335 13.280 ;
        RECT 1802.425 12.755 1802.595 13.280 ;
        RECT 1816.685 12.755 1816.855 13.280 ;
        RECT 1830.945 12.755 1831.115 13.280 ;
        RECT 1845.205 12.755 1845.375 13.280 ;
        RECT 1859.465 12.755 1859.635 13.280 ;
        RECT 1873.725 12.755 1873.895 13.280 ;
        RECT 1887.985 12.755 1888.155 13.280 ;
        RECT 1902.245 12.755 1902.415 13.280 ;
        RECT 1916.505 12.755 1916.675 13.280 ;
        RECT 1930.765 12.755 1930.935 13.280 ;
        RECT 1945.025 12.755 1945.195 13.280 ;
        RECT 1959.285 12.755 1959.455 13.280 ;
        RECT 1973.545 12.755 1973.715 13.280 ;
        RECT 1987.805 12.755 1987.975 13.280 ;
        RECT 2002.065 12.755 2002.235 13.280 ;
        RECT 2016.325 12.755 2016.495 13.280 ;
        RECT 2030.585 12.755 2030.755 13.280 ;
        RECT 2044.845 12.755 2045.015 13.280 ;
        RECT 2059.105 12.755 2059.275 13.280 ;
        RECT 2073.365 12.755 2073.535 13.280 ;
        RECT 2087.625 12.755 2087.795 13.280 ;
        RECT 2101.885 12.755 2102.055 13.280 ;
        RECT 2116.145 12.755 2116.315 13.280 ;
        RECT 2130.405 12.755 2130.575 13.280 ;
        RECT 2144.665 12.755 2144.835 13.280 ;
        RECT 2158.925 12.755 2159.095 13.280 ;
        RECT 2173.185 12.755 2173.355 13.280 ;
        RECT 2187.445 12.755 2187.615 13.280 ;
        RECT 2201.705 12.755 2201.875 13.280 ;
        RECT 2215.965 12.755 2216.135 13.280 ;
        RECT 2230.225 12.755 2230.395 13.280 ;
        RECT 2244.485 12.755 2244.655 13.280 ;
        RECT 2258.745 12.755 2258.915 13.280 ;
        RECT 2273.005 12.755 2273.175 13.280 ;
        RECT 2287.265 12.755 2287.435 13.280 ;
        RECT 2301.525 12.755 2301.695 13.280 ;
        RECT 2315.785 12.755 2315.955 13.280 ;
        RECT 2330.045 12.755 2330.215 13.280 ;
        RECT 2344.305 12.755 2344.475 13.280 ;
        RECT 2358.565 12.755 2358.735 13.280 ;
        RECT 2372.825 12.755 2372.995 13.280 ;
        RECT 2387.085 12.755 2387.255 13.280 ;
        RECT 2401.345 12.755 2401.515 13.280 ;
        RECT 2415.605 12.755 2415.775 13.280 ;
        RECT 2429.865 12.755 2430.035 13.280 ;
        RECT 2444.125 12.755 2444.295 13.280 ;
        RECT 2458.385 12.755 2458.555 13.280 ;
        RECT 2472.645 12.755 2472.815 13.280 ;
        RECT 2486.905 12.755 2487.075 13.280 ;
        RECT 2501.165 12.755 2501.335 13.280 ;
        RECT 2515.425 12.755 2515.595 13.280 ;
        RECT 2529.685 12.755 2529.855 13.280 ;
        RECT 2543.945 12.755 2544.115 13.280 ;
        RECT 2558.205 12.755 2558.375 13.280 ;
        RECT 2572.465 12.755 2572.635 13.280 ;
        RECT 2586.725 12.755 2586.895 13.280 ;
        RECT 2600.985 12.755 2601.155 13.280 ;
        RECT 2615.245 12.755 2615.415 13.280 ;
        RECT 2629.505 12.755 2629.675 13.280 ;
        RECT 2643.765 12.755 2643.935 13.280 ;
        RECT 2658.025 12.755 2658.195 13.280 ;
        RECT 2672.285 12.755 2672.455 13.280 ;
        RECT 2686.545 12.755 2686.715 13.280 ;
        RECT 2700.805 12.755 2700.975 13.280 ;
        RECT 2715.065 12.755 2715.235 13.280 ;
        RECT 2729.325 12.755 2729.495 13.280 ;
        RECT 2743.585 12.755 2743.755 13.280 ;
        RECT 2757.845 12.755 2758.015 13.280 ;
        RECT 2772.105 12.755 2772.275 13.280 ;
        RECT 2786.365 12.755 2786.535 13.280 ;
        RECT 2800.625 12.755 2800.795 13.280 ;
        RECT 2814.885 12.755 2815.055 13.280 ;
        RECT 2829.145 12.755 2829.315 13.280 ;
        RECT 2843.405 12.755 2843.575 13.280 ;
        RECT 2857.665 12.755 2857.835 13.280 ;
        RECT 2871.925 12.755 2872.095 13.280 ;
        RECT 2886.185 12.755 2886.355 13.280 ;
        RECT 2900.445 12.755 2900.615 13.280 ;
      LAYER li1 ;
        RECT 5.605 3506.915 6.125 3507.455 ;
        RECT 2913.495 3506.915 2914.015 3507.455 ;
        RECT 5.605 3506.165 6.815 3506.915 ;
        RECT 19.865 3506.300 20.155 3506.890 ;
        RECT 34.125 3506.300 34.415 3506.890 ;
        RECT 48.385 3506.300 48.675 3506.890 ;
        RECT 62.645 3506.300 62.935 3506.890 ;
        RECT 76.905 3506.300 77.195 3506.890 ;
        RECT 91.165 3506.300 91.455 3506.890 ;
        RECT 105.425 3506.300 105.715 3506.890 ;
        RECT 119.685 3506.300 119.975 3506.890 ;
        RECT 133.945 3506.300 134.235 3506.890 ;
        RECT 148.205 3506.300 148.495 3506.890 ;
        RECT 162.465 3506.300 162.755 3506.890 ;
        RECT 176.725 3506.300 177.015 3506.890 ;
        RECT 190.985 3506.300 191.275 3506.890 ;
        RECT 205.245 3506.300 205.535 3506.890 ;
        RECT 219.505 3506.300 219.795 3506.890 ;
        RECT 233.765 3506.300 234.055 3506.890 ;
        RECT 248.025 3506.300 248.315 3506.890 ;
        RECT 262.285 3506.300 262.575 3506.890 ;
        RECT 276.545 3506.300 276.835 3506.890 ;
        RECT 290.805 3506.300 291.095 3506.890 ;
        RECT 305.065 3506.300 305.355 3506.890 ;
        RECT 319.325 3506.300 319.615 3506.890 ;
        RECT 333.585 3506.300 333.875 3506.890 ;
        RECT 347.845 3506.300 348.135 3506.890 ;
        RECT 362.105 3506.300 362.395 3506.890 ;
        RECT 376.365 3506.300 376.655 3506.890 ;
        RECT 390.625 3506.300 390.915 3506.890 ;
        RECT 404.885 3506.300 405.175 3506.890 ;
        RECT 419.145 3506.300 419.435 3506.890 ;
        RECT 433.405 3506.300 433.695 3506.890 ;
        RECT 447.665 3506.300 447.955 3506.890 ;
        RECT 461.925 3506.300 462.215 3506.890 ;
        RECT 476.185 3506.300 476.475 3506.890 ;
        RECT 490.445 3506.300 490.735 3506.890 ;
        RECT 504.705 3506.300 504.995 3506.890 ;
        RECT 518.965 3506.300 519.255 3506.890 ;
        RECT 533.225 3506.300 533.515 3506.890 ;
        RECT 547.485 3506.300 547.775 3506.890 ;
        RECT 561.745 3506.300 562.035 3506.890 ;
        RECT 576.005 3506.300 576.295 3506.890 ;
        RECT 590.265 3506.300 590.555 3506.890 ;
        RECT 604.525 3506.300 604.815 3506.890 ;
        RECT 618.785 3506.300 619.075 3506.890 ;
        RECT 633.045 3506.300 633.335 3506.890 ;
        RECT 647.305 3506.300 647.595 3506.890 ;
        RECT 661.565 3506.300 661.855 3506.890 ;
        RECT 675.825 3506.300 676.115 3506.890 ;
        RECT 690.085 3506.300 690.375 3506.890 ;
        RECT 704.345 3506.300 704.635 3506.890 ;
        RECT 718.605 3506.300 718.895 3506.890 ;
        RECT 732.865 3506.300 733.155 3506.890 ;
        RECT 747.125 3506.300 747.415 3506.890 ;
        RECT 761.385 3506.300 761.675 3506.890 ;
        RECT 775.645 3506.300 775.935 3506.890 ;
        RECT 789.905 3506.300 790.195 3506.890 ;
        RECT 804.165 3506.300 804.455 3506.890 ;
        RECT 818.425 3506.300 818.715 3506.890 ;
        RECT 832.685 3506.300 832.975 3506.890 ;
        RECT 846.945 3506.300 847.235 3506.890 ;
        RECT 861.205 3506.300 861.495 3506.890 ;
        RECT 875.465 3506.300 875.755 3506.890 ;
        RECT 889.725 3506.300 890.015 3506.890 ;
        RECT 903.985 3506.300 904.275 3506.890 ;
        RECT 918.245 3506.300 918.535 3506.890 ;
        RECT 932.505 3506.300 932.795 3506.890 ;
        RECT 946.765 3506.300 947.055 3506.890 ;
        RECT 961.025 3506.300 961.315 3506.890 ;
        RECT 975.285 3506.300 975.575 3506.890 ;
        RECT 989.545 3506.300 989.835 3506.890 ;
        RECT 1003.805 3506.300 1004.095 3506.890 ;
        RECT 1018.065 3506.300 1018.355 3506.890 ;
        RECT 1032.325 3506.300 1032.615 3506.890 ;
        RECT 1046.585 3506.300 1046.875 3506.890 ;
        RECT 1060.845 3506.300 1061.135 3506.890 ;
        RECT 1075.105 3506.300 1075.395 3506.890 ;
        RECT 1089.365 3506.300 1089.655 3506.890 ;
        RECT 1103.625 3506.300 1103.915 3506.890 ;
        RECT 1117.885 3506.300 1118.175 3506.890 ;
        RECT 1132.145 3506.300 1132.435 3506.890 ;
        RECT 1146.405 3506.300 1146.695 3506.890 ;
        RECT 1160.665 3506.300 1160.955 3506.890 ;
        RECT 1174.925 3506.300 1175.215 3506.890 ;
        RECT 1189.185 3506.300 1189.475 3506.890 ;
        RECT 1203.445 3506.300 1203.735 3506.890 ;
        RECT 1217.705 3506.300 1217.995 3506.890 ;
        RECT 1231.965 3506.300 1232.255 3506.890 ;
        RECT 1246.225 3506.300 1246.515 3506.890 ;
        RECT 1260.485 3506.300 1260.775 3506.890 ;
        RECT 1274.745 3506.300 1275.035 3506.890 ;
        RECT 1289.005 3506.300 1289.295 3506.890 ;
        RECT 1303.265 3506.300 1303.555 3506.890 ;
        RECT 1317.525 3506.300 1317.815 3506.890 ;
        RECT 1331.785 3506.300 1332.075 3506.890 ;
        RECT 1346.045 3506.300 1346.335 3506.890 ;
        RECT 1360.305 3506.300 1360.595 3506.890 ;
        RECT 1374.565 3506.300 1374.855 3506.890 ;
        RECT 1388.825 3506.300 1389.115 3506.890 ;
        RECT 1403.085 3506.300 1403.375 3506.890 ;
        RECT 1417.345 3506.300 1417.635 3506.890 ;
        RECT 1431.605 3506.300 1431.895 3506.890 ;
        RECT 1445.865 3506.300 1446.155 3506.890 ;
        RECT 1460.125 3506.300 1460.415 3506.890 ;
        RECT 1474.385 3506.300 1474.675 3506.890 ;
        RECT 1488.645 3506.300 1488.935 3506.890 ;
        RECT 1502.905 3506.300 1503.195 3506.890 ;
        RECT 1517.165 3506.300 1517.455 3506.890 ;
        RECT 1531.425 3506.300 1531.715 3506.890 ;
        RECT 1545.685 3506.300 1545.975 3506.890 ;
        RECT 1559.945 3506.300 1560.235 3506.890 ;
        RECT 1574.205 3506.300 1574.495 3506.890 ;
        RECT 1588.465 3506.300 1588.755 3506.890 ;
        RECT 1602.725 3506.300 1603.015 3506.890 ;
        RECT 1616.985 3506.300 1617.275 3506.890 ;
        RECT 1631.245 3506.300 1631.535 3506.890 ;
        RECT 1645.505 3506.300 1645.795 3506.890 ;
        RECT 1659.765 3506.300 1660.055 3506.890 ;
        RECT 1674.025 3506.300 1674.315 3506.890 ;
        RECT 1688.285 3506.300 1688.575 3506.890 ;
        RECT 1702.545 3506.300 1702.835 3506.890 ;
        RECT 1716.805 3506.300 1717.095 3506.890 ;
        RECT 1731.065 3506.300 1731.355 3506.890 ;
        RECT 1745.325 3506.300 1745.615 3506.890 ;
        RECT 1759.585 3506.300 1759.875 3506.890 ;
        RECT 1773.845 3506.300 1774.135 3506.890 ;
        RECT 1788.105 3506.300 1788.395 3506.890 ;
        RECT 1802.365 3506.300 1802.655 3506.890 ;
        RECT 1816.625 3506.300 1816.915 3506.890 ;
        RECT 1830.885 3506.300 1831.175 3506.890 ;
        RECT 1845.145 3506.300 1845.435 3506.890 ;
        RECT 1859.405 3506.300 1859.695 3506.890 ;
        RECT 1873.665 3506.300 1873.955 3506.890 ;
        RECT 1887.925 3506.300 1888.215 3506.890 ;
        RECT 1902.185 3506.300 1902.475 3506.890 ;
        RECT 1916.445 3506.300 1916.735 3506.890 ;
        RECT 1930.705 3506.300 1930.995 3506.890 ;
        RECT 1944.965 3506.300 1945.255 3506.890 ;
        RECT 1959.225 3506.300 1959.515 3506.890 ;
        RECT 1973.485 3506.300 1973.775 3506.890 ;
        RECT 1987.745 3506.300 1988.035 3506.890 ;
        RECT 2002.005 3506.300 2002.295 3506.890 ;
        RECT 2016.265 3506.300 2016.555 3506.890 ;
        RECT 2030.525 3506.300 2030.815 3506.890 ;
        RECT 2044.785 3506.300 2045.075 3506.890 ;
        RECT 2059.045 3506.300 2059.335 3506.890 ;
        RECT 2073.305 3506.300 2073.595 3506.890 ;
        RECT 2087.565 3506.300 2087.855 3506.890 ;
        RECT 2101.825 3506.300 2102.115 3506.890 ;
        RECT 2116.085 3506.300 2116.375 3506.890 ;
        RECT 2130.345 3506.300 2130.635 3506.890 ;
        RECT 2144.605 3506.300 2144.895 3506.890 ;
        RECT 2158.865 3506.300 2159.155 3506.890 ;
        RECT 2173.125 3506.300 2173.415 3506.890 ;
        RECT 2187.385 3506.300 2187.675 3506.890 ;
        RECT 2201.645 3506.300 2201.935 3506.890 ;
        RECT 2215.905 3506.300 2216.195 3506.890 ;
        RECT 2230.165 3506.300 2230.455 3506.890 ;
        RECT 2244.425 3506.300 2244.715 3506.890 ;
        RECT 2258.685 3506.300 2258.975 3506.890 ;
        RECT 2272.945 3506.300 2273.235 3506.890 ;
        RECT 2287.205 3506.300 2287.495 3506.890 ;
        RECT 2301.465 3506.300 2301.755 3506.890 ;
        RECT 2315.725 3506.300 2316.015 3506.890 ;
        RECT 2329.985 3506.300 2330.275 3506.890 ;
        RECT 2344.245 3506.300 2344.535 3506.890 ;
        RECT 2358.505 3506.300 2358.795 3506.890 ;
        RECT 2372.765 3506.300 2373.055 3506.890 ;
        RECT 2387.025 3506.300 2387.315 3506.890 ;
        RECT 2401.285 3506.300 2401.575 3506.890 ;
        RECT 2415.545 3506.300 2415.835 3506.890 ;
        RECT 2429.805 3506.300 2430.095 3506.890 ;
        RECT 2444.065 3506.300 2444.355 3506.890 ;
        RECT 2458.325 3506.300 2458.615 3506.890 ;
        RECT 2472.585 3506.300 2472.875 3506.890 ;
        RECT 2486.845 3506.300 2487.135 3506.890 ;
        RECT 2501.105 3506.300 2501.395 3506.890 ;
        RECT 2515.365 3506.300 2515.655 3506.890 ;
        RECT 2529.625 3506.300 2529.915 3506.890 ;
        RECT 2543.885 3506.300 2544.175 3506.890 ;
        RECT 2558.145 3506.300 2558.435 3506.890 ;
        RECT 2572.405 3506.300 2572.695 3506.890 ;
        RECT 2586.665 3506.300 2586.955 3506.890 ;
        RECT 2600.925 3506.300 2601.215 3506.890 ;
        RECT 2615.185 3506.300 2615.475 3506.890 ;
        RECT 2629.445 3506.300 2629.735 3506.890 ;
        RECT 2643.705 3506.300 2643.995 3506.890 ;
        RECT 2657.965 3506.300 2658.255 3506.890 ;
        RECT 2672.225 3506.300 2672.515 3506.890 ;
        RECT 2686.485 3506.300 2686.775 3506.890 ;
        RECT 2700.745 3506.300 2701.035 3506.890 ;
        RECT 2715.005 3506.300 2715.295 3506.890 ;
        RECT 2729.265 3506.300 2729.555 3506.890 ;
        RECT 2743.525 3506.300 2743.815 3506.890 ;
        RECT 2757.785 3506.300 2758.075 3506.890 ;
        RECT 2772.045 3506.300 2772.335 3506.890 ;
        RECT 2786.305 3506.300 2786.595 3506.890 ;
        RECT 2800.565 3506.300 2800.855 3506.890 ;
        RECT 2814.825 3506.300 2815.115 3506.890 ;
        RECT 2829.085 3506.300 2829.375 3506.890 ;
        RECT 2843.345 3506.300 2843.635 3506.890 ;
        RECT 2857.605 3506.300 2857.895 3506.890 ;
        RECT 2871.865 3506.300 2872.155 3506.890 ;
        RECT 2886.125 3506.300 2886.415 3506.890 ;
        RECT 2900.385 3506.300 2900.675 3506.890 ;
        RECT 2912.805 3506.165 2914.015 3506.915 ;
        RECT 5.520 3505.995 6.900 3506.165 ;
        RECT 9.660 3505.995 12.420 3506.165 ;
        RECT 2909.040 3505.995 2911.800 3506.165 ;
        RECT 2912.720 3505.995 2914.100 3506.165 ;
        RECT 5.605 3505.245 6.815 3505.995 ;
        RECT 10.435 3505.335 10.775 3505.995 ;
        RECT 11.815 3505.335 12.155 3505.995 ;
        RECT 2909.815 3505.335 2910.155 3505.995 ;
        RECT 2911.195 3505.335 2911.535 3505.995 ;
        RECT 2912.805 3505.245 2914.015 3505.995 ;
        RECT 5.605 3504.705 6.125 3505.245 ;
        RECT 2913.495 3504.705 2914.015 3505.245 ;
        RECT 5.605 3501.475 6.125 3502.015 ;
        RECT 2913.495 3501.475 2914.015 3502.015 ;
        RECT 5.605 3500.725 6.815 3501.475 ;
        RECT 2910.045 3500.725 2910.335 3501.450 ;
        RECT 2912.805 3500.725 2914.015 3501.475 ;
        RECT 5.520 3500.555 6.900 3500.725 ;
        RECT 2909.960 3500.555 2910.420 3500.725 ;
        RECT 2912.720 3500.555 2914.100 3500.725 ;
        RECT 5.605 3499.805 6.815 3500.555 ;
        RECT 2912.805 3499.805 2914.015 3500.555 ;
        RECT 5.605 3499.265 6.125 3499.805 ;
        RECT 2913.495 3499.265 2914.015 3499.805 ;
        RECT 5.605 3496.035 6.125 3496.575 ;
        RECT 2913.495 3496.035 2914.015 3496.575 ;
        RECT 5.605 3495.285 6.815 3496.035 ;
        RECT 2910.045 3495.285 2910.335 3496.010 ;
        RECT 2912.805 3495.285 2914.015 3496.035 ;
        RECT 5.520 3495.115 6.900 3495.285 ;
        RECT 2909.960 3495.115 2910.420 3495.285 ;
        RECT 2912.720 3495.115 2914.100 3495.285 ;
        RECT 5.605 3494.365 6.815 3495.115 ;
        RECT 2912.805 3494.365 2914.015 3495.115 ;
        RECT 5.605 3493.825 6.125 3494.365 ;
        RECT 2913.495 3493.825 2914.015 3494.365 ;
        RECT 5.605 3490.595 6.125 3491.135 ;
        RECT 2913.495 3490.595 2914.015 3491.135 ;
        RECT 5.605 3489.845 6.815 3490.595 ;
        RECT 2910.045 3489.845 2910.335 3490.570 ;
        RECT 2912.805 3489.845 2914.015 3490.595 ;
        RECT 5.520 3489.675 6.900 3489.845 ;
        RECT 2909.960 3489.675 2910.420 3489.845 ;
        RECT 2912.720 3489.675 2914.100 3489.845 ;
        RECT 5.605 3488.925 6.815 3489.675 ;
        RECT 2912.805 3488.925 2914.015 3489.675 ;
        RECT 5.605 3488.385 6.125 3488.925 ;
        RECT 2913.495 3488.385 2914.015 3488.925 ;
        RECT 5.605 3485.155 6.125 3485.695 ;
        RECT 2913.495 3485.155 2914.015 3485.695 ;
        RECT 5.605 3484.405 6.815 3485.155 ;
        RECT 2910.045 3484.405 2910.335 3485.130 ;
        RECT 2912.805 3484.405 2914.015 3485.155 ;
        RECT 5.520 3484.235 6.900 3484.405 ;
        RECT 2909.960 3484.235 2910.420 3484.405 ;
        RECT 2912.720 3484.235 2914.100 3484.405 ;
        RECT 5.605 3483.485 6.815 3484.235 ;
        RECT 2912.805 3483.485 2914.015 3484.235 ;
        RECT 5.605 3482.945 6.125 3483.485 ;
        RECT 2913.495 3482.945 2914.015 3483.485 ;
        RECT 5.605 3479.715 6.125 3480.255 ;
        RECT 2913.495 3479.715 2914.015 3480.255 ;
        RECT 5.605 3478.965 6.815 3479.715 ;
        RECT 2910.045 3478.965 2910.335 3479.690 ;
        RECT 2912.805 3478.965 2914.015 3479.715 ;
        RECT 5.520 3478.795 6.900 3478.965 ;
        RECT 2909.960 3478.795 2910.420 3478.965 ;
        RECT 2912.720 3478.795 2914.100 3478.965 ;
        RECT 5.605 3478.045 6.815 3478.795 ;
        RECT 2912.805 3478.045 2914.015 3478.795 ;
        RECT 5.605 3477.505 6.125 3478.045 ;
        RECT 2913.495 3477.505 2914.015 3478.045 ;
        RECT 5.605 3474.275 6.125 3474.815 ;
        RECT 2913.495 3474.275 2914.015 3474.815 ;
        RECT 5.605 3473.525 6.815 3474.275 ;
        RECT 2910.045 3473.525 2910.335 3474.250 ;
        RECT 2912.805 3473.525 2914.015 3474.275 ;
        RECT 5.520 3473.355 6.900 3473.525 ;
        RECT 2909.960 3473.355 2910.420 3473.525 ;
        RECT 2912.720 3473.355 2914.100 3473.525 ;
        RECT 5.605 3472.605 6.815 3473.355 ;
        RECT 2912.805 3472.605 2914.015 3473.355 ;
        RECT 5.605 3472.065 6.125 3472.605 ;
        RECT 2913.495 3472.065 2914.015 3472.605 ;
        RECT 5.605 3468.835 6.125 3469.375 ;
        RECT 2913.495 3468.835 2914.015 3469.375 ;
        RECT 5.605 3468.085 6.815 3468.835 ;
        RECT 2910.045 3468.085 2910.335 3468.810 ;
        RECT 2912.805 3468.085 2914.015 3468.835 ;
        RECT 5.520 3467.915 6.900 3468.085 ;
        RECT 2909.960 3467.915 2910.420 3468.085 ;
        RECT 2912.720 3467.915 2914.100 3468.085 ;
        RECT 5.605 3467.165 6.815 3467.915 ;
        RECT 2912.805 3467.165 2914.015 3467.915 ;
        RECT 5.605 3466.625 6.125 3467.165 ;
        RECT 2913.495 3466.625 2914.015 3467.165 ;
        RECT 5.605 3463.395 6.125 3463.935 ;
        RECT 2913.495 3463.395 2914.015 3463.935 ;
        RECT 5.605 3462.645 6.815 3463.395 ;
        RECT 2910.045 3462.645 2910.335 3463.370 ;
        RECT 2912.805 3462.645 2914.015 3463.395 ;
        RECT 5.520 3462.475 6.900 3462.645 ;
        RECT 2909.960 3462.475 2910.420 3462.645 ;
        RECT 2912.720 3462.475 2914.100 3462.645 ;
        RECT 5.605 3461.725 6.815 3462.475 ;
        RECT 2912.805 3461.725 2914.015 3462.475 ;
        RECT 5.605 3461.185 6.125 3461.725 ;
        RECT 2913.495 3461.185 2914.015 3461.725 ;
        RECT 5.605 3457.955 6.125 3458.495 ;
        RECT 2913.495 3457.955 2914.015 3458.495 ;
        RECT 5.605 3457.205 6.815 3457.955 ;
        RECT 2910.045 3457.205 2910.335 3457.930 ;
        RECT 2912.805 3457.205 2914.015 3457.955 ;
        RECT 5.520 3457.035 6.900 3457.205 ;
        RECT 2909.960 3457.035 2910.420 3457.205 ;
        RECT 2912.720 3457.035 2914.100 3457.205 ;
        RECT 5.605 3456.285 6.815 3457.035 ;
        RECT 2912.805 3456.285 2914.015 3457.035 ;
        RECT 5.605 3455.745 6.125 3456.285 ;
        RECT 2913.495 3455.745 2914.015 3456.285 ;
        RECT 5.605 3452.515 6.125 3453.055 ;
        RECT 2913.495 3452.515 2914.015 3453.055 ;
        RECT 5.605 3451.765 6.815 3452.515 ;
        RECT 2910.045 3451.765 2910.335 3452.490 ;
        RECT 2912.805 3451.765 2914.015 3452.515 ;
        RECT 5.520 3451.595 6.900 3451.765 ;
        RECT 2909.960 3451.595 2910.420 3451.765 ;
        RECT 2912.720 3451.595 2914.100 3451.765 ;
        RECT 5.605 3450.845 6.815 3451.595 ;
        RECT 2912.805 3450.845 2914.015 3451.595 ;
        RECT 5.605 3450.305 6.125 3450.845 ;
        RECT 2913.495 3450.305 2914.015 3450.845 ;
        RECT 5.605 3447.075 6.125 3447.615 ;
        RECT 2913.495 3447.075 2914.015 3447.615 ;
        RECT 5.605 3446.325 6.815 3447.075 ;
        RECT 2910.045 3446.325 2910.335 3447.050 ;
        RECT 2912.805 3446.325 2914.015 3447.075 ;
        RECT 5.520 3446.155 6.900 3446.325 ;
        RECT 2909.960 3446.155 2910.420 3446.325 ;
        RECT 2912.720 3446.155 2914.100 3446.325 ;
        RECT 5.605 3445.405 6.815 3446.155 ;
        RECT 2912.805 3445.405 2914.015 3446.155 ;
        RECT 5.605 3444.865 6.125 3445.405 ;
        RECT 2913.495 3444.865 2914.015 3445.405 ;
        RECT 5.605 3441.635 6.125 3442.175 ;
        RECT 2913.495 3441.635 2914.015 3442.175 ;
        RECT 5.605 3440.885 6.815 3441.635 ;
        RECT 2910.045 3440.885 2910.335 3441.610 ;
        RECT 2912.805 3440.885 2914.015 3441.635 ;
        RECT 5.520 3440.715 6.900 3440.885 ;
        RECT 2909.960 3440.715 2910.420 3440.885 ;
        RECT 2912.720 3440.715 2914.100 3440.885 ;
        RECT 5.605 3439.965 6.815 3440.715 ;
        RECT 2912.805 3439.965 2914.015 3440.715 ;
        RECT 5.605 3439.425 6.125 3439.965 ;
        RECT 2913.495 3439.425 2914.015 3439.965 ;
        RECT 5.605 3436.195 6.125 3436.735 ;
        RECT 2913.495 3436.195 2914.015 3436.735 ;
        RECT 5.605 3435.445 6.815 3436.195 ;
        RECT 2910.045 3435.445 2910.335 3436.170 ;
        RECT 2912.805 3435.445 2914.015 3436.195 ;
        RECT 5.520 3435.275 6.900 3435.445 ;
        RECT 2909.960 3435.275 2910.420 3435.445 ;
        RECT 2912.720 3435.275 2914.100 3435.445 ;
        RECT 5.605 3434.525 6.815 3435.275 ;
        RECT 2912.805 3434.525 2914.015 3435.275 ;
        RECT 5.605 3433.985 6.125 3434.525 ;
        RECT 2913.495 3433.985 2914.015 3434.525 ;
        RECT 5.605 3430.755 6.125 3431.295 ;
        RECT 2913.495 3430.755 2914.015 3431.295 ;
        RECT 5.605 3430.005 6.815 3430.755 ;
        RECT 2910.045 3430.005 2910.335 3430.730 ;
        RECT 2912.805 3430.005 2914.015 3430.755 ;
        RECT 5.520 3429.835 6.900 3430.005 ;
        RECT 2909.960 3429.835 2910.420 3430.005 ;
        RECT 2912.720 3429.835 2914.100 3430.005 ;
        RECT 5.605 3429.085 6.815 3429.835 ;
        RECT 2912.805 3429.085 2914.015 3429.835 ;
        RECT 5.605 3428.545 6.125 3429.085 ;
        RECT 2913.495 3428.545 2914.015 3429.085 ;
        RECT 5.605 3425.315 6.125 3425.855 ;
        RECT 2913.495 3425.315 2914.015 3425.855 ;
        RECT 5.605 3424.565 6.815 3425.315 ;
        RECT 2910.045 3424.565 2910.335 3425.290 ;
        RECT 2912.805 3424.565 2914.015 3425.315 ;
        RECT 5.520 3424.395 6.900 3424.565 ;
        RECT 2909.960 3424.395 2910.420 3424.565 ;
        RECT 2912.720 3424.395 2914.100 3424.565 ;
        RECT 5.605 3423.645 6.815 3424.395 ;
        RECT 2912.805 3423.645 2914.015 3424.395 ;
        RECT 5.605 3423.105 6.125 3423.645 ;
        RECT 2913.495 3423.105 2914.015 3423.645 ;
        RECT 5.605 3419.875 6.125 3420.415 ;
        RECT 2913.495 3419.875 2914.015 3420.415 ;
        RECT 5.605 3419.125 6.815 3419.875 ;
        RECT 2910.045 3419.125 2910.335 3419.850 ;
        RECT 2912.805 3419.125 2914.015 3419.875 ;
        RECT 5.520 3418.955 6.900 3419.125 ;
        RECT 2909.960 3418.955 2910.420 3419.125 ;
        RECT 2912.720 3418.955 2914.100 3419.125 ;
        RECT 5.605 3418.205 6.815 3418.955 ;
        RECT 2912.805 3418.205 2914.015 3418.955 ;
        RECT 5.605 3417.665 6.125 3418.205 ;
        RECT 2913.495 3417.665 2914.015 3418.205 ;
        RECT 5.605 3414.435 6.125 3414.975 ;
        RECT 2913.495 3414.435 2914.015 3414.975 ;
        RECT 5.605 3413.685 6.815 3414.435 ;
        RECT 2910.045 3413.685 2910.335 3414.410 ;
        RECT 2912.805 3413.685 2914.015 3414.435 ;
        RECT 5.520 3413.515 6.900 3413.685 ;
        RECT 2909.960 3413.515 2910.420 3413.685 ;
        RECT 2912.720 3413.515 2914.100 3413.685 ;
        RECT 5.605 3412.765 6.815 3413.515 ;
        RECT 2912.805 3412.765 2914.015 3413.515 ;
        RECT 5.605 3412.225 6.125 3412.765 ;
        RECT 2913.495 3412.225 2914.015 3412.765 ;
        RECT 5.605 3408.995 6.125 3409.535 ;
        RECT 2913.495 3408.995 2914.015 3409.535 ;
        RECT 5.605 3408.245 6.815 3408.995 ;
        RECT 2910.045 3408.245 2910.335 3408.970 ;
        RECT 2912.805 3408.245 2914.015 3408.995 ;
        RECT 5.520 3408.075 6.900 3408.245 ;
        RECT 2909.960 3408.075 2910.420 3408.245 ;
        RECT 2912.720 3408.075 2914.100 3408.245 ;
        RECT 5.605 3407.325 6.815 3408.075 ;
        RECT 2912.805 3407.325 2914.015 3408.075 ;
        RECT 5.605 3406.785 6.125 3407.325 ;
        RECT 2913.495 3406.785 2914.015 3407.325 ;
        RECT 5.605 3403.555 6.125 3404.095 ;
        RECT 2913.495 3403.555 2914.015 3404.095 ;
        RECT 5.605 3402.805 6.815 3403.555 ;
        RECT 2910.045 3402.805 2910.335 3403.530 ;
        RECT 2912.805 3402.805 2914.015 3403.555 ;
        RECT 5.520 3402.635 6.900 3402.805 ;
        RECT 2909.040 3402.635 2910.420 3402.805 ;
        RECT 2912.720 3402.635 2914.100 3402.805 ;
        RECT 5.605 3401.885 6.815 3402.635 ;
        RECT 2909.815 3401.975 2910.155 3402.635 ;
        RECT 2912.805 3401.885 2914.015 3402.635 ;
        RECT 5.605 3401.345 6.125 3401.885 ;
        RECT 2913.495 3401.345 2914.015 3401.885 ;
        RECT 5.605 3398.115 6.125 3398.655 ;
        RECT 2913.495 3398.115 2914.015 3398.655 ;
        RECT 5.605 3397.365 6.815 3398.115 ;
        RECT 2910.045 3397.365 2910.335 3398.090 ;
        RECT 2912.805 3397.365 2914.015 3398.115 ;
        RECT 5.520 3397.195 6.900 3397.365 ;
        RECT 2909.960 3397.195 2910.420 3397.365 ;
        RECT 2912.720 3397.195 2914.100 3397.365 ;
        RECT 5.605 3396.445 6.815 3397.195 ;
        RECT 2912.805 3396.445 2914.015 3397.195 ;
        RECT 5.605 3395.905 6.125 3396.445 ;
        RECT 2913.495 3395.905 2914.015 3396.445 ;
        RECT 5.605 3392.675 6.125 3393.215 ;
        RECT 2913.495 3392.675 2914.015 3393.215 ;
        RECT 5.605 3391.925 6.815 3392.675 ;
        RECT 2910.045 3391.925 2910.335 3392.650 ;
        RECT 2912.805 3391.925 2914.015 3392.675 ;
        RECT 5.520 3391.755 6.900 3391.925 ;
        RECT 2909.960 3391.755 2910.420 3391.925 ;
        RECT 2912.720 3391.755 2914.100 3391.925 ;
        RECT 5.605 3391.005 6.815 3391.755 ;
        RECT 2912.805 3391.005 2914.015 3391.755 ;
        RECT 5.605 3390.465 6.125 3391.005 ;
        RECT 2913.495 3390.465 2914.015 3391.005 ;
        RECT 5.605 3387.235 6.125 3387.775 ;
        RECT 2913.495 3387.235 2914.015 3387.775 ;
        RECT 5.605 3386.485 6.815 3387.235 ;
        RECT 2910.045 3386.485 2910.335 3387.210 ;
        RECT 2912.805 3386.485 2914.015 3387.235 ;
        RECT 5.520 3386.315 6.900 3386.485 ;
        RECT 2909.960 3386.315 2910.420 3386.485 ;
        RECT 2912.720 3386.315 2914.100 3386.485 ;
        RECT 5.605 3385.565 6.815 3386.315 ;
        RECT 2912.805 3385.565 2914.015 3386.315 ;
        RECT 5.605 3385.025 6.125 3385.565 ;
        RECT 2913.495 3385.025 2914.015 3385.565 ;
        RECT 5.605 3381.795 6.125 3382.335 ;
        RECT 2913.495 3381.795 2914.015 3382.335 ;
        RECT 5.605 3381.045 6.815 3381.795 ;
        RECT 2910.045 3381.045 2910.335 3381.770 ;
        RECT 2912.805 3381.045 2914.015 3381.795 ;
        RECT 5.520 3380.875 6.900 3381.045 ;
        RECT 2909.960 3380.875 2910.420 3381.045 ;
        RECT 2912.720 3380.875 2914.100 3381.045 ;
        RECT 5.605 3380.125 6.815 3380.875 ;
        RECT 2912.805 3380.125 2914.015 3380.875 ;
        RECT 5.605 3379.585 6.125 3380.125 ;
        RECT 2913.495 3379.585 2914.015 3380.125 ;
        RECT 5.605 3376.355 6.125 3376.895 ;
        RECT 2913.495 3376.355 2914.015 3376.895 ;
        RECT 5.605 3375.605 6.815 3376.355 ;
        RECT 2910.045 3375.605 2910.335 3376.330 ;
        RECT 2912.805 3375.605 2914.015 3376.355 ;
        RECT 5.520 3375.435 6.900 3375.605 ;
        RECT 2909.960 3375.435 2910.420 3375.605 ;
        RECT 2912.720 3375.435 2914.100 3375.605 ;
        RECT 5.605 3374.685 6.815 3375.435 ;
        RECT 2912.805 3374.685 2914.015 3375.435 ;
        RECT 5.605 3374.145 6.125 3374.685 ;
        RECT 2913.495 3374.145 2914.015 3374.685 ;
        RECT 5.605 3370.915 6.125 3371.455 ;
        RECT 2913.495 3370.915 2914.015 3371.455 ;
        RECT 5.605 3370.165 6.815 3370.915 ;
        RECT 2910.045 3370.165 2910.335 3370.890 ;
        RECT 2912.805 3370.165 2914.015 3370.915 ;
        RECT 5.520 3369.995 6.900 3370.165 ;
        RECT 2909.960 3369.995 2910.420 3370.165 ;
        RECT 2912.720 3369.995 2914.100 3370.165 ;
        RECT 5.605 3369.245 6.815 3369.995 ;
        RECT 2912.805 3369.245 2914.015 3369.995 ;
        RECT 5.605 3368.705 6.125 3369.245 ;
        RECT 2913.495 3368.705 2914.015 3369.245 ;
        RECT 5.605 3365.475 6.125 3366.015 ;
        RECT 2913.495 3365.475 2914.015 3366.015 ;
        RECT 5.605 3364.725 6.815 3365.475 ;
        RECT 2910.045 3364.725 2910.335 3365.450 ;
        RECT 2911.195 3364.725 2911.535 3365.385 ;
        RECT 2912.805 3364.725 2914.015 3365.475 ;
        RECT 5.520 3364.555 6.900 3364.725 ;
        RECT 2909.960 3364.555 2911.800 3364.725 ;
        RECT 2912.720 3364.555 2914.100 3364.725 ;
        RECT 5.605 3363.805 6.815 3364.555 ;
        RECT 2912.805 3363.805 2914.015 3364.555 ;
        RECT 5.605 3363.265 6.125 3363.805 ;
        RECT 2913.495 3363.265 2914.015 3363.805 ;
        RECT 5.605 3360.035 6.125 3360.575 ;
        RECT 2913.495 3360.035 2914.015 3360.575 ;
        RECT 5.605 3359.285 6.815 3360.035 ;
        RECT 2910.045 3359.285 2910.335 3360.010 ;
        RECT 2912.805 3359.285 2914.015 3360.035 ;
        RECT 5.520 3359.115 6.900 3359.285 ;
        RECT 2909.960 3359.115 2910.420 3359.285 ;
        RECT 2912.720 3359.115 2914.100 3359.285 ;
        RECT 5.605 3358.365 6.815 3359.115 ;
        RECT 2912.805 3358.365 2914.015 3359.115 ;
        RECT 5.605 3357.825 6.125 3358.365 ;
        RECT 2913.495 3357.825 2914.015 3358.365 ;
        RECT 5.605 3354.595 6.125 3355.135 ;
        RECT 2913.495 3354.595 2914.015 3355.135 ;
        RECT 5.605 3353.845 6.815 3354.595 ;
        RECT 2910.045 3353.845 2910.335 3354.570 ;
        RECT 2912.805 3353.845 2914.015 3354.595 ;
        RECT 5.520 3353.675 6.900 3353.845 ;
        RECT 2909.960 3353.675 2910.420 3353.845 ;
        RECT 2912.720 3353.675 2914.100 3353.845 ;
        RECT 5.605 3352.925 6.815 3353.675 ;
        RECT 2912.805 3352.925 2914.015 3353.675 ;
        RECT 5.605 3352.385 6.125 3352.925 ;
        RECT 2913.495 3352.385 2914.015 3352.925 ;
        RECT 5.605 3349.155 6.125 3349.695 ;
        RECT 2913.495 3349.155 2914.015 3349.695 ;
        RECT 5.605 3348.405 6.815 3349.155 ;
        RECT 2910.045 3348.405 2910.335 3349.130 ;
        RECT 2912.805 3348.405 2914.015 3349.155 ;
        RECT 5.520 3348.235 6.900 3348.405 ;
        RECT 2909.960 3348.235 2910.420 3348.405 ;
        RECT 2912.720 3348.235 2914.100 3348.405 ;
        RECT 5.605 3347.485 6.815 3348.235 ;
        RECT 2912.805 3347.485 2914.015 3348.235 ;
        RECT 5.605 3346.945 6.125 3347.485 ;
        RECT 2913.495 3346.945 2914.015 3347.485 ;
        RECT 5.605 3343.715 6.125 3344.255 ;
        RECT 2913.495 3343.715 2914.015 3344.255 ;
        RECT 5.605 3342.965 6.815 3343.715 ;
        RECT 2910.045 3342.965 2910.335 3343.690 ;
        RECT 2912.805 3342.965 2914.015 3343.715 ;
        RECT 5.520 3342.795 6.900 3342.965 ;
        RECT 2909.960 3342.795 2910.420 3342.965 ;
        RECT 2912.720 3342.795 2914.100 3342.965 ;
        RECT 5.605 3342.045 6.815 3342.795 ;
        RECT 2912.805 3342.045 2914.015 3342.795 ;
        RECT 5.605 3341.505 6.125 3342.045 ;
        RECT 2913.495 3341.505 2914.015 3342.045 ;
        RECT 5.605 3338.275 6.125 3338.815 ;
        RECT 2913.495 3338.275 2914.015 3338.815 ;
        RECT 5.605 3337.525 6.815 3338.275 ;
        RECT 2910.045 3337.525 2910.335 3338.250 ;
        RECT 2912.805 3337.525 2914.015 3338.275 ;
        RECT 5.520 3337.355 6.900 3337.525 ;
        RECT 2909.960 3337.355 2910.420 3337.525 ;
        RECT 2912.720 3337.355 2914.100 3337.525 ;
        RECT 5.605 3336.605 6.815 3337.355 ;
        RECT 2912.805 3336.605 2914.015 3337.355 ;
        RECT 5.605 3336.065 6.125 3336.605 ;
        RECT 2913.495 3336.065 2914.015 3336.605 ;
        RECT 5.605 3332.835 6.125 3333.375 ;
        RECT 2913.495 3332.835 2914.015 3333.375 ;
        RECT 5.605 3332.085 6.815 3332.835 ;
        RECT 2910.045 3332.085 2910.335 3332.810 ;
        RECT 2912.805 3332.085 2914.015 3332.835 ;
        RECT 5.520 3331.915 6.900 3332.085 ;
        RECT 2909.960 3331.915 2910.420 3332.085 ;
        RECT 2912.720 3331.915 2914.100 3332.085 ;
        RECT 5.605 3331.165 6.815 3331.915 ;
        RECT 2912.805 3331.165 2914.015 3331.915 ;
        RECT 5.605 3330.625 6.125 3331.165 ;
        RECT 2913.495 3330.625 2914.015 3331.165 ;
        RECT 5.605 3327.395 6.125 3327.935 ;
        RECT 2913.495 3327.395 2914.015 3327.935 ;
        RECT 5.605 3326.645 6.815 3327.395 ;
        RECT 2910.045 3326.645 2910.335 3327.370 ;
        RECT 2912.805 3326.645 2914.015 3327.395 ;
        RECT 5.520 3326.475 6.900 3326.645 ;
        RECT 2909.960 3326.475 2910.420 3326.645 ;
        RECT 2912.720 3326.475 2914.100 3326.645 ;
        RECT 5.605 3325.725 6.815 3326.475 ;
        RECT 2912.805 3325.725 2914.015 3326.475 ;
        RECT 5.605 3325.185 6.125 3325.725 ;
        RECT 2913.495 3325.185 2914.015 3325.725 ;
        RECT 5.605 3321.955 6.125 3322.495 ;
        RECT 2913.495 3321.955 2914.015 3322.495 ;
        RECT 5.605 3321.205 6.815 3321.955 ;
        RECT 2910.045 3321.205 2910.335 3321.930 ;
        RECT 2912.805 3321.205 2914.015 3321.955 ;
        RECT 5.520 3321.035 6.900 3321.205 ;
        RECT 2909.960 3321.035 2910.420 3321.205 ;
        RECT 2912.720 3321.035 2914.100 3321.205 ;
        RECT 5.605 3320.285 6.815 3321.035 ;
        RECT 2912.805 3320.285 2914.015 3321.035 ;
        RECT 5.605 3319.745 6.125 3320.285 ;
        RECT 2913.495 3319.745 2914.015 3320.285 ;
        RECT 5.605 3316.515 6.125 3317.055 ;
        RECT 2913.495 3316.515 2914.015 3317.055 ;
        RECT 5.605 3315.765 6.815 3316.515 ;
        RECT 2910.045 3315.765 2910.335 3316.490 ;
        RECT 2912.805 3315.765 2914.015 3316.515 ;
        RECT 5.520 3315.595 6.900 3315.765 ;
        RECT 2909.960 3315.595 2910.420 3315.765 ;
        RECT 2912.720 3315.595 2914.100 3315.765 ;
        RECT 5.605 3314.845 6.815 3315.595 ;
        RECT 2912.805 3314.845 2914.015 3315.595 ;
        RECT 5.605 3314.305 6.125 3314.845 ;
        RECT 2913.495 3314.305 2914.015 3314.845 ;
        RECT 5.605 3311.075 6.125 3311.615 ;
        RECT 2913.495 3311.075 2914.015 3311.615 ;
        RECT 5.605 3310.325 6.815 3311.075 ;
        RECT 2910.045 3310.325 2910.335 3311.050 ;
        RECT 2912.805 3310.325 2914.015 3311.075 ;
        RECT 5.520 3310.155 6.900 3310.325 ;
        RECT 2909.960 3310.155 2910.420 3310.325 ;
        RECT 2912.720 3310.155 2914.100 3310.325 ;
        RECT 5.605 3309.405 6.815 3310.155 ;
        RECT 2912.805 3309.405 2914.015 3310.155 ;
        RECT 5.605 3308.865 6.125 3309.405 ;
        RECT 2913.495 3308.865 2914.015 3309.405 ;
        RECT 5.605 3305.635 6.125 3306.175 ;
        RECT 2913.495 3305.635 2914.015 3306.175 ;
        RECT 5.605 3304.885 6.815 3305.635 ;
        RECT 2910.045 3304.885 2910.335 3305.610 ;
        RECT 2912.805 3304.885 2914.015 3305.635 ;
        RECT 5.520 3304.715 6.900 3304.885 ;
        RECT 2909.960 3304.715 2910.420 3304.885 ;
        RECT 2912.720 3304.715 2914.100 3304.885 ;
        RECT 5.605 3303.965 6.815 3304.715 ;
        RECT 2912.805 3303.965 2914.015 3304.715 ;
        RECT 5.605 3303.425 6.125 3303.965 ;
        RECT 2913.495 3303.425 2914.015 3303.965 ;
        RECT 5.605 3300.195 6.125 3300.735 ;
        RECT 2913.495 3300.195 2914.015 3300.735 ;
        RECT 5.605 3299.445 6.815 3300.195 ;
        RECT 2910.045 3299.445 2910.335 3300.170 ;
        RECT 2912.805 3299.445 2914.015 3300.195 ;
        RECT 5.520 3299.275 6.900 3299.445 ;
        RECT 2909.960 3299.275 2910.420 3299.445 ;
        RECT 2912.720 3299.275 2914.100 3299.445 ;
        RECT 5.605 3298.525 6.815 3299.275 ;
        RECT 2912.805 3298.525 2914.015 3299.275 ;
        RECT 5.605 3297.985 6.125 3298.525 ;
        RECT 2913.495 3297.985 2914.015 3298.525 ;
        RECT 5.605 3294.755 6.125 3295.295 ;
        RECT 2913.495 3294.755 2914.015 3295.295 ;
        RECT 5.605 3294.005 6.815 3294.755 ;
        RECT 2910.045 3294.005 2910.335 3294.730 ;
        RECT 2912.805 3294.005 2914.015 3294.755 ;
        RECT 5.520 3293.835 6.900 3294.005 ;
        RECT 2909.960 3293.835 2910.420 3294.005 ;
        RECT 2912.720 3293.835 2914.100 3294.005 ;
        RECT 5.605 3293.085 6.815 3293.835 ;
        RECT 2912.805 3293.085 2914.015 3293.835 ;
        RECT 5.605 3292.545 6.125 3293.085 ;
        RECT 2913.495 3292.545 2914.015 3293.085 ;
        RECT 5.605 3289.315 6.125 3289.855 ;
        RECT 2913.495 3289.315 2914.015 3289.855 ;
        RECT 5.605 3288.565 6.815 3289.315 ;
        RECT 2910.045 3288.565 2910.335 3289.290 ;
        RECT 2912.805 3288.565 2914.015 3289.315 ;
        RECT 5.520 3288.395 6.900 3288.565 ;
        RECT 2909.960 3288.395 2910.420 3288.565 ;
        RECT 2912.720 3288.395 2914.100 3288.565 ;
        RECT 5.605 3287.645 6.815 3288.395 ;
        RECT 2912.805 3287.645 2914.015 3288.395 ;
        RECT 5.605 3287.105 6.125 3287.645 ;
        RECT 2913.495 3287.105 2914.015 3287.645 ;
        RECT 5.605 3283.875 6.125 3284.415 ;
        RECT 2913.495 3283.875 2914.015 3284.415 ;
        RECT 5.605 3283.125 6.815 3283.875 ;
        RECT 2910.045 3283.125 2910.335 3283.850 ;
        RECT 2912.805 3283.125 2914.015 3283.875 ;
        RECT 5.520 3282.955 6.900 3283.125 ;
        RECT 2909.960 3282.955 2910.420 3283.125 ;
        RECT 2912.720 3282.955 2914.100 3283.125 ;
        RECT 5.605 3282.205 6.815 3282.955 ;
        RECT 2912.805 3282.205 2914.015 3282.955 ;
        RECT 5.605 3281.665 6.125 3282.205 ;
        RECT 2913.495 3281.665 2914.015 3282.205 ;
        RECT 5.605 3278.435 6.125 3278.975 ;
        RECT 2913.495 3278.435 2914.015 3278.975 ;
        RECT 5.605 3277.685 6.815 3278.435 ;
        RECT 2910.045 3277.685 2910.335 3278.410 ;
        RECT 2912.805 3277.685 2914.015 3278.435 ;
        RECT 5.520 3277.515 6.900 3277.685 ;
        RECT 2909.960 3277.515 2910.420 3277.685 ;
        RECT 2912.720 3277.515 2914.100 3277.685 ;
        RECT 5.605 3276.765 6.815 3277.515 ;
        RECT 2912.805 3276.765 2914.015 3277.515 ;
        RECT 5.605 3276.225 6.125 3276.765 ;
        RECT 2913.495 3276.225 2914.015 3276.765 ;
        RECT 5.605 3272.995 6.125 3273.535 ;
        RECT 2913.495 3272.995 2914.015 3273.535 ;
        RECT 5.605 3272.245 6.815 3272.995 ;
        RECT 2910.045 3272.245 2910.335 3272.970 ;
        RECT 2912.805 3272.245 2914.015 3272.995 ;
        RECT 5.520 3272.075 6.900 3272.245 ;
        RECT 2909.960 3272.075 2910.420 3272.245 ;
        RECT 2912.720 3272.075 2914.100 3272.245 ;
        RECT 5.605 3271.325 6.815 3272.075 ;
        RECT 2912.805 3271.325 2914.015 3272.075 ;
        RECT 5.605 3270.785 6.125 3271.325 ;
        RECT 2913.495 3270.785 2914.015 3271.325 ;
        RECT 5.605 3267.555 6.125 3268.095 ;
        RECT 2913.495 3267.555 2914.015 3268.095 ;
        RECT 5.605 3266.805 6.815 3267.555 ;
        RECT 2910.045 3266.805 2910.335 3267.530 ;
        RECT 2912.805 3266.805 2914.015 3267.555 ;
        RECT 5.520 3266.635 6.900 3266.805 ;
        RECT 2909.960 3266.635 2910.420 3266.805 ;
        RECT 2912.720 3266.635 2914.100 3266.805 ;
        RECT 5.605 3265.885 6.815 3266.635 ;
        RECT 2912.805 3265.885 2914.015 3266.635 ;
        RECT 5.605 3265.345 6.125 3265.885 ;
        RECT 2913.495 3265.345 2914.015 3265.885 ;
        RECT 5.605 3262.115 6.125 3262.655 ;
        RECT 2913.495 3262.115 2914.015 3262.655 ;
        RECT 5.605 3261.365 6.815 3262.115 ;
        RECT 2910.045 3261.365 2910.335 3262.090 ;
        RECT 2912.805 3261.365 2914.015 3262.115 ;
        RECT 5.520 3261.195 6.900 3261.365 ;
        RECT 2909.960 3261.195 2910.420 3261.365 ;
        RECT 2912.720 3261.195 2914.100 3261.365 ;
        RECT 5.605 3260.445 6.815 3261.195 ;
        RECT 2912.805 3260.445 2914.015 3261.195 ;
        RECT 5.605 3259.905 6.125 3260.445 ;
        RECT 2913.495 3259.905 2914.015 3260.445 ;
        RECT 5.605 3256.675 6.125 3257.215 ;
        RECT 2913.495 3256.675 2914.015 3257.215 ;
        RECT 5.605 3255.925 6.815 3256.675 ;
        RECT 2910.045 3255.925 2910.335 3256.650 ;
        RECT 2912.805 3255.925 2914.015 3256.675 ;
        RECT 5.520 3255.755 6.900 3255.925 ;
        RECT 2909.960 3255.755 2910.420 3255.925 ;
        RECT 2912.720 3255.755 2914.100 3255.925 ;
        RECT 5.605 3255.005 6.815 3255.755 ;
        RECT 2912.805 3255.005 2914.015 3255.755 ;
        RECT 5.605 3254.465 6.125 3255.005 ;
        RECT 2913.495 3254.465 2914.015 3255.005 ;
        RECT 5.605 3251.235 6.125 3251.775 ;
        RECT 2913.495 3251.235 2914.015 3251.775 ;
        RECT 5.605 3250.485 6.815 3251.235 ;
        RECT 2910.045 3250.485 2910.335 3251.210 ;
        RECT 2912.805 3250.485 2914.015 3251.235 ;
        RECT 5.520 3250.315 6.900 3250.485 ;
        RECT 2909.960 3250.315 2910.420 3250.485 ;
        RECT 2912.720 3250.315 2914.100 3250.485 ;
        RECT 5.605 3249.565 6.815 3250.315 ;
        RECT 2912.805 3249.565 2914.015 3250.315 ;
        RECT 5.605 3249.025 6.125 3249.565 ;
        RECT 2913.495 3249.025 2914.015 3249.565 ;
        RECT 5.605 3245.795 6.125 3246.335 ;
        RECT 2913.495 3245.795 2914.015 3246.335 ;
        RECT 5.605 3245.045 6.815 3245.795 ;
        RECT 2910.045 3245.045 2910.335 3245.770 ;
        RECT 2912.805 3245.045 2914.015 3245.795 ;
        RECT 5.520 3244.875 6.900 3245.045 ;
        RECT 2909.960 3244.875 2910.420 3245.045 ;
        RECT 2912.720 3244.875 2914.100 3245.045 ;
        RECT 5.605 3244.125 6.815 3244.875 ;
        RECT 2912.805 3244.125 2914.015 3244.875 ;
        RECT 5.605 3243.585 6.125 3244.125 ;
        RECT 2913.495 3243.585 2914.015 3244.125 ;
        RECT 5.605 3240.355 6.125 3240.895 ;
        RECT 2913.495 3240.355 2914.015 3240.895 ;
        RECT 5.605 3239.605 6.815 3240.355 ;
        RECT 2910.045 3239.605 2910.335 3240.330 ;
        RECT 2912.805 3239.605 2914.015 3240.355 ;
        RECT 5.520 3239.435 6.900 3239.605 ;
        RECT 2909.960 3239.435 2910.420 3239.605 ;
        RECT 2912.720 3239.435 2914.100 3239.605 ;
        RECT 5.605 3238.685 6.815 3239.435 ;
        RECT 2912.805 3238.685 2914.015 3239.435 ;
        RECT 5.605 3238.145 6.125 3238.685 ;
        RECT 2913.495 3238.145 2914.015 3238.685 ;
        RECT 5.605 3234.915 6.125 3235.455 ;
        RECT 2913.495 3234.915 2914.015 3235.455 ;
        RECT 5.605 3234.165 6.815 3234.915 ;
        RECT 2910.045 3234.165 2910.335 3234.890 ;
        RECT 2912.805 3234.165 2914.015 3234.915 ;
        RECT 5.520 3233.995 6.900 3234.165 ;
        RECT 2909.960 3233.995 2910.420 3234.165 ;
        RECT 2912.720 3233.995 2914.100 3234.165 ;
        RECT 5.605 3233.245 6.815 3233.995 ;
        RECT 2912.805 3233.245 2914.015 3233.995 ;
        RECT 5.605 3232.705 6.125 3233.245 ;
        RECT 2913.495 3232.705 2914.015 3233.245 ;
        RECT 5.605 3229.475 6.125 3230.015 ;
        RECT 2913.495 3229.475 2914.015 3230.015 ;
        RECT 5.605 3228.725 6.815 3229.475 ;
        RECT 2910.045 3228.725 2910.335 3229.450 ;
        RECT 2912.805 3228.725 2914.015 3229.475 ;
        RECT 5.520 3228.555 6.900 3228.725 ;
        RECT 2909.960 3228.555 2910.420 3228.725 ;
        RECT 2912.720 3228.555 2914.100 3228.725 ;
        RECT 5.605 3227.805 6.815 3228.555 ;
        RECT 2912.805 3227.805 2914.015 3228.555 ;
        RECT 5.605 3227.265 6.125 3227.805 ;
        RECT 2913.495 3227.265 2914.015 3227.805 ;
        RECT 5.605 3224.035 6.125 3224.575 ;
        RECT 2913.495 3224.035 2914.015 3224.575 ;
        RECT 5.605 3223.285 6.815 3224.035 ;
        RECT 9.515 3223.285 9.855 3223.945 ;
        RECT 2910.045 3223.285 2910.335 3224.010 ;
        RECT 2912.805 3223.285 2914.015 3224.035 ;
        RECT 5.520 3223.115 6.900 3223.285 ;
        RECT 8.740 3223.115 10.120 3223.285 ;
        RECT 2909.960 3223.115 2910.420 3223.285 ;
        RECT 2912.720 3223.115 2914.100 3223.285 ;
        RECT 5.605 3222.365 6.815 3223.115 ;
        RECT 2912.805 3222.365 2914.015 3223.115 ;
        RECT 5.605 3221.825 6.125 3222.365 ;
        RECT 2913.495 3221.825 2914.015 3222.365 ;
        RECT 5.605 3218.595 6.125 3219.135 ;
        RECT 2913.495 3218.595 2914.015 3219.135 ;
        RECT 5.605 3217.845 6.815 3218.595 ;
        RECT 2910.045 3217.845 2910.335 3218.570 ;
        RECT 2912.805 3217.845 2914.015 3218.595 ;
        RECT 5.520 3217.675 6.900 3217.845 ;
        RECT 2909.960 3217.675 2910.420 3217.845 ;
        RECT 2912.720 3217.675 2914.100 3217.845 ;
        RECT 5.605 3216.925 6.815 3217.675 ;
        RECT 2912.805 3216.925 2914.015 3217.675 ;
        RECT 5.605 3216.385 6.125 3216.925 ;
        RECT 2913.495 3216.385 2914.015 3216.925 ;
        RECT 5.605 3213.155 6.125 3213.695 ;
        RECT 2913.495 3213.155 2914.015 3213.695 ;
        RECT 5.605 3212.405 6.815 3213.155 ;
        RECT 2910.045 3212.405 2910.335 3213.130 ;
        RECT 2912.805 3212.405 2914.015 3213.155 ;
        RECT 5.520 3212.235 6.900 3212.405 ;
        RECT 2909.960 3212.235 2910.420 3212.405 ;
        RECT 2912.720 3212.235 2914.100 3212.405 ;
        RECT 5.605 3211.485 6.815 3212.235 ;
        RECT 2912.805 3211.485 2914.015 3212.235 ;
        RECT 5.605 3210.945 6.125 3211.485 ;
        RECT 2913.495 3210.945 2914.015 3211.485 ;
        RECT 5.605 3207.715 6.125 3208.255 ;
        RECT 2913.495 3207.715 2914.015 3208.255 ;
        RECT 5.605 3206.965 6.815 3207.715 ;
        RECT 2910.045 3206.965 2910.335 3207.690 ;
        RECT 2912.805 3206.965 2914.015 3207.715 ;
        RECT 5.520 3206.795 6.900 3206.965 ;
        RECT 2909.960 3206.795 2910.420 3206.965 ;
        RECT 2912.720 3206.795 2914.100 3206.965 ;
        RECT 5.605 3206.045 6.815 3206.795 ;
        RECT 2912.805 3206.045 2914.015 3206.795 ;
        RECT 5.605 3205.505 6.125 3206.045 ;
        RECT 2913.495 3205.505 2914.015 3206.045 ;
        RECT 5.605 3202.275 6.125 3202.815 ;
        RECT 2913.495 3202.275 2914.015 3202.815 ;
        RECT 5.605 3201.525 6.815 3202.275 ;
        RECT 2910.045 3201.525 2910.335 3202.250 ;
        RECT 2911.195 3201.525 2911.535 3202.185 ;
        RECT 2912.805 3201.525 2914.015 3202.275 ;
        RECT 5.520 3201.355 6.900 3201.525 ;
        RECT 2909.960 3201.355 2911.800 3201.525 ;
        RECT 2912.720 3201.355 2914.100 3201.525 ;
        RECT 5.605 3200.605 6.815 3201.355 ;
        RECT 2912.805 3200.605 2914.015 3201.355 ;
        RECT 5.605 3200.065 6.125 3200.605 ;
        RECT 2913.495 3200.065 2914.015 3200.605 ;
        RECT 5.605 3196.835 6.125 3197.375 ;
        RECT 2913.495 3196.835 2914.015 3197.375 ;
        RECT 5.605 3196.085 6.815 3196.835 ;
        RECT 2910.045 3196.085 2910.335 3196.810 ;
        RECT 2912.805 3196.085 2914.015 3196.835 ;
        RECT 5.520 3195.915 6.900 3196.085 ;
        RECT 2909.960 3195.915 2910.420 3196.085 ;
        RECT 2912.720 3195.915 2914.100 3196.085 ;
        RECT 5.605 3195.165 6.815 3195.915 ;
        RECT 2912.805 3195.165 2914.015 3195.915 ;
        RECT 5.605 3194.625 6.125 3195.165 ;
        RECT 2913.495 3194.625 2914.015 3195.165 ;
        RECT 5.605 3191.395 6.125 3191.935 ;
        RECT 2913.495 3191.395 2914.015 3191.935 ;
        RECT 5.605 3190.645 6.815 3191.395 ;
        RECT 2910.045 3190.645 2910.335 3191.370 ;
        RECT 2912.805 3190.645 2914.015 3191.395 ;
        RECT 5.520 3190.475 6.900 3190.645 ;
        RECT 2909.960 3190.475 2910.420 3190.645 ;
        RECT 2912.720 3190.475 2914.100 3190.645 ;
        RECT 5.605 3189.725 6.815 3190.475 ;
        RECT 2912.805 3189.725 2914.015 3190.475 ;
        RECT 5.605 3189.185 6.125 3189.725 ;
        RECT 2913.495 3189.185 2914.015 3189.725 ;
        RECT 5.605 3185.955 6.125 3186.495 ;
        RECT 2913.495 3185.955 2914.015 3186.495 ;
        RECT 5.605 3185.205 6.815 3185.955 ;
        RECT 2910.045 3185.205 2910.335 3185.930 ;
        RECT 2912.805 3185.205 2914.015 3185.955 ;
        RECT 5.520 3185.035 6.900 3185.205 ;
        RECT 2909.960 3185.035 2910.420 3185.205 ;
        RECT 2912.720 3185.035 2914.100 3185.205 ;
        RECT 5.605 3184.285 6.815 3185.035 ;
        RECT 2912.805 3184.285 2914.015 3185.035 ;
        RECT 5.605 3183.745 6.125 3184.285 ;
        RECT 2913.495 3183.745 2914.015 3184.285 ;
        RECT 5.605 3180.515 6.125 3181.055 ;
        RECT 2913.495 3180.515 2914.015 3181.055 ;
        RECT 5.605 3179.765 6.815 3180.515 ;
        RECT 2910.045 3179.765 2910.335 3180.490 ;
        RECT 2912.805 3179.765 2914.015 3180.515 ;
        RECT 5.520 3179.595 6.900 3179.765 ;
        RECT 2909.960 3179.595 2910.420 3179.765 ;
        RECT 2912.720 3179.595 2914.100 3179.765 ;
        RECT 5.605 3178.845 6.815 3179.595 ;
        RECT 2912.805 3178.845 2914.015 3179.595 ;
        RECT 5.605 3178.305 6.125 3178.845 ;
        RECT 2913.495 3178.305 2914.015 3178.845 ;
        RECT 5.605 3175.075 6.125 3175.615 ;
        RECT 2913.495 3175.075 2914.015 3175.615 ;
        RECT 5.605 3174.325 6.815 3175.075 ;
        RECT 2910.045 3174.325 2910.335 3175.050 ;
        RECT 2912.805 3174.325 2914.015 3175.075 ;
        RECT 5.520 3174.155 6.900 3174.325 ;
        RECT 2909.960 3174.155 2910.420 3174.325 ;
        RECT 2912.720 3174.155 2914.100 3174.325 ;
        RECT 5.605 3173.405 6.815 3174.155 ;
        RECT 2912.805 3173.405 2914.015 3174.155 ;
        RECT 5.605 3172.865 6.125 3173.405 ;
        RECT 2913.495 3172.865 2914.015 3173.405 ;
        RECT 5.605 3169.635 6.125 3170.175 ;
        RECT 2913.495 3169.635 2914.015 3170.175 ;
        RECT 5.605 3168.885 6.815 3169.635 ;
        RECT 2910.045 3168.885 2910.335 3169.610 ;
        RECT 2912.805 3168.885 2914.015 3169.635 ;
        RECT 5.520 3168.715 6.900 3168.885 ;
        RECT 2909.960 3168.715 2910.420 3168.885 ;
        RECT 2912.720 3168.715 2914.100 3168.885 ;
        RECT 5.605 3167.965 6.815 3168.715 ;
        RECT 2912.805 3167.965 2914.015 3168.715 ;
        RECT 5.605 3167.425 6.125 3167.965 ;
        RECT 2913.495 3167.425 2914.015 3167.965 ;
        RECT 5.605 3164.195 6.125 3164.735 ;
        RECT 2913.495 3164.195 2914.015 3164.735 ;
        RECT 5.605 3163.445 6.815 3164.195 ;
        RECT 2910.045 3163.445 2910.335 3164.170 ;
        RECT 2912.805 3163.445 2914.015 3164.195 ;
        RECT 5.520 3163.275 6.900 3163.445 ;
        RECT 2909.960 3163.275 2910.420 3163.445 ;
        RECT 2912.720 3163.275 2914.100 3163.445 ;
        RECT 5.605 3162.525 6.815 3163.275 ;
        RECT 2912.805 3162.525 2914.015 3163.275 ;
        RECT 5.605 3161.985 6.125 3162.525 ;
        RECT 2913.495 3161.985 2914.015 3162.525 ;
        RECT 5.605 3158.755 6.125 3159.295 ;
        RECT 2913.495 3158.755 2914.015 3159.295 ;
        RECT 5.605 3158.005 6.815 3158.755 ;
        RECT 2910.045 3158.005 2910.335 3158.730 ;
        RECT 2912.805 3158.005 2914.015 3158.755 ;
        RECT 5.520 3157.835 6.900 3158.005 ;
        RECT 2909.960 3157.835 2910.420 3158.005 ;
        RECT 2912.720 3157.835 2914.100 3158.005 ;
        RECT 5.605 3157.085 6.815 3157.835 ;
        RECT 2912.805 3157.085 2914.015 3157.835 ;
        RECT 5.605 3156.545 6.125 3157.085 ;
        RECT 2913.495 3156.545 2914.015 3157.085 ;
        RECT 5.605 3153.315 6.125 3153.855 ;
        RECT 2913.495 3153.315 2914.015 3153.855 ;
        RECT 5.605 3152.565 6.815 3153.315 ;
        RECT 2910.045 3152.565 2910.335 3153.290 ;
        RECT 2912.805 3152.565 2914.015 3153.315 ;
        RECT 5.520 3152.395 6.900 3152.565 ;
        RECT 2909.960 3152.395 2910.420 3152.565 ;
        RECT 2912.720 3152.395 2914.100 3152.565 ;
        RECT 5.605 3151.645 6.815 3152.395 ;
        RECT 2912.805 3151.645 2914.015 3152.395 ;
        RECT 5.605 3151.105 6.125 3151.645 ;
        RECT 2913.495 3151.105 2914.015 3151.645 ;
        RECT 5.605 3147.875 6.125 3148.415 ;
        RECT 2913.495 3147.875 2914.015 3148.415 ;
        RECT 5.605 3147.125 6.815 3147.875 ;
        RECT 2910.045 3147.125 2910.335 3147.850 ;
        RECT 2912.805 3147.125 2914.015 3147.875 ;
        RECT 5.520 3146.955 6.900 3147.125 ;
        RECT 2909.960 3146.955 2910.420 3147.125 ;
        RECT 2912.720 3146.955 2914.100 3147.125 ;
        RECT 5.605 3146.205 6.815 3146.955 ;
        RECT 2912.805 3146.205 2914.015 3146.955 ;
        RECT 5.605 3145.665 6.125 3146.205 ;
        RECT 2913.495 3145.665 2914.015 3146.205 ;
        RECT 5.605 3142.435 6.125 3142.975 ;
        RECT 2913.495 3142.435 2914.015 3142.975 ;
        RECT 5.605 3141.685 6.815 3142.435 ;
        RECT 2910.045 3141.685 2910.335 3142.410 ;
        RECT 2912.805 3141.685 2914.015 3142.435 ;
        RECT 5.520 3141.515 6.900 3141.685 ;
        RECT 2909.960 3141.515 2910.420 3141.685 ;
        RECT 2912.720 3141.515 2914.100 3141.685 ;
        RECT 5.605 3140.765 6.815 3141.515 ;
        RECT 2912.805 3140.765 2914.015 3141.515 ;
        RECT 5.605 3140.225 6.125 3140.765 ;
        RECT 2913.495 3140.225 2914.015 3140.765 ;
        RECT 5.605 3136.995 6.125 3137.535 ;
        RECT 2913.495 3136.995 2914.015 3137.535 ;
        RECT 5.605 3136.245 6.815 3136.995 ;
        RECT 2910.045 3136.245 2910.335 3136.970 ;
        RECT 2912.805 3136.245 2914.015 3136.995 ;
        RECT 5.520 3136.075 6.900 3136.245 ;
        RECT 2909.960 3136.075 2910.420 3136.245 ;
        RECT 2912.720 3136.075 2914.100 3136.245 ;
        RECT 5.605 3135.325 6.815 3136.075 ;
        RECT 2912.805 3135.325 2914.015 3136.075 ;
        RECT 5.605 3134.785 6.125 3135.325 ;
        RECT 2913.495 3134.785 2914.015 3135.325 ;
        RECT 5.605 3131.555 6.125 3132.095 ;
        RECT 2913.495 3131.555 2914.015 3132.095 ;
        RECT 5.605 3130.805 6.815 3131.555 ;
        RECT 2910.045 3130.805 2910.335 3131.530 ;
        RECT 2912.805 3130.805 2914.015 3131.555 ;
        RECT 5.520 3130.635 6.900 3130.805 ;
        RECT 2909.960 3130.635 2910.420 3130.805 ;
        RECT 2912.720 3130.635 2914.100 3130.805 ;
        RECT 5.605 3129.885 6.815 3130.635 ;
        RECT 2912.805 3129.885 2914.015 3130.635 ;
        RECT 5.605 3129.345 6.125 3129.885 ;
        RECT 2913.495 3129.345 2914.015 3129.885 ;
        RECT 5.605 3126.115 6.125 3126.655 ;
        RECT 2913.495 3126.115 2914.015 3126.655 ;
        RECT 5.605 3125.365 6.815 3126.115 ;
        RECT 2910.045 3125.365 2910.335 3126.090 ;
        RECT 2912.805 3125.365 2914.015 3126.115 ;
        RECT 5.520 3125.195 6.900 3125.365 ;
        RECT 2909.960 3125.195 2910.420 3125.365 ;
        RECT 2912.720 3125.195 2914.100 3125.365 ;
        RECT 5.605 3124.445 6.815 3125.195 ;
        RECT 2912.805 3124.445 2914.015 3125.195 ;
        RECT 5.605 3123.905 6.125 3124.445 ;
        RECT 2913.495 3123.905 2914.015 3124.445 ;
        RECT 5.605 3120.675 6.125 3121.215 ;
        RECT 2913.495 3120.675 2914.015 3121.215 ;
        RECT 5.605 3119.925 6.815 3120.675 ;
        RECT 2910.045 3119.925 2910.335 3120.650 ;
        RECT 2912.805 3119.925 2914.015 3120.675 ;
        RECT 5.520 3119.755 6.900 3119.925 ;
        RECT 2909.960 3119.755 2910.420 3119.925 ;
        RECT 2912.720 3119.755 2914.100 3119.925 ;
        RECT 5.605 3119.005 6.815 3119.755 ;
        RECT 2912.805 3119.005 2914.015 3119.755 ;
        RECT 5.605 3118.465 6.125 3119.005 ;
        RECT 2913.495 3118.465 2914.015 3119.005 ;
        RECT 5.605 3115.235 6.125 3115.775 ;
        RECT 2913.495 3115.235 2914.015 3115.775 ;
        RECT 5.605 3114.485 6.815 3115.235 ;
        RECT 2910.045 3114.485 2910.335 3115.210 ;
        RECT 2912.805 3114.485 2914.015 3115.235 ;
        RECT 5.520 3114.315 6.900 3114.485 ;
        RECT 2909.960 3114.315 2910.420 3114.485 ;
        RECT 2912.720 3114.315 2914.100 3114.485 ;
        RECT 5.605 3113.565 6.815 3114.315 ;
        RECT 2912.805 3113.565 2914.015 3114.315 ;
        RECT 5.605 3113.025 6.125 3113.565 ;
        RECT 2913.495 3113.025 2914.015 3113.565 ;
        RECT 5.605 3109.795 6.125 3110.335 ;
        RECT 2913.495 3109.795 2914.015 3110.335 ;
        RECT 5.605 3109.045 6.815 3109.795 ;
        RECT 2910.045 3109.045 2910.335 3109.770 ;
        RECT 2912.805 3109.045 2914.015 3109.795 ;
        RECT 5.520 3108.875 6.900 3109.045 ;
        RECT 2909.960 3108.875 2910.420 3109.045 ;
        RECT 2912.720 3108.875 2914.100 3109.045 ;
        RECT 5.605 3108.125 6.815 3108.875 ;
        RECT 2912.805 3108.125 2914.015 3108.875 ;
        RECT 5.605 3107.585 6.125 3108.125 ;
        RECT 2913.495 3107.585 2914.015 3108.125 ;
        RECT 5.605 3104.355 6.125 3104.895 ;
        RECT 2913.495 3104.355 2914.015 3104.895 ;
        RECT 5.605 3103.605 6.815 3104.355 ;
        RECT 2910.045 3103.605 2910.335 3104.330 ;
        RECT 2912.805 3103.605 2914.015 3104.355 ;
        RECT 5.520 3103.435 6.900 3103.605 ;
        RECT 2909.960 3103.435 2910.420 3103.605 ;
        RECT 2912.720 3103.435 2914.100 3103.605 ;
        RECT 5.605 3102.685 6.815 3103.435 ;
        RECT 2912.805 3102.685 2914.015 3103.435 ;
        RECT 5.605 3102.145 6.125 3102.685 ;
        RECT 2913.495 3102.145 2914.015 3102.685 ;
        RECT 5.605 3098.915 6.125 3099.455 ;
        RECT 2913.495 3098.915 2914.015 3099.455 ;
        RECT 5.605 3098.165 6.815 3098.915 ;
        RECT 2910.045 3098.165 2910.335 3098.890 ;
        RECT 2912.805 3098.165 2914.015 3098.915 ;
        RECT 5.520 3097.995 6.900 3098.165 ;
        RECT 2909.040 3097.995 2910.420 3098.165 ;
        RECT 2912.720 3097.995 2914.100 3098.165 ;
        RECT 5.605 3097.245 6.815 3097.995 ;
        RECT 2909.815 3097.335 2910.155 3097.995 ;
        RECT 2912.805 3097.245 2914.015 3097.995 ;
        RECT 5.605 3096.705 6.125 3097.245 ;
        RECT 2913.495 3096.705 2914.015 3097.245 ;
        RECT 5.605 3093.475 6.125 3094.015 ;
        RECT 2913.495 3093.475 2914.015 3094.015 ;
        RECT 5.605 3092.725 6.815 3093.475 ;
        RECT 2910.045 3092.725 2910.335 3093.450 ;
        RECT 2912.805 3092.725 2914.015 3093.475 ;
        RECT 5.520 3092.555 6.900 3092.725 ;
        RECT 2909.960 3092.555 2910.420 3092.725 ;
        RECT 2912.720 3092.555 2914.100 3092.725 ;
        RECT 5.605 3091.805 6.815 3092.555 ;
        RECT 2912.805 3091.805 2914.015 3092.555 ;
        RECT 5.605 3091.265 6.125 3091.805 ;
        RECT 2913.495 3091.265 2914.015 3091.805 ;
        RECT 5.605 3088.035 6.125 3088.575 ;
        RECT 2913.495 3088.035 2914.015 3088.575 ;
        RECT 5.605 3087.285 6.815 3088.035 ;
        RECT 2910.045 3087.285 2910.335 3088.010 ;
        RECT 2912.805 3087.285 2914.015 3088.035 ;
        RECT 5.520 3087.115 6.900 3087.285 ;
        RECT 2909.960 3087.115 2910.420 3087.285 ;
        RECT 2912.720 3087.115 2914.100 3087.285 ;
        RECT 5.605 3086.365 6.815 3087.115 ;
        RECT 2912.805 3086.365 2914.015 3087.115 ;
        RECT 5.605 3085.825 6.125 3086.365 ;
        RECT 2913.495 3085.825 2914.015 3086.365 ;
        RECT 5.605 3082.595 6.125 3083.135 ;
        RECT 2913.495 3082.595 2914.015 3083.135 ;
        RECT 5.605 3081.845 6.815 3082.595 ;
        RECT 2910.045 3081.845 2910.335 3082.570 ;
        RECT 2912.805 3081.845 2914.015 3082.595 ;
        RECT 5.520 3081.675 6.900 3081.845 ;
        RECT 2909.960 3081.675 2910.420 3081.845 ;
        RECT 2912.720 3081.675 2914.100 3081.845 ;
        RECT 5.605 3080.925 6.815 3081.675 ;
        RECT 2912.805 3080.925 2914.015 3081.675 ;
        RECT 5.605 3080.385 6.125 3080.925 ;
        RECT 2913.495 3080.385 2914.015 3080.925 ;
        RECT 5.605 3077.155 6.125 3077.695 ;
        RECT 2913.495 3077.155 2914.015 3077.695 ;
        RECT 5.605 3076.405 6.815 3077.155 ;
        RECT 2910.045 3076.405 2910.335 3077.130 ;
        RECT 2912.805 3076.405 2914.015 3077.155 ;
        RECT 5.520 3076.235 6.900 3076.405 ;
        RECT 2909.960 3076.235 2910.420 3076.405 ;
        RECT 2912.720 3076.235 2914.100 3076.405 ;
        RECT 5.605 3075.485 6.815 3076.235 ;
        RECT 2912.805 3075.485 2914.015 3076.235 ;
        RECT 5.605 3074.945 6.125 3075.485 ;
        RECT 2913.495 3074.945 2914.015 3075.485 ;
        RECT 5.605 3071.715 6.125 3072.255 ;
        RECT 2913.495 3071.715 2914.015 3072.255 ;
        RECT 5.605 3070.965 6.815 3071.715 ;
        RECT 2910.045 3070.965 2910.335 3071.690 ;
        RECT 2912.805 3070.965 2914.015 3071.715 ;
        RECT 5.520 3070.795 6.900 3070.965 ;
        RECT 2909.960 3070.795 2910.420 3070.965 ;
        RECT 2912.720 3070.795 2914.100 3070.965 ;
        RECT 5.605 3070.045 6.815 3070.795 ;
        RECT 2912.805 3070.045 2914.015 3070.795 ;
        RECT 5.605 3069.505 6.125 3070.045 ;
        RECT 2913.495 3069.505 2914.015 3070.045 ;
        RECT 5.605 3066.275 6.125 3066.815 ;
        RECT 2913.495 3066.275 2914.015 3066.815 ;
        RECT 5.605 3065.525 6.815 3066.275 ;
        RECT 2910.045 3065.525 2910.335 3066.250 ;
        RECT 2912.805 3065.525 2914.015 3066.275 ;
        RECT 5.520 3065.355 6.900 3065.525 ;
        RECT 2909.960 3065.355 2910.420 3065.525 ;
        RECT 2912.720 3065.355 2914.100 3065.525 ;
        RECT 5.605 3064.605 6.815 3065.355 ;
        RECT 2912.805 3064.605 2914.015 3065.355 ;
        RECT 5.605 3064.065 6.125 3064.605 ;
        RECT 2913.495 3064.065 2914.015 3064.605 ;
        RECT 5.605 3060.835 6.125 3061.375 ;
        RECT 2913.495 3060.835 2914.015 3061.375 ;
        RECT 5.605 3060.085 6.815 3060.835 ;
        RECT 2910.045 3060.085 2910.335 3060.810 ;
        RECT 2912.805 3060.085 2914.015 3060.835 ;
        RECT 5.520 3059.915 6.900 3060.085 ;
        RECT 2909.960 3059.915 2910.420 3060.085 ;
        RECT 2912.720 3059.915 2914.100 3060.085 ;
        RECT 5.605 3059.165 6.815 3059.915 ;
        RECT 2912.805 3059.165 2914.015 3059.915 ;
        RECT 5.605 3058.625 6.125 3059.165 ;
        RECT 2913.495 3058.625 2914.015 3059.165 ;
        RECT 5.605 3055.395 6.125 3055.935 ;
        RECT 2913.495 3055.395 2914.015 3055.935 ;
        RECT 5.605 3054.645 6.815 3055.395 ;
        RECT 2910.045 3054.645 2910.335 3055.370 ;
        RECT 2912.805 3054.645 2914.015 3055.395 ;
        RECT 5.520 3054.475 6.900 3054.645 ;
        RECT 2909.960 3054.475 2910.420 3054.645 ;
        RECT 2912.720 3054.475 2914.100 3054.645 ;
        RECT 5.605 3053.725 6.815 3054.475 ;
        RECT 2912.805 3053.725 2914.015 3054.475 ;
        RECT 5.605 3053.185 6.125 3053.725 ;
        RECT 2913.495 3053.185 2914.015 3053.725 ;
        RECT 5.605 3049.955 6.125 3050.495 ;
        RECT 2913.495 3049.955 2914.015 3050.495 ;
        RECT 5.605 3049.205 6.815 3049.955 ;
        RECT 2910.045 3049.205 2910.335 3049.930 ;
        RECT 2912.805 3049.205 2914.015 3049.955 ;
        RECT 5.520 3049.035 6.900 3049.205 ;
        RECT 2909.960 3049.035 2910.420 3049.205 ;
        RECT 2912.720 3049.035 2914.100 3049.205 ;
        RECT 5.605 3048.285 6.815 3049.035 ;
        RECT 2912.805 3048.285 2914.015 3049.035 ;
        RECT 5.605 3047.745 6.125 3048.285 ;
        RECT 2913.495 3047.745 2914.015 3048.285 ;
        RECT 5.605 3044.515 6.125 3045.055 ;
        RECT 2913.495 3044.515 2914.015 3045.055 ;
        RECT 5.605 3043.765 6.815 3044.515 ;
        RECT 2910.045 3043.765 2910.335 3044.490 ;
        RECT 2912.805 3043.765 2914.015 3044.515 ;
        RECT 5.520 3043.595 6.900 3043.765 ;
        RECT 2909.960 3043.595 2910.420 3043.765 ;
        RECT 2912.720 3043.595 2914.100 3043.765 ;
        RECT 5.605 3042.845 6.815 3043.595 ;
        RECT 2912.805 3042.845 2914.015 3043.595 ;
        RECT 5.605 3042.305 6.125 3042.845 ;
        RECT 2913.495 3042.305 2914.015 3042.845 ;
        RECT 5.605 3039.075 6.125 3039.615 ;
        RECT 2913.495 3039.075 2914.015 3039.615 ;
        RECT 5.605 3038.325 6.815 3039.075 ;
        RECT 2910.045 3038.325 2910.335 3039.050 ;
        RECT 2912.805 3038.325 2914.015 3039.075 ;
        RECT 5.520 3038.155 6.900 3038.325 ;
        RECT 2909.960 3038.155 2910.420 3038.325 ;
        RECT 2912.720 3038.155 2914.100 3038.325 ;
        RECT 5.605 3037.405 6.815 3038.155 ;
        RECT 2912.805 3037.405 2914.015 3038.155 ;
        RECT 5.605 3036.865 6.125 3037.405 ;
        RECT 2913.495 3036.865 2914.015 3037.405 ;
        RECT 5.605 3033.635 6.125 3034.175 ;
        RECT 2913.495 3033.635 2914.015 3034.175 ;
        RECT 5.605 3032.885 6.815 3033.635 ;
        RECT 2910.045 3032.885 2910.335 3033.610 ;
        RECT 2912.805 3032.885 2914.015 3033.635 ;
        RECT 5.520 3032.715 6.900 3032.885 ;
        RECT 2909.960 3032.715 2910.420 3032.885 ;
        RECT 2912.720 3032.715 2914.100 3032.885 ;
        RECT 5.605 3031.965 6.815 3032.715 ;
        RECT 2912.805 3031.965 2914.015 3032.715 ;
        RECT 5.605 3031.425 6.125 3031.965 ;
        RECT 2913.495 3031.425 2914.015 3031.965 ;
        RECT 5.605 3028.195 6.125 3028.735 ;
        RECT 2913.495 3028.195 2914.015 3028.735 ;
        RECT 5.605 3027.445 6.815 3028.195 ;
        RECT 2910.045 3027.445 2910.335 3028.170 ;
        RECT 2912.805 3027.445 2914.015 3028.195 ;
        RECT 5.520 3027.275 6.900 3027.445 ;
        RECT 2909.960 3027.275 2910.420 3027.445 ;
        RECT 2912.720 3027.275 2914.100 3027.445 ;
        RECT 5.605 3026.525 6.815 3027.275 ;
        RECT 2912.805 3026.525 2914.015 3027.275 ;
        RECT 5.605 3025.985 6.125 3026.525 ;
        RECT 2913.495 3025.985 2914.015 3026.525 ;
        RECT 5.605 3022.755 6.125 3023.295 ;
        RECT 2913.495 3022.755 2914.015 3023.295 ;
        RECT 5.605 3022.005 6.815 3022.755 ;
        RECT 2910.045 3022.005 2910.335 3022.730 ;
        RECT 2912.805 3022.005 2914.015 3022.755 ;
        RECT 5.520 3021.835 6.900 3022.005 ;
        RECT 2909.960 3021.835 2910.420 3022.005 ;
        RECT 2912.720 3021.835 2914.100 3022.005 ;
        RECT 5.605 3021.085 6.815 3021.835 ;
        RECT 2912.805 3021.085 2914.015 3021.835 ;
        RECT 5.605 3020.545 6.125 3021.085 ;
        RECT 2913.495 3020.545 2914.015 3021.085 ;
        RECT 5.605 3017.315 6.125 3017.855 ;
        RECT 2913.495 3017.315 2914.015 3017.855 ;
        RECT 5.605 3016.565 6.815 3017.315 ;
        RECT 2910.045 3016.565 2910.335 3017.290 ;
        RECT 2912.805 3016.565 2914.015 3017.315 ;
        RECT 5.520 3016.395 6.900 3016.565 ;
        RECT 2909.960 3016.395 2910.420 3016.565 ;
        RECT 2912.720 3016.395 2914.100 3016.565 ;
        RECT 5.605 3015.645 6.815 3016.395 ;
        RECT 2912.805 3015.645 2914.015 3016.395 ;
        RECT 5.605 3015.105 6.125 3015.645 ;
        RECT 2913.495 3015.105 2914.015 3015.645 ;
        RECT 5.605 3011.875 6.125 3012.415 ;
        RECT 2913.495 3011.875 2914.015 3012.415 ;
        RECT 5.605 3011.125 6.815 3011.875 ;
        RECT 9.515 3011.125 9.855 3011.785 ;
        RECT 2910.045 3011.125 2910.335 3011.850 ;
        RECT 2912.805 3011.125 2914.015 3011.875 ;
        RECT 5.520 3010.955 6.900 3011.125 ;
        RECT 8.740 3010.955 10.120 3011.125 ;
        RECT 2909.960 3010.955 2910.420 3011.125 ;
        RECT 2912.720 3010.955 2914.100 3011.125 ;
        RECT 5.605 3010.205 6.815 3010.955 ;
        RECT 2912.805 3010.205 2914.015 3010.955 ;
        RECT 5.605 3009.665 6.125 3010.205 ;
        RECT 2913.495 3009.665 2914.015 3010.205 ;
        RECT 5.605 3006.435 6.125 3006.975 ;
        RECT 2913.495 3006.435 2914.015 3006.975 ;
        RECT 5.605 3005.685 6.815 3006.435 ;
        RECT 2910.045 3005.685 2910.335 3006.410 ;
        RECT 2912.805 3005.685 2914.015 3006.435 ;
        RECT 5.520 3005.515 6.900 3005.685 ;
        RECT 2909.960 3005.515 2910.420 3005.685 ;
        RECT 2912.720 3005.515 2914.100 3005.685 ;
        RECT 5.605 3004.765 6.815 3005.515 ;
        RECT 2912.805 3004.765 2914.015 3005.515 ;
        RECT 5.605 3004.225 6.125 3004.765 ;
        RECT 2913.495 3004.225 2914.015 3004.765 ;
        RECT 5.605 3000.995 6.125 3001.535 ;
        RECT 2913.495 3000.995 2914.015 3001.535 ;
        RECT 5.605 3000.245 6.815 3000.995 ;
        RECT 2910.045 3000.245 2910.335 3000.970 ;
        RECT 2912.805 3000.245 2914.015 3000.995 ;
        RECT 5.520 3000.075 6.900 3000.245 ;
        RECT 2909.960 3000.075 2910.420 3000.245 ;
        RECT 2912.720 3000.075 2914.100 3000.245 ;
        RECT 5.605 2999.325 6.815 3000.075 ;
        RECT 2912.805 2999.325 2914.015 3000.075 ;
        RECT 5.605 2998.785 6.125 2999.325 ;
        RECT 2913.495 2998.785 2914.015 2999.325 ;
        RECT 5.605 2995.555 6.125 2996.095 ;
        RECT 2913.495 2995.555 2914.015 2996.095 ;
        RECT 5.605 2994.805 6.815 2995.555 ;
        RECT 2910.045 2994.805 2910.335 2995.530 ;
        RECT 2912.805 2994.805 2914.015 2995.555 ;
        RECT 5.520 2994.635 6.900 2994.805 ;
        RECT 2909.960 2994.635 2910.420 2994.805 ;
        RECT 2912.720 2994.635 2914.100 2994.805 ;
        RECT 5.605 2993.885 6.815 2994.635 ;
        RECT 2912.805 2993.885 2914.015 2994.635 ;
        RECT 5.605 2993.345 6.125 2993.885 ;
        RECT 2913.495 2993.345 2914.015 2993.885 ;
        RECT 5.605 2990.115 6.125 2990.655 ;
        RECT 2913.495 2990.115 2914.015 2990.655 ;
        RECT 5.605 2989.365 6.815 2990.115 ;
        RECT 2910.045 2989.365 2910.335 2990.090 ;
        RECT 2912.805 2989.365 2914.015 2990.115 ;
        RECT 5.520 2989.195 6.900 2989.365 ;
        RECT 2909.960 2989.195 2910.420 2989.365 ;
        RECT 2912.720 2989.195 2914.100 2989.365 ;
        RECT 5.605 2988.445 6.815 2989.195 ;
        RECT 2912.805 2988.445 2914.015 2989.195 ;
        RECT 5.605 2987.905 6.125 2988.445 ;
        RECT 2913.495 2987.905 2914.015 2988.445 ;
        RECT 5.605 2984.675 6.125 2985.215 ;
        RECT 2913.495 2984.675 2914.015 2985.215 ;
        RECT 5.605 2983.925 6.815 2984.675 ;
        RECT 2910.045 2983.925 2910.335 2984.650 ;
        RECT 2912.805 2983.925 2914.015 2984.675 ;
        RECT 5.520 2983.755 6.900 2983.925 ;
        RECT 2909.960 2983.755 2910.420 2983.925 ;
        RECT 2912.720 2983.755 2914.100 2983.925 ;
        RECT 5.605 2983.005 6.815 2983.755 ;
        RECT 2912.805 2983.005 2914.015 2983.755 ;
        RECT 5.605 2982.465 6.125 2983.005 ;
        RECT 2913.495 2982.465 2914.015 2983.005 ;
        RECT 5.605 2979.235 6.125 2979.775 ;
        RECT 2913.495 2979.235 2914.015 2979.775 ;
        RECT 5.605 2978.485 6.815 2979.235 ;
        RECT 2910.045 2978.485 2910.335 2979.210 ;
        RECT 2912.805 2978.485 2914.015 2979.235 ;
        RECT 5.520 2978.315 6.900 2978.485 ;
        RECT 2909.960 2978.315 2910.420 2978.485 ;
        RECT 2912.720 2978.315 2914.100 2978.485 ;
        RECT 5.605 2977.565 6.815 2978.315 ;
        RECT 2912.805 2977.565 2914.015 2978.315 ;
        RECT 5.605 2977.025 6.125 2977.565 ;
        RECT 2913.495 2977.025 2914.015 2977.565 ;
        RECT 5.605 2973.795 6.125 2974.335 ;
        RECT 2913.495 2973.795 2914.015 2974.335 ;
        RECT 5.605 2973.045 6.815 2973.795 ;
        RECT 2910.045 2973.045 2910.335 2973.770 ;
        RECT 2912.805 2973.045 2914.015 2973.795 ;
        RECT 5.520 2972.875 6.900 2973.045 ;
        RECT 8.740 2972.875 10.120 2973.045 ;
        RECT 2909.960 2972.875 2910.420 2973.045 ;
        RECT 2912.720 2972.875 2914.100 2973.045 ;
        RECT 5.605 2972.125 6.815 2972.875 ;
        RECT 9.515 2972.215 9.855 2972.875 ;
        RECT 2912.805 2972.125 2914.015 2972.875 ;
        RECT 5.605 2971.585 6.125 2972.125 ;
        RECT 2913.495 2971.585 2914.015 2972.125 ;
        RECT 5.605 2968.355 6.125 2968.895 ;
        RECT 2913.495 2968.355 2914.015 2968.895 ;
        RECT 5.605 2967.605 6.815 2968.355 ;
        RECT 2910.045 2967.605 2910.335 2968.330 ;
        RECT 2912.805 2967.605 2914.015 2968.355 ;
        RECT 5.520 2967.435 6.900 2967.605 ;
        RECT 2909.960 2967.435 2910.420 2967.605 ;
        RECT 2912.720 2967.435 2914.100 2967.605 ;
        RECT 5.605 2966.685 6.815 2967.435 ;
        RECT 2912.805 2966.685 2914.015 2967.435 ;
        RECT 5.605 2966.145 6.125 2966.685 ;
        RECT 2913.495 2966.145 2914.015 2966.685 ;
        RECT 5.605 2962.915 6.125 2963.455 ;
        RECT 2913.495 2962.915 2914.015 2963.455 ;
        RECT 5.605 2962.165 6.815 2962.915 ;
        RECT 2910.045 2962.165 2910.335 2962.890 ;
        RECT 2912.805 2962.165 2914.015 2962.915 ;
        RECT 5.520 2961.995 6.900 2962.165 ;
        RECT 2909.960 2961.995 2910.420 2962.165 ;
        RECT 2912.720 2961.995 2914.100 2962.165 ;
        RECT 5.605 2961.245 6.815 2961.995 ;
        RECT 2912.805 2961.245 2914.015 2961.995 ;
        RECT 5.605 2960.705 6.125 2961.245 ;
        RECT 2913.495 2960.705 2914.015 2961.245 ;
        RECT 5.605 2957.475 6.125 2958.015 ;
        RECT 2913.495 2957.475 2914.015 2958.015 ;
        RECT 5.605 2956.725 6.815 2957.475 ;
        RECT 2910.045 2956.725 2910.335 2957.450 ;
        RECT 2912.805 2956.725 2914.015 2957.475 ;
        RECT 5.520 2956.555 6.900 2956.725 ;
        RECT 8.740 2956.555 10.120 2956.725 ;
        RECT 2909.960 2956.555 2910.420 2956.725 ;
        RECT 2912.720 2956.555 2914.100 2956.725 ;
        RECT 5.605 2955.805 6.815 2956.555 ;
        RECT 9.515 2955.895 9.855 2956.555 ;
        RECT 2912.805 2955.805 2914.015 2956.555 ;
        RECT 5.605 2955.265 6.125 2955.805 ;
        RECT 2913.495 2955.265 2914.015 2955.805 ;
        RECT 5.605 2952.035 6.125 2952.575 ;
        RECT 2913.495 2952.035 2914.015 2952.575 ;
        RECT 5.605 2951.285 6.815 2952.035 ;
        RECT 2910.045 2951.285 2910.335 2952.010 ;
        RECT 2912.805 2951.285 2914.015 2952.035 ;
        RECT 5.520 2951.115 6.900 2951.285 ;
        RECT 2909.960 2951.115 2910.420 2951.285 ;
        RECT 2912.720 2951.115 2914.100 2951.285 ;
        RECT 5.605 2950.365 6.815 2951.115 ;
        RECT 2912.805 2950.365 2914.015 2951.115 ;
        RECT 5.605 2949.825 6.125 2950.365 ;
        RECT 2913.495 2949.825 2914.015 2950.365 ;
        RECT 5.605 2946.595 6.125 2947.135 ;
        RECT 2913.495 2946.595 2914.015 2947.135 ;
        RECT 5.605 2945.845 6.815 2946.595 ;
        RECT 2910.045 2945.845 2910.335 2946.570 ;
        RECT 2912.805 2945.845 2914.015 2946.595 ;
        RECT 5.520 2945.675 6.900 2945.845 ;
        RECT 2909.960 2945.675 2910.420 2945.845 ;
        RECT 2912.720 2945.675 2914.100 2945.845 ;
        RECT 5.605 2944.925 6.815 2945.675 ;
        RECT 2912.805 2944.925 2914.015 2945.675 ;
        RECT 5.605 2944.385 6.125 2944.925 ;
        RECT 2913.495 2944.385 2914.015 2944.925 ;
        RECT 5.605 2941.155 6.125 2941.695 ;
        RECT 2913.495 2941.155 2914.015 2941.695 ;
        RECT 5.605 2940.405 6.815 2941.155 ;
        RECT 2910.045 2940.405 2910.335 2941.130 ;
        RECT 2912.805 2940.405 2914.015 2941.155 ;
        RECT 5.520 2940.235 6.900 2940.405 ;
        RECT 2909.960 2940.235 2910.420 2940.405 ;
        RECT 2912.720 2940.235 2914.100 2940.405 ;
        RECT 5.605 2939.485 6.815 2940.235 ;
        RECT 2912.805 2939.485 2914.015 2940.235 ;
        RECT 5.605 2938.945 6.125 2939.485 ;
        RECT 2913.495 2938.945 2914.015 2939.485 ;
        RECT 5.605 2935.715 6.125 2936.255 ;
        RECT 2913.495 2935.715 2914.015 2936.255 ;
        RECT 5.605 2934.965 6.815 2935.715 ;
        RECT 2910.045 2934.965 2910.335 2935.690 ;
        RECT 2912.805 2934.965 2914.015 2935.715 ;
        RECT 5.520 2934.795 6.900 2934.965 ;
        RECT 2909.960 2934.795 2910.420 2934.965 ;
        RECT 2912.720 2934.795 2914.100 2934.965 ;
        RECT 5.605 2934.045 6.815 2934.795 ;
        RECT 2912.805 2934.045 2914.015 2934.795 ;
        RECT 5.605 2933.505 6.125 2934.045 ;
        RECT 2913.495 2933.505 2914.015 2934.045 ;
        RECT 5.605 2930.275 6.125 2930.815 ;
        RECT 2913.495 2930.275 2914.015 2930.815 ;
        RECT 5.605 2929.525 6.815 2930.275 ;
        RECT 2910.045 2929.525 2910.335 2930.250 ;
        RECT 2912.805 2929.525 2914.015 2930.275 ;
        RECT 5.520 2929.355 6.900 2929.525 ;
        RECT 2909.960 2929.355 2910.420 2929.525 ;
        RECT 2912.720 2929.355 2914.100 2929.525 ;
        RECT 5.605 2928.605 6.815 2929.355 ;
        RECT 2912.805 2928.605 2914.015 2929.355 ;
        RECT 5.605 2928.065 6.125 2928.605 ;
        RECT 2913.495 2928.065 2914.015 2928.605 ;
        RECT 5.605 2924.835 6.125 2925.375 ;
        RECT 2913.495 2924.835 2914.015 2925.375 ;
        RECT 5.605 2924.085 6.815 2924.835 ;
        RECT 2910.045 2924.085 2910.335 2924.810 ;
        RECT 2912.805 2924.085 2914.015 2924.835 ;
        RECT 5.520 2923.915 6.900 2924.085 ;
        RECT 2909.960 2923.915 2910.420 2924.085 ;
        RECT 2912.720 2923.915 2914.100 2924.085 ;
        RECT 5.605 2923.165 6.815 2923.915 ;
        RECT 2912.805 2923.165 2914.015 2923.915 ;
        RECT 5.605 2922.625 6.125 2923.165 ;
        RECT 2913.495 2922.625 2914.015 2923.165 ;
        RECT 5.605 2919.395 6.125 2919.935 ;
        RECT 2913.495 2919.395 2914.015 2919.935 ;
        RECT 5.605 2918.645 6.815 2919.395 ;
        RECT 2910.045 2918.645 2910.335 2919.370 ;
        RECT 2912.805 2918.645 2914.015 2919.395 ;
        RECT 5.520 2918.475 6.900 2918.645 ;
        RECT 2909.960 2918.475 2910.420 2918.645 ;
        RECT 2912.720 2918.475 2914.100 2918.645 ;
        RECT 5.605 2917.725 6.815 2918.475 ;
        RECT 2912.805 2917.725 2914.015 2918.475 ;
        RECT 5.605 2917.185 6.125 2917.725 ;
        RECT 2913.495 2917.185 2914.015 2917.725 ;
        RECT 5.605 2913.955 6.125 2914.495 ;
        RECT 2913.495 2913.955 2914.015 2914.495 ;
        RECT 5.605 2913.205 6.815 2913.955 ;
        RECT 2910.045 2913.205 2910.335 2913.930 ;
        RECT 2911.195 2913.205 2911.535 2913.865 ;
        RECT 2912.805 2913.205 2914.015 2913.955 ;
        RECT 5.520 2913.035 6.900 2913.205 ;
        RECT 2909.960 2913.035 2911.800 2913.205 ;
        RECT 2912.720 2913.035 2914.100 2913.205 ;
        RECT 5.605 2912.285 6.815 2913.035 ;
        RECT 2912.805 2912.285 2914.015 2913.035 ;
        RECT 5.605 2911.745 6.125 2912.285 ;
        RECT 2913.495 2911.745 2914.015 2912.285 ;
        RECT 5.605 2908.515 6.125 2909.055 ;
        RECT 2913.495 2908.515 2914.015 2909.055 ;
        RECT 5.605 2907.765 6.815 2908.515 ;
        RECT 2910.045 2907.765 2910.335 2908.490 ;
        RECT 2912.805 2907.765 2914.015 2908.515 ;
        RECT 5.520 2907.595 6.900 2907.765 ;
        RECT 2909.960 2907.595 2910.420 2907.765 ;
        RECT 2912.720 2907.595 2914.100 2907.765 ;
        RECT 5.605 2906.845 6.815 2907.595 ;
        RECT 2912.805 2906.845 2914.015 2907.595 ;
        RECT 5.605 2906.305 6.125 2906.845 ;
        RECT 2913.495 2906.305 2914.015 2906.845 ;
        RECT 5.605 2903.075 6.125 2903.615 ;
        RECT 2913.495 2903.075 2914.015 2903.615 ;
        RECT 5.605 2902.325 6.815 2903.075 ;
        RECT 2910.045 2902.325 2910.335 2903.050 ;
        RECT 2912.805 2902.325 2914.015 2903.075 ;
        RECT 5.520 2902.155 6.900 2902.325 ;
        RECT 2909.960 2902.155 2910.420 2902.325 ;
        RECT 2912.720 2902.155 2914.100 2902.325 ;
        RECT 5.605 2901.405 6.815 2902.155 ;
        RECT 2912.805 2901.405 2914.015 2902.155 ;
        RECT 5.605 2900.865 6.125 2901.405 ;
        RECT 2913.495 2900.865 2914.015 2901.405 ;
        RECT 5.605 2897.635 6.125 2898.175 ;
        RECT 2913.495 2897.635 2914.015 2898.175 ;
        RECT 5.605 2896.885 6.815 2897.635 ;
        RECT 2910.045 2896.885 2910.335 2897.610 ;
        RECT 2912.805 2896.885 2914.015 2897.635 ;
        RECT 5.520 2896.715 6.900 2896.885 ;
        RECT 2909.960 2896.715 2910.420 2896.885 ;
        RECT 2912.720 2896.715 2914.100 2896.885 ;
        RECT 5.605 2895.965 6.815 2896.715 ;
        RECT 2912.805 2895.965 2914.015 2896.715 ;
        RECT 5.605 2895.425 6.125 2895.965 ;
        RECT 2913.495 2895.425 2914.015 2895.965 ;
        RECT 5.605 2892.195 6.125 2892.735 ;
        RECT 2913.495 2892.195 2914.015 2892.735 ;
        RECT 5.605 2891.445 6.815 2892.195 ;
        RECT 2910.045 2891.445 2910.335 2892.170 ;
        RECT 2912.805 2891.445 2914.015 2892.195 ;
        RECT 5.520 2891.275 6.900 2891.445 ;
        RECT 2909.960 2891.275 2910.420 2891.445 ;
        RECT 2912.720 2891.275 2914.100 2891.445 ;
        RECT 5.605 2890.525 6.815 2891.275 ;
        RECT 2912.805 2890.525 2914.015 2891.275 ;
        RECT 5.605 2889.985 6.125 2890.525 ;
        RECT 2913.495 2889.985 2914.015 2890.525 ;
        RECT 5.605 2886.755 6.125 2887.295 ;
        RECT 2913.495 2886.755 2914.015 2887.295 ;
        RECT 5.605 2886.005 6.815 2886.755 ;
        RECT 2910.045 2886.005 2910.335 2886.730 ;
        RECT 2912.805 2886.005 2914.015 2886.755 ;
        RECT 5.520 2885.835 6.900 2886.005 ;
        RECT 8.740 2885.835 10.120 2886.005 ;
        RECT 2909.960 2885.835 2910.420 2886.005 ;
        RECT 2912.720 2885.835 2914.100 2886.005 ;
        RECT 5.605 2885.085 6.815 2885.835 ;
        RECT 9.515 2885.175 9.855 2885.835 ;
        RECT 2912.805 2885.085 2914.015 2885.835 ;
        RECT 5.605 2884.545 6.125 2885.085 ;
        RECT 2913.495 2884.545 2914.015 2885.085 ;
        RECT 5.605 2881.315 6.125 2881.855 ;
        RECT 2913.495 2881.315 2914.015 2881.855 ;
        RECT 5.605 2880.565 6.815 2881.315 ;
        RECT 2910.045 2880.565 2910.335 2881.290 ;
        RECT 2912.805 2880.565 2914.015 2881.315 ;
        RECT 5.520 2880.395 6.900 2880.565 ;
        RECT 2909.960 2880.395 2910.420 2880.565 ;
        RECT 2912.720 2880.395 2914.100 2880.565 ;
        RECT 5.605 2879.645 6.815 2880.395 ;
        RECT 2912.805 2879.645 2914.015 2880.395 ;
        RECT 5.605 2879.105 6.125 2879.645 ;
        RECT 2913.495 2879.105 2914.015 2879.645 ;
        RECT 5.605 2875.875 6.125 2876.415 ;
        RECT 2913.495 2875.875 2914.015 2876.415 ;
        RECT 5.605 2875.125 6.815 2875.875 ;
        RECT 2910.045 2875.125 2910.335 2875.850 ;
        RECT 2912.805 2875.125 2914.015 2875.875 ;
        RECT 5.520 2874.955 6.900 2875.125 ;
        RECT 2909.960 2874.955 2910.420 2875.125 ;
        RECT 2912.720 2874.955 2914.100 2875.125 ;
        RECT 5.605 2874.205 6.815 2874.955 ;
        RECT 2912.805 2874.205 2914.015 2874.955 ;
        RECT 5.605 2873.665 6.125 2874.205 ;
        RECT 2913.495 2873.665 2914.015 2874.205 ;
        RECT 5.605 2870.435 6.125 2870.975 ;
        RECT 2913.495 2870.435 2914.015 2870.975 ;
        RECT 5.605 2869.685 6.815 2870.435 ;
        RECT 9.515 2869.685 9.855 2870.345 ;
        RECT 2910.045 2869.685 2910.335 2870.410 ;
        RECT 2912.805 2869.685 2914.015 2870.435 ;
        RECT 5.520 2869.515 6.900 2869.685 ;
        RECT 8.740 2869.515 10.120 2869.685 ;
        RECT 2909.960 2869.515 2910.420 2869.685 ;
        RECT 2912.720 2869.515 2914.100 2869.685 ;
        RECT 5.605 2868.765 6.815 2869.515 ;
        RECT 2912.805 2868.765 2914.015 2869.515 ;
        RECT 5.605 2868.225 6.125 2868.765 ;
        RECT 2913.495 2868.225 2914.015 2868.765 ;
        RECT 5.605 2864.995 6.125 2865.535 ;
        RECT 2913.495 2864.995 2914.015 2865.535 ;
        RECT 5.605 2864.245 6.815 2864.995 ;
        RECT 2910.045 2864.245 2910.335 2864.970 ;
        RECT 2912.805 2864.245 2914.015 2864.995 ;
        RECT 5.520 2864.075 6.900 2864.245 ;
        RECT 2909.960 2864.075 2910.420 2864.245 ;
        RECT 2912.720 2864.075 2914.100 2864.245 ;
        RECT 5.605 2863.325 6.815 2864.075 ;
        RECT 2912.805 2863.325 2914.015 2864.075 ;
        RECT 5.605 2862.785 6.125 2863.325 ;
        RECT 2913.495 2862.785 2914.015 2863.325 ;
        RECT 5.605 2859.555 6.125 2860.095 ;
        RECT 2913.495 2859.555 2914.015 2860.095 ;
        RECT 5.605 2858.805 6.815 2859.555 ;
        RECT 2910.045 2858.805 2910.335 2859.530 ;
        RECT 2912.805 2858.805 2914.015 2859.555 ;
        RECT 5.520 2858.635 6.900 2858.805 ;
        RECT 2909.960 2858.635 2910.420 2858.805 ;
        RECT 2912.720 2858.635 2914.100 2858.805 ;
        RECT 5.605 2857.885 6.815 2858.635 ;
        RECT 2912.805 2857.885 2914.015 2858.635 ;
        RECT 5.605 2857.345 6.125 2857.885 ;
        RECT 2913.495 2857.345 2914.015 2857.885 ;
        RECT 5.605 2854.115 6.125 2854.655 ;
        RECT 2913.495 2854.115 2914.015 2854.655 ;
        RECT 5.605 2853.365 6.815 2854.115 ;
        RECT 2910.045 2853.365 2910.335 2854.090 ;
        RECT 2912.805 2853.365 2914.015 2854.115 ;
        RECT 5.520 2853.195 6.900 2853.365 ;
        RECT 2909.960 2853.195 2910.420 2853.365 ;
        RECT 2912.720 2853.195 2914.100 2853.365 ;
        RECT 5.605 2852.445 6.815 2853.195 ;
        RECT 2912.805 2852.445 2914.015 2853.195 ;
        RECT 5.605 2851.905 6.125 2852.445 ;
        RECT 2913.495 2851.905 2914.015 2852.445 ;
        RECT 5.605 2848.675 6.125 2849.215 ;
        RECT 2913.495 2848.675 2914.015 2849.215 ;
        RECT 5.605 2847.925 6.815 2848.675 ;
        RECT 2910.045 2847.925 2910.335 2848.650 ;
        RECT 2912.805 2847.925 2914.015 2848.675 ;
        RECT 5.520 2847.755 6.900 2847.925 ;
        RECT 2909.960 2847.755 2910.420 2847.925 ;
        RECT 2912.720 2847.755 2914.100 2847.925 ;
        RECT 5.605 2847.005 6.815 2847.755 ;
        RECT 2912.805 2847.005 2914.015 2847.755 ;
        RECT 5.605 2846.465 6.125 2847.005 ;
        RECT 2913.495 2846.465 2914.015 2847.005 ;
        RECT 5.605 2843.235 6.125 2843.775 ;
        RECT 2913.495 2843.235 2914.015 2843.775 ;
        RECT 5.605 2842.485 6.815 2843.235 ;
        RECT 2910.045 2842.485 2910.335 2843.210 ;
        RECT 2912.805 2842.485 2914.015 2843.235 ;
        RECT 5.520 2842.315 6.900 2842.485 ;
        RECT 2909.960 2842.315 2910.420 2842.485 ;
        RECT 2912.720 2842.315 2914.100 2842.485 ;
        RECT 5.605 2841.565 6.815 2842.315 ;
        RECT 2912.805 2841.565 2914.015 2842.315 ;
        RECT 5.605 2841.025 6.125 2841.565 ;
        RECT 2913.495 2841.025 2914.015 2841.565 ;
        RECT 5.605 2837.795 6.125 2838.335 ;
        RECT 2913.495 2837.795 2914.015 2838.335 ;
        RECT 5.605 2837.045 6.815 2837.795 ;
        RECT 2910.045 2837.045 2910.335 2837.770 ;
        RECT 2912.805 2837.045 2914.015 2837.795 ;
        RECT 5.520 2836.875 6.900 2837.045 ;
        RECT 2909.960 2836.875 2910.420 2837.045 ;
        RECT 2912.720 2836.875 2914.100 2837.045 ;
        RECT 5.605 2836.125 6.815 2836.875 ;
        RECT 2912.805 2836.125 2914.015 2836.875 ;
        RECT 5.605 2835.585 6.125 2836.125 ;
        RECT 2913.495 2835.585 2914.015 2836.125 ;
        RECT 5.605 2832.355 6.125 2832.895 ;
        RECT 2913.495 2832.355 2914.015 2832.895 ;
        RECT 5.605 2831.605 6.815 2832.355 ;
        RECT 2910.045 2831.605 2910.335 2832.330 ;
        RECT 2912.805 2831.605 2914.015 2832.355 ;
        RECT 5.520 2831.435 6.900 2831.605 ;
        RECT 2909.960 2831.435 2910.420 2831.605 ;
        RECT 2912.720 2831.435 2914.100 2831.605 ;
        RECT 5.605 2830.685 6.815 2831.435 ;
        RECT 2912.805 2830.685 2914.015 2831.435 ;
        RECT 5.605 2830.145 6.125 2830.685 ;
        RECT 2913.495 2830.145 2914.015 2830.685 ;
        RECT 5.605 2826.915 6.125 2827.455 ;
        RECT 2913.495 2826.915 2914.015 2827.455 ;
        RECT 5.605 2826.165 6.815 2826.915 ;
        RECT 2910.045 2826.165 2910.335 2826.890 ;
        RECT 2912.805 2826.165 2914.015 2826.915 ;
        RECT 5.520 2825.995 6.900 2826.165 ;
        RECT 2909.960 2825.995 2910.420 2826.165 ;
        RECT 2912.720 2825.995 2914.100 2826.165 ;
        RECT 5.605 2825.245 6.815 2825.995 ;
        RECT 2912.805 2825.245 2914.015 2825.995 ;
        RECT 5.605 2824.705 6.125 2825.245 ;
        RECT 2913.495 2824.705 2914.015 2825.245 ;
        RECT 5.605 2821.475 6.125 2822.015 ;
        RECT 2913.495 2821.475 2914.015 2822.015 ;
        RECT 5.605 2820.725 6.815 2821.475 ;
        RECT 2910.045 2820.725 2910.335 2821.450 ;
        RECT 2912.805 2820.725 2914.015 2821.475 ;
        RECT 5.520 2820.555 6.900 2820.725 ;
        RECT 2909.960 2820.555 2910.420 2820.725 ;
        RECT 2912.720 2820.555 2914.100 2820.725 ;
        RECT 5.605 2819.805 6.815 2820.555 ;
        RECT 2912.805 2819.805 2914.015 2820.555 ;
        RECT 5.605 2819.265 6.125 2819.805 ;
        RECT 2913.495 2819.265 2914.015 2819.805 ;
        RECT 5.605 2816.035 6.125 2816.575 ;
        RECT 2913.495 2816.035 2914.015 2816.575 ;
        RECT 5.605 2815.285 6.815 2816.035 ;
        RECT 2910.045 2815.285 2910.335 2816.010 ;
        RECT 2912.805 2815.285 2914.015 2816.035 ;
        RECT 5.520 2815.115 6.900 2815.285 ;
        RECT 2909.960 2815.115 2910.420 2815.285 ;
        RECT 2912.720 2815.115 2914.100 2815.285 ;
        RECT 5.605 2814.365 6.815 2815.115 ;
        RECT 2912.805 2814.365 2914.015 2815.115 ;
        RECT 5.605 2813.825 6.125 2814.365 ;
        RECT 2913.495 2813.825 2914.015 2814.365 ;
        RECT 5.605 2810.595 6.125 2811.135 ;
        RECT 2913.495 2810.595 2914.015 2811.135 ;
        RECT 5.605 2809.845 6.815 2810.595 ;
        RECT 2910.045 2809.845 2910.335 2810.570 ;
        RECT 2912.805 2809.845 2914.015 2810.595 ;
        RECT 5.520 2809.675 6.900 2809.845 ;
        RECT 2909.960 2809.675 2910.420 2809.845 ;
        RECT 2912.720 2809.675 2914.100 2809.845 ;
        RECT 5.605 2808.925 6.815 2809.675 ;
        RECT 2912.805 2808.925 2914.015 2809.675 ;
        RECT 5.605 2808.385 6.125 2808.925 ;
        RECT 2913.495 2808.385 2914.015 2808.925 ;
        RECT 5.605 2805.155 6.125 2805.695 ;
        RECT 2913.495 2805.155 2914.015 2805.695 ;
        RECT 5.605 2804.405 6.815 2805.155 ;
        RECT 2910.045 2804.405 2910.335 2805.130 ;
        RECT 2912.805 2804.405 2914.015 2805.155 ;
        RECT 5.520 2804.235 6.900 2804.405 ;
        RECT 2909.960 2804.235 2910.420 2804.405 ;
        RECT 2912.720 2804.235 2914.100 2804.405 ;
        RECT 5.605 2803.485 6.815 2804.235 ;
        RECT 2912.805 2803.485 2914.015 2804.235 ;
        RECT 5.605 2802.945 6.125 2803.485 ;
        RECT 2913.495 2802.945 2914.015 2803.485 ;
        RECT 5.605 2799.715 6.125 2800.255 ;
        RECT 2913.495 2799.715 2914.015 2800.255 ;
        RECT 5.605 2798.965 6.815 2799.715 ;
        RECT 2910.045 2798.965 2910.335 2799.690 ;
        RECT 2912.805 2798.965 2914.015 2799.715 ;
        RECT 5.520 2798.795 6.900 2798.965 ;
        RECT 2909.960 2798.795 2910.420 2798.965 ;
        RECT 2912.720 2798.795 2914.100 2798.965 ;
        RECT 5.605 2798.045 6.815 2798.795 ;
        RECT 2912.805 2798.045 2914.015 2798.795 ;
        RECT 5.605 2797.505 6.125 2798.045 ;
        RECT 2913.495 2797.505 2914.015 2798.045 ;
        RECT 5.605 2794.275 6.125 2794.815 ;
        RECT 2913.495 2794.275 2914.015 2794.815 ;
        RECT 5.605 2793.525 6.815 2794.275 ;
        RECT 2910.045 2793.525 2910.335 2794.250 ;
        RECT 2912.805 2793.525 2914.015 2794.275 ;
        RECT 5.520 2793.355 6.900 2793.525 ;
        RECT 2909.960 2793.355 2910.420 2793.525 ;
        RECT 2912.720 2793.355 2914.100 2793.525 ;
        RECT 5.605 2792.605 6.815 2793.355 ;
        RECT 2912.805 2792.605 2914.015 2793.355 ;
        RECT 5.605 2792.065 6.125 2792.605 ;
        RECT 2913.495 2792.065 2914.015 2792.605 ;
        RECT 5.605 2788.835 6.125 2789.375 ;
        RECT 2913.495 2788.835 2914.015 2789.375 ;
        RECT 5.605 2788.085 6.815 2788.835 ;
        RECT 2910.045 2788.085 2910.335 2788.810 ;
        RECT 2912.805 2788.085 2914.015 2788.835 ;
        RECT 5.520 2787.915 6.900 2788.085 ;
        RECT 2909.960 2787.915 2910.420 2788.085 ;
        RECT 2912.720 2787.915 2914.100 2788.085 ;
        RECT 5.605 2787.165 6.815 2787.915 ;
        RECT 2912.805 2787.165 2914.015 2787.915 ;
        RECT 5.605 2786.625 6.125 2787.165 ;
        RECT 2913.495 2786.625 2914.015 2787.165 ;
        RECT 5.605 2783.395 6.125 2783.935 ;
        RECT 2913.495 2783.395 2914.015 2783.935 ;
        RECT 5.605 2782.645 6.815 2783.395 ;
        RECT 2910.045 2782.645 2910.335 2783.370 ;
        RECT 2912.805 2782.645 2914.015 2783.395 ;
        RECT 5.520 2782.475 6.900 2782.645 ;
        RECT 2909.960 2782.475 2910.420 2782.645 ;
        RECT 2912.720 2782.475 2914.100 2782.645 ;
        RECT 5.605 2781.725 6.815 2782.475 ;
        RECT 2912.805 2781.725 2914.015 2782.475 ;
        RECT 5.605 2781.185 6.125 2781.725 ;
        RECT 2913.495 2781.185 2914.015 2781.725 ;
        RECT 5.605 2777.955 6.125 2778.495 ;
        RECT 2913.495 2777.955 2914.015 2778.495 ;
        RECT 5.605 2777.205 6.815 2777.955 ;
        RECT 2910.045 2777.205 2910.335 2777.930 ;
        RECT 2912.805 2777.205 2914.015 2777.955 ;
        RECT 5.520 2777.035 6.900 2777.205 ;
        RECT 2909.040 2777.035 2910.420 2777.205 ;
        RECT 2912.720 2777.035 2914.100 2777.205 ;
        RECT 5.605 2776.285 6.815 2777.035 ;
        RECT 2909.815 2776.375 2910.155 2777.035 ;
        RECT 2912.805 2776.285 2914.015 2777.035 ;
        RECT 5.605 2775.745 6.125 2776.285 ;
        RECT 2913.495 2775.745 2914.015 2776.285 ;
        RECT 5.605 2772.515 6.125 2773.055 ;
        RECT 2913.495 2772.515 2914.015 2773.055 ;
        RECT 5.605 2771.765 6.815 2772.515 ;
        RECT 2910.045 2771.765 2910.335 2772.490 ;
        RECT 2912.805 2771.765 2914.015 2772.515 ;
        RECT 5.520 2771.595 6.900 2771.765 ;
        RECT 2909.960 2771.595 2910.420 2771.765 ;
        RECT 2912.720 2771.595 2914.100 2771.765 ;
        RECT 5.605 2770.845 6.815 2771.595 ;
        RECT 2912.805 2770.845 2914.015 2771.595 ;
        RECT 5.605 2770.305 6.125 2770.845 ;
        RECT 2913.495 2770.305 2914.015 2770.845 ;
        RECT 5.605 2767.075 6.125 2767.615 ;
        RECT 2913.495 2767.075 2914.015 2767.615 ;
        RECT 5.605 2766.325 6.815 2767.075 ;
        RECT 2910.045 2766.325 2910.335 2767.050 ;
        RECT 2912.805 2766.325 2914.015 2767.075 ;
        RECT 5.520 2766.155 6.900 2766.325 ;
        RECT 2909.960 2766.155 2910.420 2766.325 ;
        RECT 2912.720 2766.155 2914.100 2766.325 ;
        RECT 5.605 2765.405 6.815 2766.155 ;
        RECT 2912.805 2765.405 2914.015 2766.155 ;
        RECT 5.605 2764.865 6.125 2765.405 ;
        RECT 2913.495 2764.865 2914.015 2765.405 ;
        RECT 5.605 2761.635 6.125 2762.175 ;
        RECT 2913.495 2761.635 2914.015 2762.175 ;
        RECT 5.605 2760.885 6.815 2761.635 ;
        RECT 2910.045 2760.885 2910.335 2761.610 ;
        RECT 2912.805 2760.885 2914.015 2761.635 ;
        RECT 5.520 2760.715 6.900 2760.885 ;
        RECT 2909.960 2760.715 2910.420 2760.885 ;
        RECT 2912.720 2760.715 2914.100 2760.885 ;
        RECT 5.605 2759.965 6.815 2760.715 ;
        RECT 2912.805 2759.965 2914.015 2760.715 ;
        RECT 5.605 2759.425 6.125 2759.965 ;
        RECT 2913.495 2759.425 2914.015 2759.965 ;
        RECT 5.605 2756.195 6.125 2756.735 ;
        RECT 2913.495 2756.195 2914.015 2756.735 ;
        RECT 5.605 2755.445 6.815 2756.195 ;
        RECT 2910.045 2755.445 2910.335 2756.170 ;
        RECT 2912.805 2755.445 2914.015 2756.195 ;
        RECT 5.520 2755.275 6.900 2755.445 ;
        RECT 2909.960 2755.275 2910.420 2755.445 ;
        RECT 2912.720 2755.275 2914.100 2755.445 ;
        RECT 5.605 2754.525 6.815 2755.275 ;
        RECT 2912.805 2754.525 2914.015 2755.275 ;
        RECT 5.605 2753.985 6.125 2754.525 ;
        RECT 2913.495 2753.985 2914.015 2754.525 ;
        RECT 5.605 2750.755 6.125 2751.295 ;
        RECT 2913.495 2750.755 2914.015 2751.295 ;
        RECT 5.605 2750.005 6.815 2750.755 ;
        RECT 2910.045 2750.005 2910.335 2750.730 ;
        RECT 2912.805 2750.005 2914.015 2750.755 ;
        RECT 5.520 2749.835 6.900 2750.005 ;
        RECT 2909.960 2749.835 2910.420 2750.005 ;
        RECT 2912.720 2749.835 2914.100 2750.005 ;
        RECT 5.605 2749.085 6.815 2749.835 ;
        RECT 2912.805 2749.085 2914.015 2749.835 ;
        RECT 5.605 2748.545 6.125 2749.085 ;
        RECT 2913.495 2748.545 2914.015 2749.085 ;
        RECT 5.605 2745.315 6.125 2745.855 ;
        RECT 2913.495 2745.315 2914.015 2745.855 ;
        RECT 5.605 2744.565 6.815 2745.315 ;
        RECT 2910.045 2744.565 2910.335 2745.290 ;
        RECT 2912.805 2744.565 2914.015 2745.315 ;
        RECT 5.520 2744.395 6.900 2744.565 ;
        RECT 2909.960 2744.395 2910.420 2744.565 ;
        RECT 2912.720 2744.395 2914.100 2744.565 ;
        RECT 5.605 2743.645 6.815 2744.395 ;
        RECT 2912.805 2743.645 2914.015 2744.395 ;
        RECT 5.605 2743.105 6.125 2743.645 ;
        RECT 2913.495 2743.105 2914.015 2743.645 ;
        RECT 5.605 2739.875 6.125 2740.415 ;
        RECT 2913.495 2739.875 2914.015 2740.415 ;
        RECT 5.605 2739.125 6.815 2739.875 ;
        RECT 2910.045 2739.125 2910.335 2739.850 ;
        RECT 2912.805 2739.125 2914.015 2739.875 ;
        RECT 5.520 2738.955 6.900 2739.125 ;
        RECT 2909.960 2738.955 2910.420 2739.125 ;
        RECT 2912.720 2738.955 2914.100 2739.125 ;
        RECT 5.605 2738.205 6.815 2738.955 ;
        RECT 2912.805 2738.205 2914.015 2738.955 ;
        RECT 5.605 2737.665 6.125 2738.205 ;
        RECT 2913.495 2737.665 2914.015 2738.205 ;
        RECT 5.605 2734.435 6.125 2734.975 ;
        RECT 2913.495 2734.435 2914.015 2734.975 ;
        RECT 5.605 2733.685 6.815 2734.435 ;
        RECT 2910.045 2733.685 2910.335 2734.410 ;
        RECT 2912.805 2733.685 2914.015 2734.435 ;
        RECT 5.520 2733.515 6.900 2733.685 ;
        RECT 2909.960 2733.515 2910.420 2733.685 ;
        RECT 2912.720 2733.515 2914.100 2733.685 ;
        RECT 5.605 2732.765 6.815 2733.515 ;
        RECT 2912.805 2732.765 2914.015 2733.515 ;
        RECT 5.605 2732.225 6.125 2732.765 ;
        RECT 2913.495 2732.225 2914.015 2732.765 ;
        RECT 5.605 2728.995 6.125 2729.535 ;
        RECT 2913.495 2728.995 2914.015 2729.535 ;
        RECT 5.605 2728.245 6.815 2728.995 ;
        RECT 2910.045 2728.245 2910.335 2728.970 ;
        RECT 2912.805 2728.245 2914.015 2728.995 ;
        RECT 5.520 2728.075 6.900 2728.245 ;
        RECT 2909.960 2728.075 2910.420 2728.245 ;
        RECT 2912.720 2728.075 2914.100 2728.245 ;
        RECT 5.605 2727.325 6.815 2728.075 ;
        RECT 2912.805 2727.325 2914.015 2728.075 ;
        RECT 5.605 2726.785 6.125 2727.325 ;
        RECT 2913.495 2726.785 2914.015 2727.325 ;
        RECT 5.605 2723.555 6.125 2724.095 ;
        RECT 2913.495 2723.555 2914.015 2724.095 ;
        RECT 5.605 2722.805 6.815 2723.555 ;
        RECT 2910.045 2722.805 2910.335 2723.530 ;
        RECT 2912.805 2722.805 2914.015 2723.555 ;
        RECT 5.520 2722.635 6.900 2722.805 ;
        RECT 2909.960 2722.635 2910.420 2722.805 ;
        RECT 2912.720 2722.635 2914.100 2722.805 ;
        RECT 5.605 2721.885 6.815 2722.635 ;
        RECT 2912.805 2721.885 2914.015 2722.635 ;
        RECT 5.605 2721.345 6.125 2721.885 ;
        RECT 2913.495 2721.345 2914.015 2721.885 ;
        RECT 5.605 2718.115 6.125 2718.655 ;
        RECT 2913.495 2718.115 2914.015 2718.655 ;
        RECT 5.605 2717.365 6.815 2718.115 ;
        RECT 2910.045 2717.365 2910.335 2718.090 ;
        RECT 2912.805 2717.365 2914.015 2718.115 ;
        RECT 5.520 2717.195 6.900 2717.365 ;
        RECT 2909.960 2717.195 2910.420 2717.365 ;
        RECT 2912.720 2717.195 2914.100 2717.365 ;
        RECT 5.605 2716.445 6.815 2717.195 ;
        RECT 2912.805 2716.445 2914.015 2717.195 ;
        RECT 5.605 2715.905 6.125 2716.445 ;
        RECT 2913.495 2715.905 2914.015 2716.445 ;
        RECT 5.605 2712.675 6.125 2713.215 ;
        RECT 2913.495 2712.675 2914.015 2713.215 ;
        RECT 5.605 2711.925 6.815 2712.675 ;
        RECT 2910.045 2711.925 2910.335 2712.650 ;
        RECT 2912.805 2711.925 2914.015 2712.675 ;
        RECT 5.520 2711.755 6.900 2711.925 ;
        RECT 2909.960 2711.755 2910.420 2711.925 ;
        RECT 2912.720 2711.755 2914.100 2711.925 ;
        RECT 5.605 2711.005 6.815 2711.755 ;
        RECT 2912.805 2711.005 2914.015 2711.755 ;
        RECT 5.605 2710.465 6.125 2711.005 ;
        RECT 2913.495 2710.465 2914.015 2711.005 ;
        RECT 5.605 2707.235 6.125 2707.775 ;
        RECT 2913.495 2707.235 2914.015 2707.775 ;
        RECT 5.605 2706.485 6.815 2707.235 ;
        RECT 2910.045 2706.485 2910.335 2707.210 ;
        RECT 2912.805 2706.485 2914.015 2707.235 ;
        RECT 5.520 2706.315 6.900 2706.485 ;
        RECT 2909.960 2706.315 2910.420 2706.485 ;
        RECT 2912.720 2706.315 2914.100 2706.485 ;
        RECT 5.605 2705.565 6.815 2706.315 ;
        RECT 2912.805 2705.565 2914.015 2706.315 ;
        RECT 5.605 2705.025 6.125 2705.565 ;
        RECT 2913.495 2705.025 2914.015 2705.565 ;
        RECT 5.605 2701.795 6.125 2702.335 ;
        RECT 2913.495 2701.795 2914.015 2702.335 ;
        RECT 5.605 2701.045 6.815 2701.795 ;
        RECT 2910.045 2701.045 2910.335 2701.770 ;
        RECT 2912.805 2701.045 2914.015 2701.795 ;
        RECT 5.520 2700.875 6.900 2701.045 ;
        RECT 2909.960 2700.875 2910.420 2701.045 ;
        RECT 2912.720 2700.875 2914.100 2701.045 ;
        RECT 5.605 2700.125 6.815 2700.875 ;
        RECT 2912.805 2700.125 2914.015 2700.875 ;
        RECT 5.605 2699.585 6.125 2700.125 ;
        RECT 2913.495 2699.585 2914.015 2700.125 ;
        RECT 5.605 2696.355 6.125 2696.895 ;
        RECT 2913.495 2696.355 2914.015 2696.895 ;
        RECT 5.605 2695.605 6.815 2696.355 ;
        RECT 2910.045 2695.605 2910.335 2696.330 ;
        RECT 2912.805 2695.605 2914.015 2696.355 ;
        RECT 5.520 2695.435 6.900 2695.605 ;
        RECT 2909.960 2695.435 2910.420 2695.605 ;
        RECT 2912.720 2695.435 2914.100 2695.605 ;
        RECT 5.605 2694.685 6.815 2695.435 ;
        RECT 2912.805 2694.685 2914.015 2695.435 ;
        RECT 5.605 2694.145 6.125 2694.685 ;
        RECT 2913.495 2694.145 2914.015 2694.685 ;
        RECT 5.605 2690.915 6.125 2691.455 ;
        RECT 2913.495 2690.915 2914.015 2691.455 ;
        RECT 5.605 2690.165 6.815 2690.915 ;
        RECT 2912.805 2690.165 2914.015 2690.915 ;
        RECT 5.520 2689.995 6.900 2690.165 ;
        RECT 2906.300 2689.995 2906.740 2690.165 ;
        RECT 2912.720 2689.995 2914.100 2690.165 ;
        RECT 5.605 2689.245 6.815 2689.995 ;
        RECT 2906.365 2689.270 2906.655 2689.995 ;
        RECT 2912.805 2689.245 2914.015 2689.995 ;
        RECT 5.605 2688.705 6.125 2689.245 ;
        RECT 2913.495 2688.705 2914.015 2689.245 ;
        RECT 5.605 2685.475 6.125 2686.015 ;
        RECT 2913.495 2685.475 2914.015 2686.015 ;
        RECT 5.605 2684.725 6.815 2685.475 ;
        RECT 2912.805 2684.725 2914.015 2685.475 ;
        RECT 5.520 2684.555 6.900 2684.725 ;
        RECT 2906.300 2684.555 2906.740 2684.725 ;
        RECT 2912.720 2684.555 2914.100 2684.725 ;
        RECT 5.605 2683.805 6.815 2684.555 ;
        RECT 2906.365 2683.830 2906.655 2684.555 ;
        RECT 2912.805 2683.805 2914.015 2684.555 ;
        RECT 5.605 2683.265 6.125 2683.805 ;
        RECT 2913.495 2683.265 2914.015 2683.805 ;
        RECT 5.605 2680.035 6.125 2680.575 ;
        RECT 2913.495 2680.035 2914.015 2680.575 ;
        RECT 5.605 2679.285 6.815 2680.035 ;
        RECT 2912.805 2679.285 2914.015 2680.035 ;
        RECT 5.520 2679.115 6.900 2679.285 ;
        RECT 2906.300 2679.115 2906.740 2679.285 ;
        RECT 2912.720 2679.115 2914.100 2679.285 ;
        RECT 5.605 2678.365 6.815 2679.115 ;
        RECT 2906.365 2678.390 2906.655 2679.115 ;
        RECT 2912.805 2678.365 2914.015 2679.115 ;
        RECT 5.605 2677.825 6.125 2678.365 ;
        RECT 2913.495 2677.825 2914.015 2678.365 ;
        RECT 5.605 2674.595 6.125 2675.135 ;
        RECT 2913.495 2674.595 2914.015 2675.135 ;
        RECT 5.605 2673.845 6.815 2674.595 ;
        RECT 2912.805 2673.845 2914.015 2674.595 ;
        RECT 5.520 2673.675 6.900 2673.845 ;
        RECT 2906.300 2673.675 2906.740 2673.845 ;
        RECT 2912.720 2673.675 2914.100 2673.845 ;
        RECT 5.605 2672.925 6.815 2673.675 ;
        RECT 2906.365 2672.950 2906.655 2673.675 ;
        RECT 2912.805 2672.925 2914.015 2673.675 ;
        RECT 5.605 2672.385 6.125 2672.925 ;
        RECT 2913.495 2672.385 2914.015 2672.925 ;
        RECT 5.605 2669.155 6.125 2669.695 ;
        RECT 2913.495 2669.155 2914.015 2669.695 ;
        RECT 5.605 2668.405 6.815 2669.155 ;
        RECT 2912.805 2668.405 2914.015 2669.155 ;
        RECT 5.520 2668.235 6.900 2668.405 ;
        RECT 2906.300 2668.235 2906.740 2668.405 ;
        RECT 2912.720 2668.235 2914.100 2668.405 ;
        RECT 5.605 2667.485 6.815 2668.235 ;
        RECT 2906.365 2667.510 2906.655 2668.235 ;
        RECT 2912.805 2667.485 2914.015 2668.235 ;
        RECT 5.605 2666.945 6.125 2667.485 ;
        RECT 2913.495 2666.945 2914.015 2667.485 ;
        RECT 5.605 2663.715 6.125 2664.255 ;
        RECT 2913.495 2663.715 2914.015 2664.255 ;
        RECT 5.605 2662.965 6.815 2663.715 ;
        RECT 2912.805 2662.965 2914.015 2663.715 ;
        RECT 5.520 2662.795 6.900 2662.965 ;
        RECT 2906.300 2662.795 2906.740 2662.965 ;
        RECT 2912.720 2662.795 2914.100 2662.965 ;
        RECT 5.605 2662.045 6.815 2662.795 ;
        RECT 2906.365 2662.070 2906.655 2662.795 ;
        RECT 2912.805 2662.045 2914.015 2662.795 ;
        RECT 5.605 2661.505 6.125 2662.045 ;
        RECT 2913.495 2661.505 2914.015 2662.045 ;
        RECT 5.605 2658.275 6.125 2658.815 ;
        RECT 2913.495 2658.275 2914.015 2658.815 ;
        RECT 5.605 2657.525 6.815 2658.275 ;
        RECT 2912.805 2657.525 2914.015 2658.275 ;
        RECT 5.520 2657.355 6.900 2657.525 ;
        RECT 2906.300 2657.355 2906.740 2657.525 ;
        RECT 2912.720 2657.355 2914.100 2657.525 ;
        RECT 5.605 2656.605 6.815 2657.355 ;
        RECT 2906.365 2656.630 2906.655 2657.355 ;
        RECT 2912.805 2656.605 2914.015 2657.355 ;
        RECT 5.605 2656.065 6.125 2656.605 ;
        RECT 2913.495 2656.065 2914.015 2656.605 ;
        RECT 5.605 2652.835 6.125 2653.375 ;
        RECT 2913.495 2652.835 2914.015 2653.375 ;
        RECT 5.605 2652.085 6.815 2652.835 ;
        RECT 2912.805 2652.085 2914.015 2652.835 ;
        RECT 5.520 2651.915 6.900 2652.085 ;
        RECT 2906.300 2651.915 2906.740 2652.085 ;
        RECT 2912.720 2651.915 2914.100 2652.085 ;
        RECT 5.605 2651.165 6.815 2651.915 ;
        RECT 2906.365 2651.190 2906.655 2651.915 ;
        RECT 2912.805 2651.165 2914.015 2651.915 ;
        RECT 5.605 2650.625 6.125 2651.165 ;
        RECT 2913.495 2650.625 2914.015 2651.165 ;
        RECT 5.605 2647.395 6.125 2647.935 ;
        RECT 2913.495 2647.395 2914.015 2647.935 ;
        RECT 5.605 2646.645 6.815 2647.395 ;
        RECT 2912.805 2646.645 2914.015 2647.395 ;
        RECT 5.520 2646.475 6.900 2646.645 ;
        RECT 2906.300 2646.475 2906.740 2646.645 ;
        RECT 2912.720 2646.475 2914.100 2646.645 ;
        RECT 5.605 2645.725 6.815 2646.475 ;
        RECT 2906.365 2645.750 2906.655 2646.475 ;
        RECT 2912.805 2645.725 2914.015 2646.475 ;
        RECT 5.605 2645.185 6.125 2645.725 ;
        RECT 2913.495 2645.185 2914.015 2645.725 ;
        RECT 5.605 2641.955 6.125 2642.495 ;
        RECT 2913.495 2641.955 2914.015 2642.495 ;
        RECT 5.605 2641.205 6.815 2641.955 ;
        RECT 2912.805 2641.205 2914.015 2641.955 ;
        RECT 5.520 2641.035 6.900 2641.205 ;
        RECT 2906.300 2641.035 2906.740 2641.205 ;
        RECT 2912.720 2641.035 2914.100 2641.205 ;
        RECT 5.605 2640.285 6.815 2641.035 ;
        RECT 2906.365 2640.310 2906.655 2641.035 ;
        RECT 2912.805 2640.285 2914.015 2641.035 ;
        RECT 5.605 2639.745 6.125 2640.285 ;
        RECT 2913.495 2639.745 2914.015 2640.285 ;
        RECT 5.605 2636.515 6.125 2637.055 ;
        RECT 2913.495 2636.515 2914.015 2637.055 ;
        RECT 5.605 2635.765 6.815 2636.515 ;
        RECT 2912.805 2635.765 2914.015 2636.515 ;
        RECT 5.520 2635.595 6.900 2635.765 ;
        RECT 2906.300 2635.595 2906.740 2635.765 ;
        RECT 2912.720 2635.595 2914.100 2635.765 ;
        RECT 5.605 2634.845 6.815 2635.595 ;
        RECT 2906.365 2634.870 2906.655 2635.595 ;
        RECT 2912.805 2634.845 2914.015 2635.595 ;
        RECT 5.605 2634.305 6.125 2634.845 ;
        RECT 2913.495 2634.305 2914.015 2634.845 ;
        RECT 5.605 2631.075 6.125 2631.615 ;
        RECT 2913.495 2631.075 2914.015 2631.615 ;
        RECT 5.605 2630.325 6.815 2631.075 ;
        RECT 2912.805 2630.325 2914.015 2631.075 ;
        RECT 5.520 2630.155 6.900 2630.325 ;
        RECT 2906.300 2630.155 2906.740 2630.325 ;
        RECT 2909.040 2630.155 2910.420 2630.325 ;
        RECT 2912.720 2630.155 2914.100 2630.325 ;
        RECT 5.605 2629.405 6.815 2630.155 ;
        RECT 2906.365 2629.430 2906.655 2630.155 ;
        RECT 2909.815 2629.495 2910.155 2630.155 ;
        RECT 2912.805 2629.405 2914.015 2630.155 ;
        RECT 5.605 2628.865 6.125 2629.405 ;
        RECT 2913.495 2628.865 2914.015 2629.405 ;
        RECT 5.605 2625.635 6.125 2626.175 ;
        RECT 2913.495 2625.635 2914.015 2626.175 ;
        RECT 5.605 2624.885 6.815 2625.635 ;
        RECT 2912.805 2624.885 2914.015 2625.635 ;
        RECT 5.520 2624.715 6.900 2624.885 ;
        RECT 2906.300 2624.715 2906.740 2624.885 ;
        RECT 2912.720 2624.715 2914.100 2624.885 ;
        RECT 5.605 2623.965 6.815 2624.715 ;
        RECT 2906.365 2623.990 2906.655 2624.715 ;
        RECT 2912.805 2623.965 2914.015 2624.715 ;
        RECT 5.605 2623.425 6.125 2623.965 ;
        RECT 2913.495 2623.425 2914.015 2623.965 ;
        RECT 5.605 2620.195 6.125 2620.735 ;
        RECT 2913.495 2620.195 2914.015 2620.735 ;
        RECT 5.605 2619.445 6.815 2620.195 ;
        RECT 2912.805 2619.445 2914.015 2620.195 ;
        RECT 5.520 2619.275 6.900 2619.445 ;
        RECT 2906.300 2619.275 2906.740 2619.445 ;
        RECT 2912.720 2619.275 2914.100 2619.445 ;
        RECT 5.605 2618.525 6.815 2619.275 ;
        RECT 2906.365 2618.550 2906.655 2619.275 ;
        RECT 2912.805 2618.525 2914.015 2619.275 ;
        RECT 5.605 2617.985 6.125 2618.525 ;
        RECT 2913.495 2617.985 2914.015 2618.525 ;
        RECT 5.605 2614.755 6.125 2615.295 ;
        RECT 2913.495 2614.755 2914.015 2615.295 ;
        RECT 5.605 2614.005 6.815 2614.755 ;
        RECT 2912.805 2614.005 2914.015 2614.755 ;
        RECT 5.520 2613.835 6.900 2614.005 ;
        RECT 2906.300 2613.835 2906.740 2614.005 ;
        RECT 2912.720 2613.835 2914.100 2614.005 ;
        RECT 5.605 2613.085 6.815 2613.835 ;
        RECT 2906.365 2613.110 2906.655 2613.835 ;
        RECT 2912.805 2613.085 2914.015 2613.835 ;
        RECT 5.605 2612.545 6.125 2613.085 ;
        RECT 2913.495 2612.545 2914.015 2613.085 ;
        RECT 5.605 2609.315 6.125 2609.855 ;
        RECT 2913.495 2609.315 2914.015 2609.855 ;
        RECT 5.605 2608.565 6.815 2609.315 ;
        RECT 2912.805 2608.565 2914.015 2609.315 ;
        RECT 5.520 2608.395 6.900 2608.565 ;
        RECT 2906.300 2608.395 2906.740 2608.565 ;
        RECT 2912.720 2608.395 2914.100 2608.565 ;
        RECT 5.605 2607.645 6.815 2608.395 ;
        RECT 2906.365 2607.670 2906.655 2608.395 ;
        RECT 2912.805 2607.645 2914.015 2608.395 ;
        RECT 5.605 2607.105 6.125 2607.645 ;
        RECT 2913.495 2607.105 2914.015 2607.645 ;
        RECT 5.605 2603.875 6.125 2604.415 ;
        RECT 2913.495 2603.875 2914.015 2604.415 ;
        RECT 5.605 2603.125 6.815 2603.875 ;
        RECT 2912.805 2603.125 2914.015 2603.875 ;
        RECT 5.520 2602.955 6.900 2603.125 ;
        RECT 2906.300 2602.955 2906.740 2603.125 ;
        RECT 2909.040 2602.955 2910.420 2603.125 ;
        RECT 2912.720 2602.955 2914.100 2603.125 ;
        RECT 5.605 2602.205 6.815 2602.955 ;
        RECT 2906.365 2602.230 2906.655 2602.955 ;
        RECT 2909.815 2602.295 2910.155 2602.955 ;
        RECT 2912.805 2602.205 2914.015 2602.955 ;
        RECT 5.605 2601.665 6.125 2602.205 ;
        RECT 2913.495 2601.665 2914.015 2602.205 ;
        RECT 5.605 2598.435 6.125 2598.975 ;
        RECT 2913.495 2598.435 2914.015 2598.975 ;
        RECT 5.605 2597.685 6.815 2598.435 ;
        RECT 2912.805 2597.685 2914.015 2598.435 ;
        RECT 5.520 2597.515 6.900 2597.685 ;
        RECT 2906.300 2597.515 2906.740 2597.685 ;
        RECT 2912.720 2597.515 2914.100 2597.685 ;
        RECT 5.605 2596.765 6.815 2597.515 ;
        RECT 2906.365 2596.790 2906.655 2597.515 ;
        RECT 2912.805 2596.765 2914.015 2597.515 ;
        RECT 5.605 2596.225 6.125 2596.765 ;
        RECT 2913.495 2596.225 2914.015 2596.765 ;
        RECT 5.605 2592.995 6.125 2593.535 ;
        RECT 2913.495 2592.995 2914.015 2593.535 ;
        RECT 5.605 2592.245 6.815 2592.995 ;
        RECT 2912.805 2592.245 2914.015 2592.995 ;
        RECT 5.520 2592.075 6.900 2592.245 ;
        RECT 2906.300 2592.075 2906.740 2592.245 ;
        RECT 2912.720 2592.075 2914.100 2592.245 ;
        RECT 5.605 2591.325 6.815 2592.075 ;
        RECT 2906.365 2591.350 2906.655 2592.075 ;
        RECT 2912.805 2591.325 2914.015 2592.075 ;
        RECT 5.605 2590.785 6.125 2591.325 ;
        RECT 2913.495 2590.785 2914.015 2591.325 ;
        RECT 5.605 2587.555 6.125 2588.095 ;
        RECT 2913.495 2587.555 2914.015 2588.095 ;
        RECT 5.605 2586.805 6.815 2587.555 ;
        RECT 2912.805 2586.805 2914.015 2587.555 ;
        RECT 5.520 2586.635 6.900 2586.805 ;
        RECT 2906.300 2586.635 2906.740 2586.805 ;
        RECT 2912.720 2586.635 2914.100 2586.805 ;
        RECT 5.605 2585.885 6.815 2586.635 ;
        RECT 2906.365 2585.910 2906.655 2586.635 ;
        RECT 2912.805 2585.885 2914.015 2586.635 ;
        RECT 5.605 2585.345 6.125 2585.885 ;
        RECT 2913.495 2585.345 2914.015 2585.885 ;
        RECT 5.605 2582.115 6.125 2582.655 ;
        RECT 2913.495 2582.115 2914.015 2582.655 ;
        RECT 5.605 2581.365 6.815 2582.115 ;
        RECT 2912.805 2581.365 2914.015 2582.115 ;
        RECT 5.520 2581.195 6.900 2581.365 ;
        RECT 2906.300 2581.195 2906.740 2581.365 ;
        RECT 2912.720 2581.195 2914.100 2581.365 ;
        RECT 5.605 2580.445 6.815 2581.195 ;
        RECT 2906.365 2580.470 2906.655 2581.195 ;
        RECT 2912.805 2580.445 2914.015 2581.195 ;
        RECT 5.605 2579.905 6.125 2580.445 ;
        RECT 2913.495 2579.905 2914.015 2580.445 ;
        RECT 5.605 2576.675 6.125 2577.215 ;
        RECT 2913.495 2576.675 2914.015 2577.215 ;
        RECT 5.605 2575.925 6.815 2576.675 ;
        RECT 2912.805 2575.925 2914.015 2576.675 ;
        RECT 5.520 2575.755 6.900 2575.925 ;
        RECT 2906.300 2575.755 2906.740 2575.925 ;
        RECT 2912.720 2575.755 2914.100 2575.925 ;
        RECT 5.605 2575.005 6.815 2575.755 ;
        RECT 2906.365 2575.030 2906.655 2575.755 ;
        RECT 2912.805 2575.005 2914.015 2575.755 ;
        RECT 5.605 2574.465 6.125 2575.005 ;
        RECT 2913.495 2574.465 2914.015 2575.005 ;
        RECT 5.605 2571.235 6.125 2571.775 ;
        RECT 2913.495 2571.235 2914.015 2571.775 ;
        RECT 5.605 2570.485 6.815 2571.235 ;
        RECT 2912.805 2570.485 2914.015 2571.235 ;
        RECT 5.520 2570.315 6.900 2570.485 ;
        RECT 2906.300 2570.315 2906.740 2570.485 ;
        RECT 2912.720 2570.315 2914.100 2570.485 ;
        RECT 5.605 2569.565 6.815 2570.315 ;
        RECT 2906.365 2569.590 2906.655 2570.315 ;
        RECT 2912.805 2569.565 2914.015 2570.315 ;
        RECT 5.605 2569.025 6.125 2569.565 ;
        RECT 2913.495 2569.025 2914.015 2569.565 ;
        RECT 5.605 2565.795 6.125 2566.335 ;
        RECT 2913.495 2565.795 2914.015 2566.335 ;
        RECT 5.605 2565.045 6.815 2565.795 ;
        RECT 2912.805 2565.045 2914.015 2565.795 ;
        RECT 5.520 2564.875 6.900 2565.045 ;
        RECT 2906.300 2564.875 2906.740 2565.045 ;
        RECT 2912.720 2564.875 2914.100 2565.045 ;
        RECT 5.605 2564.125 6.815 2564.875 ;
        RECT 2906.365 2564.150 2906.655 2564.875 ;
        RECT 2912.805 2564.125 2914.015 2564.875 ;
        RECT 5.605 2563.585 6.125 2564.125 ;
        RECT 2913.495 2563.585 2914.015 2564.125 ;
        RECT 5.605 2560.355 6.125 2560.895 ;
        RECT 2913.495 2560.355 2914.015 2560.895 ;
        RECT 5.605 2559.605 6.815 2560.355 ;
        RECT 2912.805 2559.605 2914.015 2560.355 ;
        RECT 5.520 2559.435 6.900 2559.605 ;
        RECT 2906.300 2559.435 2906.740 2559.605 ;
        RECT 2912.720 2559.435 2914.100 2559.605 ;
        RECT 5.605 2558.685 6.815 2559.435 ;
        RECT 2906.365 2558.710 2906.655 2559.435 ;
        RECT 2912.805 2558.685 2914.015 2559.435 ;
        RECT 5.605 2558.145 6.125 2558.685 ;
        RECT 2913.495 2558.145 2914.015 2558.685 ;
        RECT 5.605 2554.915 6.125 2555.455 ;
        RECT 2913.495 2554.915 2914.015 2555.455 ;
        RECT 5.605 2554.165 6.815 2554.915 ;
        RECT 2912.805 2554.165 2914.015 2554.915 ;
        RECT 5.520 2553.995 6.900 2554.165 ;
        RECT 2906.300 2553.995 2906.740 2554.165 ;
        RECT 2912.720 2553.995 2914.100 2554.165 ;
        RECT 5.605 2553.245 6.815 2553.995 ;
        RECT 2906.365 2553.270 2906.655 2553.995 ;
        RECT 2912.805 2553.245 2914.015 2553.995 ;
        RECT 5.605 2552.705 6.125 2553.245 ;
        RECT 2913.495 2552.705 2914.015 2553.245 ;
        RECT 5.605 2549.475 6.125 2550.015 ;
        RECT 2913.495 2549.475 2914.015 2550.015 ;
        RECT 5.605 2548.725 6.815 2549.475 ;
        RECT 2912.805 2548.725 2914.015 2549.475 ;
        RECT 5.520 2548.555 6.900 2548.725 ;
        RECT 2906.300 2548.555 2906.740 2548.725 ;
        RECT 2912.720 2548.555 2914.100 2548.725 ;
        RECT 5.605 2547.805 6.815 2548.555 ;
        RECT 2906.365 2547.830 2906.655 2548.555 ;
        RECT 2912.805 2547.805 2914.015 2548.555 ;
        RECT 5.605 2547.265 6.125 2547.805 ;
        RECT 2913.495 2547.265 2914.015 2547.805 ;
        RECT 5.605 2544.035 6.125 2544.575 ;
        RECT 2913.495 2544.035 2914.015 2544.575 ;
        RECT 5.605 2543.285 6.815 2544.035 ;
        RECT 2912.805 2543.285 2914.015 2544.035 ;
        RECT 5.520 2543.115 6.900 2543.285 ;
        RECT 2906.300 2543.115 2906.740 2543.285 ;
        RECT 2912.720 2543.115 2914.100 2543.285 ;
        RECT 5.605 2542.365 6.815 2543.115 ;
        RECT 2906.365 2542.390 2906.655 2543.115 ;
        RECT 2912.805 2542.365 2914.015 2543.115 ;
        RECT 5.605 2541.825 6.125 2542.365 ;
        RECT 2913.495 2541.825 2914.015 2542.365 ;
        RECT 5.605 2538.595 6.125 2539.135 ;
        RECT 2913.495 2538.595 2914.015 2539.135 ;
        RECT 5.605 2537.845 6.815 2538.595 ;
        RECT 2912.805 2537.845 2914.015 2538.595 ;
        RECT 5.520 2537.675 6.900 2537.845 ;
        RECT 2906.300 2537.675 2906.740 2537.845 ;
        RECT 2912.720 2537.675 2914.100 2537.845 ;
        RECT 5.605 2536.925 6.815 2537.675 ;
        RECT 2906.365 2536.950 2906.655 2537.675 ;
        RECT 2912.805 2536.925 2914.015 2537.675 ;
        RECT 5.605 2536.385 6.125 2536.925 ;
        RECT 2913.495 2536.385 2914.015 2536.925 ;
        RECT 5.605 2533.155 6.125 2533.695 ;
        RECT 2913.495 2533.155 2914.015 2533.695 ;
        RECT 5.605 2532.405 6.815 2533.155 ;
        RECT 2912.805 2532.405 2914.015 2533.155 ;
        RECT 5.520 2532.235 6.900 2532.405 ;
        RECT 2906.300 2532.235 2906.740 2532.405 ;
        RECT 2912.720 2532.235 2914.100 2532.405 ;
        RECT 5.605 2531.485 6.815 2532.235 ;
        RECT 2906.365 2531.510 2906.655 2532.235 ;
        RECT 2912.805 2531.485 2914.015 2532.235 ;
        RECT 5.605 2530.945 6.125 2531.485 ;
        RECT 2913.495 2530.945 2914.015 2531.485 ;
        RECT 5.605 2527.715 6.125 2528.255 ;
        RECT 2913.495 2527.715 2914.015 2528.255 ;
        RECT 5.605 2526.965 6.815 2527.715 ;
        RECT 2912.805 2526.965 2914.015 2527.715 ;
        RECT 5.520 2526.795 6.900 2526.965 ;
        RECT 2906.300 2526.795 2906.740 2526.965 ;
        RECT 2912.720 2526.795 2914.100 2526.965 ;
        RECT 5.605 2526.045 6.815 2526.795 ;
        RECT 2906.365 2526.070 2906.655 2526.795 ;
        RECT 2912.805 2526.045 2914.015 2526.795 ;
        RECT 5.605 2525.505 6.125 2526.045 ;
        RECT 2913.495 2525.505 2914.015 2526.045 ;
        RECT 5.605 2522.275 6.125 2522.815 ;
        RECT 2913.495 2522.275 2914.015 2522.815 ;
        RECT 5.605 2521.525 6.815 2522.275 ;
        RECT 2912.805 2521.525 2914.015 2522.275 ;
        RECT 5.520 2521.355 6.900 2521.525 ;
        RECT 2906.300 2521.355 2906.740 2521.525 ;
        RECT 2912.720 2521.355 2914.100 2521.525 ;
        RECT 5.605 2520.605 6.815 2521.355 ;
        RECT 2906.365 2520.630 2906.655 2521.355 ;
        RECT 2912.805 2520.605 2914.015 2521.355 ;
        RECT 5.605 2520.065 6.125 2520.605 ;
        RECT 2913.495 2520.065 2914.015 2520.605 ;
        RECT 5.605 2516.835 6.125 2517.375 ;
        RECT 2913.495 2516.835 2914.015 2517.375 ;
        RECT 5.605 2516.085 6.815 2516.835 ;
        RECT 2912.805 2516.085 2914.015 2516.835 ;
        RECT 5.520 2515.915 6.900 2516.085 ;
        RECT 2906.300 2515.915 2906.740 2516.085 ;
        RECT 2912.720 2515.915 2914.100 2516.085 ;
        RECT 5.605 2515.165 6.815 2515.915 ;
        RECT 2906.365 2515.190 2906.655 2515.915 ;
        RECT 2912.805 2515.165 2914.015 2515.915 ;
        RECT 5.605 2514.625 6.125 2515.165 ;
        RECT 2913.495 2514.625 2914.015 2515.165 ;
        RECT 5.605 2511.395 6.125 2511.935 ;
        RECT 2913.495 2511.395 2914.015 2511.935 ;
        RECT 5.605 2510.645 6.815 2511.395 ;
        RECT 2912.805 2510.645 2914.015 2511.395 ;
        RECT 5.520 2510.475 6.900 2510.645 ;
        RECT 2906.300 2510.475 2906.740 2510.645 ;
        RECT 2912.720 2510.475 2914.100 2510.645 ;
        RECT 5.605 2509.725 6.815 2510.475 ;
        RECT 2906.365 2509.750 2906.655 2510.475 ;
        RECT 2912.805 2509.725 2914.015 2510.475 ;
        RECT 5.605 2509.185 6.125 2509.725 ;
        RECT 2913.495 2509.185 2914.015 2509.725 ;
        RECT 5.605 2505.955 6.125 2506.495 ;
        RECT 2913.495 2505.955 2914.015 2506.495 ;
        RECT 5.605 2505.205 6.815 2505.955 ;
        RECT 2912.805 2505.205 2914.015 2505.955 ;
        RECT 5.520 2505.035 6.900 2505.205 ;
        RECT 2906.300 2505.035 2906.740 2505.205 ;
        RECT 2912.720 2505.035 2914.100 2505.205 ;
        RECT 5.605 2504.285 6.815 2505.035 ;
        RECT 2906.365 2504.310 2906.655 2505.035 ;
        RECT 2912.805 2504.285 2914.015 2505.035 ;
        RECT 5.605 2503.745 6.125 2504.285 ;
        RECT 2913.495 2503.745 2914.015 2504.285 ;
        RECT 5.605 2500.515 6.125 2501.055 ;
        RECT 2913.495 2500.515 2914.015 2501.055 ;
        RECT 5.605 2499.765 6.815 2500.515 ;
        RECT 9.515 2499.765 9.855 2500.425 ;
        RECT 2912.805 2499.765 2914.015 2500.515 ;
        RECT 5.520 2499.595 6.900 2499.765 ;
        RECT 8.740 2499.595 10.120 2499.765 ;
        RECT 2906.300 2499.595 2906.740 2499.765 ;
        RECT 2912.720 2499.595 2914.100 2499.765 ;
        RECT 5.605 2498.845 6.815 2499.595 ;
        RECT 2906.365 2498.870 2906.655 2499.595 ;
        RECT 2912.805 2498.845 2914.015 2499.595 ;
        RECT 5.605 2498.305 6.125 2498.845 ;
        RECT 2913.495 2498.305 2914.015 2498.845 ;
        RECT 5.605 2495.075 6.125 2495.615 ;
        RECT 2913.495 2495.075 2914.015 2495.615 ;
        RECT 5.605 2494.325 6.815 2495.075 ;
        RECT 2912.805 2494.325 2914.015 2495.075 ;
        RECT 5.520 2494.155 6.900 2494.325 ;
        RECT 2906.300 2494.155 2906.740 2494.325 ;
        RECT 2912.720 2494.155 2914.100 2494.325 ;
        RECT 5.605 2493.405 6.815 2494.155 ;
        RECT 2906.365 2493.430 2906.655 2494.155 ;
        RECT 2912.805 2493.405 2914.015 2494.155 ;
        RECT 5.605 2492.865 6.125 2493.405 ;
        RECT 2913.495 2492.865 2914.015 2493.405 ;
        RECT 5.605 2489.635 6.125 2490.175 ;
        RECT 2913.495 2489.635 2914.015 2490.175 ;
        RECT 5.605 2488.885 6.815 2489.635 ;
        RECT 2912.805 2488.885 2914.015 2489.635 ;
        RECT 5.520 2488.715 6.900 2488.885 ;
        RECT 2906.300 2488.715 2906.740 2488.885 ;
        RECT 2912.720 2488.715 2914.100 2488.885 ;
        RECT 5.605 2487.965 6.815 2488.715 ;
        RECT 2906.365 2487.990 2906.655 2488.715 ;
        RECT 2912.805 2487.965 2914.015 2488.715 ;
        RECT 5.605 2487.425 6.125 2487.965 ;
        RECT 2913.495 2487.425 2914.015 2487.965 ;
        RECT 5.605 2484.195 6.125 2484.735 ;
        RECT 2913.495 2484.195 2914.015 2484.735 ;
        RECT 5.605 2483.445 6.815 2484.195 ;
        RECT 2912.805 2483.445 2914.015 2484.195 ;
        RECT 5.520 2483.275 6.900 2483.445 ;
        RECT 2906.300 2483.275 2906.740 2483.445 ;
        RECT 2912.720 2483.275 2914.100 2483.445 ;
        RECT 5.605 2482.525 6.815 2483.275 ;
        RECT 2906.365 2482.550 2906.655 2483.275 ;
        RECT 2912.805 2482.525 2914.015 2483.275 ;
        RECT 5.605 2481.985 6.125 2482.525 ;
        RECT 2913.495 2481.985 2914.015 2482.525 ;
        RECT 5.605 2478.755 6.125 2479.295 ;
        RECT 2913.495 2478.755 2914.015 2479.295 ;
        RECT 5.605 2478.005 6.815 2478.755 ;
        RECT 2912.805 2478.005 2914.015 2478.755 ;
        RECT 5.520 2477.835 6.900 2478.005 ;
        RECT 2906.300 2477.835 2906.740 2478.005 ;
        RECT 2912.720 2477.835 2914.100 2478.005 ;
        RECT 5.605 2477.085 6.815 2477.835 ;
        RECT 2906.365 2477.110 2906.655 2477.835 ;
        RECT 2912.805 2477.085 2914.015 2477.835 ;
        RECT 5.605 2476.545 6.125 2477.085 ;
        RECT 2913.495 2476.545 2914.015 2477.085 ;
        RECT 5.605 2473.315 6.125 2473.855 ;
        RECT 2913.495 2473.315 2914.015 2473.855 ;
        RECT 5.605 2472.565 6.815 2473.315 ;
        RECT 2912.805 2472.565 2914.015 2473.315 ;
        RECT 5.520 2472.395 6.900 2472.565 ;
        RECT 2906.300 2472.395 2906.740 2472.565 ;
        RECT 2912.720 2472.395 2914.100 2472.565 ;
        RECT 5.605 2471.645 6.815 2472.395 ;
        RECT 2906.365 2471.670 2906.655 2472.395 ;
        RECT 2912.805 2471.645 2914.015 2472.395 ;
        RECT 5.605 2471.105 6.125 2471.645 ;
        RECT 2913.495 2471.105 2914.015 2471.645 ;
        RECT 5.605 2467.875 6.125 2468.415 ;
        RECT 2913.495 2467.875 2914.015 2468.415 ;
        RECT 5.605 2467.125 6.815 2467.875 ;
        RECT 2912.805 2467.125 2914.015 2467.875 ;
        RECT 5.520 2466.955 6.900 2467.125 ;
        RECT 2906.300 2466.955 2906.740 2467.125 ;
        RECT 2912.720 2466.955 2914.100 2467.125 ;
        RECT 5.605 2466.205 6.815 2466.955 ;
        RECT 2906.365 2466.230 2906.655 2466.955 ;
        RECT 2912.805 2466.205 2914.015 2466.955 ;
        RECT 5.605 2465.665 6.125 2466.205 ;
        RECT 2913.495 2465.665 2914.015 2466.205 ;
        RECT 5.605 2462.435 6.125 2462.975 ;
        RECT 2913.495 2462.435 2914.015 2462.975 ;
        RECT 5.605 2461.685 6.815 2462.435 ;
        RECT 2909.815 2461.685 2910.155 2462.345 ;
        RECT 2912.805 2461.685 2914.015 2462.435 ;
        RECT 5.520 2461.515 6.900 2461.685 ;
        RECT 2906.300 2461.515 2906.740 2461.685 ;
        RECT 2909.040 2461.515 2910.420 2461.685 ;
        RECT 2912.720 2461.515 2914.100 2461.685 ;
        RECT 5.605 2460.765 6.815 2461.515 ;
        RECT 2906.365 2460.790 2906.655 2461.515 ;
        RECT 2912.805 2460.765 2914.015 2461.515 ;
        RECT 5.605 2460.225 6.125 2460.765 ;
        RECT 2913.495 2460.225 2914.015 2460.765 ;
        RECT 5.605 2456.995 6.125 2457.535 ;
        RECT 2913.495 2456.995 2914.015 2457.535 ;
        RECT 5.605 2456.245 6.815 2456.995 ;
        RECT 2912.805 2456.245 2914.015 2456.995 ;
        RECT 5.520 2456.075 6.900 2456.245 ;
        RECT 2906.300 2456.075 2906.740 2456.245 ;
        RECT 2912.720 2456.075 2914.100 2456.245 ;
        RECT 5.605 2455.325 6.815 2456.075 ;
        RECT 2906.365 2455.350 2906.655 2456.075 ;
        RECT 2912.805 2455.325 2914.015 2456.075 ;
        RECT 5.605 2454.785 6.125 2455.325 ;
        RECT 2913.495 2454.785 2914.015 2455.325 ;
        RECT 5.605 2451.555 6.125 2452.095 ;
        RECT 2913.495 2451.555 2914.015 2452.095 ;
        RECT 5.605 2450.805 6.815 2451.555 ;
        RECT 2912.805 2450.805 2914.015 2451.555 ;
        RECT 5.520 2450.635 6.900 2450.805 ;
        RECT 2906.300 2450.635 2906.740 2450.805 ;
        RECT 2912.720 2450.635 2914.100 2450.805 ;
        RECT 5.605 2449.885 6.815 2450.635 ;
        RECT 2906.365 2449.910 2906.655 2450.635 ;
        RECT 2912.805 2449.885 2914.015 2450.635 ;
        RECT 5.605 2449.345 6.125 2449.885 ;
        RECT 2913.495 2449.345 2914.015 2449.885 ;
        RECT 5.605 2446.115 6.125 2446.655 ;
        RECT 2913.495 2446.115 2914.015 2446.655 ;
        RECT 5.605 2445.365 6.815 2446.115 ;
        RECT 2912.805 2445.365 2914.015 2446.115 ;
        RECT 5.520 2445.195 6.900 2445.365 ;
        RECT 2906.300 2445.195 2906.740 2445.365 ;
        RECT 2912.720 2445.195 2914.100 2445.365 ;
        RECT 5.605 2444.445 6.815 2445.195 ;
        RECT 2906.365 2444.470 2906.655 2445.195 ;
        RECT 2912.805 2444.445 2914.015 2445.195 ;
        RECT 5.605 2443.905 6.125 2444.445 ;
        RECT 2913.495 2443.905 2914.015 2444.445 ;
        RECT 5.605 2440.675 6.125 2441.215 ;
        RECT 2913.495 2440.675 2914.015 2441.215 ;
        RECT 5.605 2439.925 6.815 2440.675 ;
        RECT 2912.805 2439.925 2914.015 2440.675 ;
        RECT 5.520 2439.755 6.900 2439.925 ;
        RECT 2906.300 2439.755 2906.740 2439.925 ;
        RECT 2912.720 2439.755 2914.100 2439.925 ;
        RECT 5.605 2439.005 6.815 2439.755 ;
        RECT 2906.365 2439.030 2906.655 2439.755 ;
        RECT 2912.805 2439.005 2914.015 2439.755 ;
        RECT 5.605 2438.465 6.125 2439.005 ;
        RECT 2913.495 2438.465 2914.015 2439.005 ;
        RECT 5.605 2435.235 6.125 2435.775 ;
        RECT 2913.495 2435.235 2914.015 2435.775 ;
        RECT 5.605 2434.485 6.815 2435.235 ;
        RECT 2912.805 2434.485 2914.015 2435.235 ;
        RECT 5.520 2434.315 6.900 2434.485 ;
        RECT 2906.300 2434.315 2906.740 2434.485 ;
        RECT 2909.040 2434.315 2910.420 2434.485 ;
        RECT 2912.720 2434.315 2914.100 2434.485 ;
        RECT 5.605 2433.565 6.815 2434.315 ;
        RECT 2906.365 2433.590 2906.655 2434.315 ;
        RECT 2909.815 2433.655 2910.155 2434.315 ;
        RECT 2912.805 2433.565 2914.015 2434.315 ;
        RECT 5.605 2433.025 6.125 2433.565 ;
        RECT 2913.495 2433.025 2914.015 2433.565 ;
        RECT 5.605 2429.795 6.125 2430.335 ;
        RECT 2913.495 2429.795 2914.015 2430.335 ;
        RECT 5.605 2429.045 6.815 2429.795 ;
        RECT 2912.805 2429.045 2914.015 2429.795 ;
        RECT 5.520 2428.875 6.900 2429.045 ;
        RECT 2906.300 2428.875 2906.740 2429.045 ;
        RECT 2912.720 2428.875 2914.100 2429.045 ;
        RECT 5.605 2428.125 6.815 2428.875 ;
        RECT 2906.365 2428.150 2906.655 2428.875 ;
        RECT 2912.805 2428.125 2914.015 2428.875 ;
        RECT 5.605 2427.585 6.125 2428.125 ;
        RECT 2913.495 2427.585 2914.015 2428.125 ;
        RECT 5.605 2424.355 6.125 2424.895 ;
        RECT 2913.495 2424.355 2914.015 2424.895 ;
        RECT 5.605 2423.605 6.815 2424.355 ;
        RECT 2912.805 2423.605 2914.015 2424.355 ;
        RECT 5.520 2423.435 6.900 2423.605 ;
        RECT 2906.300 2423.435 2906.740 2423.605 ;
        RECT 2912.720 2423.435 2914.100 2423.605 ;
        RECT 5.605 2422.685 6.815 2423.435 ;
        RECT 2906.365 2422.710 2906.655 2423.435 ;
        RECT 2912.805 2422.685 2914.015 2423.435 ;
        RECT 5.605 2422.145 6.125 2422.685 ;
        RECT 2913.495 2422.145 2914.015 2422.685 ;
        RECT 5.605 2418.915 6.125 2419.455 ;
        RECT 2913.495 2418.915 2914.015 2419.455 ;
        RECT 5.605 2418.165 6.815 2418.915 ;
        RECT 2912.805 2418.165 2914.015 2418.915 ;
        RECT 5.520 2417.995 6.900 2418.165 ;
        RECT 2906.300 2417.995 2906.740 2418.165 ;
        RECT 2912.720 2417.995 2914.100 2418.165 ;
        RECT 5.605 2417.245 6.815 2417.995 ;
        RECT 2906.365 2417.270 2906.655 2417.995 ;
        RECT 2912.805 2417.245 2914.015 2417.995 ;
        RECT 5.605 2416.705 6.125 2417.245 ;
        RECT 2913.495 2416.705 2914.015 2417.245 ;
        RECT 5.605 2413.475 6.125 2414.015 ;
        RECT 2913.495 2413.475 2914.015 2414.015 ;
        RECT 5.605 2412.725 6.815 2413.475 ;
        RECT 2912.805 2412.725 2914.015 2413.475 ;
        RECT 5.520 2412.555 6.900 2412.725 ;
        RECT 2906.300 2412.555 2906.740 2412.725 ;
        RECT 2912.720 2412.555 2914.100 2412.725 ;
        RECT 5.605 2411.805 6.815 2412.555 ;
        RECT 2906.365 2411.830 2906.655 2412.555 ;
        RECT 2912.805 2411.805 2914.015 2412.555 ;
        RECT 5.605 2411.265 6.125 2411.805 ;
        RECT 2913.495 2411.265 2914.015 2411.805 ;
        RECT 5.605 2408.035 6.125 2408.575 ;
        RECT 2913.495 2408.035 2914.015 2408.575 ;
        RECT 5.605 2407.285 6.815 2408.035 ;
        RECT 2912.805 2407.285 2914.015 2408.035 ;
        RECT 5.520 2407.115 6.900 2407.285 ;
        RECT 2906.300 2407.115 2906.740 2407.285 ;
        RECT 2912.720 2407.115 2914.100 2407.285 ;
        RECT 5.605 2406.365 6.815 2407.115 ;
        RECT 2906.365 2406.390 2906.655 2407.115 ;
        RECT 2912.805 2406.365 2914.015 2407.115 ;
        RECT 5.605 2405.825 6.125 2406.365 ;
        RECT 2913.495 2405.825 2914.015 2406.365 ;
        RECT 5.605 2402.595 6.125 2403.135 ;
        RECT 2913.495 2402.595 2914.015 2403.135 ;
        RECT 5.605 2401.845 6.815 2402.595 ;
        RECT 2912.805 2401.845 2914.015 2402.595 ;
        RECT 5.520 2401.675 6.900 2401.845 ;
        RECT 2906.300 2401.675 2906.740 2401.845 ;
        RECT 2912.720 2401.675 2914.100 2401.845 ;
        RECT 5.605 2400.925 6.815 2401.675 ;
        RECT 2906.365 2400.950 2906.655 2401.675 ;
        RECT 2912.805 2400.925 2914.015 2401.675 ;
        RECT 5.605 2400.385 6.125 2400.925 ;
        RECT 2913.495 2400.385 2914.015 2400.925 ;
        RECT 5.605 2397.155 6.125 2397.695 ;
        RECT 2913.495 2397.155 2914.015 2397.695 ;
        RECT 5.605 2396.405 6.815 2397.155 ;
        RECT 2912.805 2396.405 2914.015 2397.155 ;
        RECT 5.520 2396.235 6.900 2396.405 ;
        RECT 2906.300 2396.235 2906.740 2396.405 ;
        RECT 2912.720 2396.235 2914.100 2396.405 ;
        RECT 5.605 2395.485 6.815 2396.235 ;
        RECT 2906.365 2395.510 2906.655 2396.235 ;
        RECT 2912.805 2395.485 2914.015 2396.235 ;
        RECT 5.605 2394.945 6.125 2395.485 ;
        RECT 2913.495 2394.945 2914.015 2395.485 ;
        RECT 5.605 2391.715 6.125 2392.255 ;
        RECT 2913.495 2391.715 2914.015 2392.255 ;
        RECT 5.605 2390.965 6.815 2391.715 ;
        RECT 2912.805 2390.965 2914.015 2391.715 ;
        RECT 5.520 2390.795 6.900 2390.965 ;
        RECT 2906.300 2390.795 2906.740 2390.965 ;
        RECT 2912.720 2390.795 2914.100 2390.965 ;
        RECT 5.605 2390.045 6.815 2390.795 ;
        RECT 2906.365 2390.070 2906.655 2390.795 ;
        RECT 2912.805 2390.045 2914.015 2390.795 ;
        RECT 5.605 2389.505 6.125 2390.045 ;
        RECT 2913.495 2389.505 2914.015 2390.045 ;
        RECT 5.605 2386.275 6.125 2386.815 ;
        RECT 2913.495 2386.275 2914.015 2386.815 ;
        RECT 5.605 2385.525 6.815 2386.275 ;
        RECT 2909.815 2385.525 2910.155 2386.185 ;
        RECT 2912.805 2385.525 2914.015 2386.275 ;
        RECT 5.520 2385.355 6.900 2385.525 ;
        RECT 2906.300 2385.355 2906.740 2385.525 ;
        RECT 2909.040 2385.355 2910.420 2385.525 ;
        RECT 2912.720 2385.355 2914.100 2385.525 ;
        RECT 5.605 2384.605 6.815 2385.355 ;
        RECT 2906.365 2384.630 2906.655 2385.355 ;
        RECT 2912.805 2384.605 2914.015 2385.355 ;
        RECT 5.605 2384.065 6.125 2384.605 ;
        RECT 2913.495 2384.065 2914.015 2384.605 ;
        RECT 5.605 2380.835 6.125 2381.375 ;
        RECT 2913.495 2380.835 2914.015 2381.375 ;
        RECT 5.605 2380.085 6.815 2380.835 ;
        RECT 9.515 2380.085 9.855 2380.745 ;
        RECT 2912.805 2380.085 2914.015 2380.835 ;
        RECT 5.520 2379.915 6.900 2380.085 ;
        RECT 8.740 2379.915 10.120 2380.085 ;
        RECT 2906.300 2379.915 2906.740 2380.085 ;
        RECT 2912.720 2379.915 2914.100 2380.085 ;
        RECT 5.605 2379.165 6.815 2379.915 ;
        RECT 2906.365 2379.190 2906.655 2379.915 ;
        RECT 2912.805 2379.165 2914.015 2379.915 ;
        RECT 5.605 2378.625 6.125 2379.165 ;
        RECT 2913.495 2378.625 2914.015 2379.165 ;
        RECT 5.605 2375.395 6.125 2375.935 ;
        RECT 2913.495 2375.395 2914.015 2375.935 ;
        RECT 5.605 2374.645 6.815 2375.395 ;
        RECT 2912.805 2374.645 2914.015 2375.395 ;
        RECT 5.520 2374.475 6.900 2374.645 ;
        RECT 2906.300 2374.475 2906.740 2374.645 ;
        RECT 2912.720 2374.475 2914.100 2374.645 ;
        RECT 5.605 2373.725 6.815 2374.475 ;
        RECT 2906.365 2373.750 2906.655 2374.475 ;
        RECT 2912.805 2373.725 2914.015 2374.475 ;
        RECT 5.605 2373.185 6.125 2373.725 ;
        RECT 2913.495 2373.185 2914.015 2373.725 ;
        RECT 5.605 2369.955 6.125 2370.495 ;
        RECT 2913.495 2369.955 2914.015 2370.495 ;
        RECT 5.605 2369.205 6.815 2369.955 ;
        RECT 2912.805 2369.205 2914.015 2369.955 ;
        RECT 5.520 2369.035 6.900 2369.205 ;
        RECT 2906.300 2369.035 2906.740 2369.205 ;
        RECT 2912.720 2369.035 2914.100 2369.205 ;
        RECT 5.605 2368.285 6.815 2369.035 ;
        RECT 2906.365 2368.310 2906.655 2369.035 ;
        RECT 2912.805 2368.285 2914.015 2369.035 ;
        RECT 5.605 2367.745 6.125 2368.285 ;
        RECT 2913.495 2367.745 2914.015 2368.285 ;
        RECT 5.605 2364.515 6.125 2365.055 ;
        RECT 2913.495 2364.515 2914.015 2365.055 ;
        RECT 5.605 2363.765 6.815 2364.515 ;
        RECT 2912.805 2363.765 2914.015 2364.515 ;
        RECT 5.520 2363.595 6.900 2363.765 ;
        RECT 2906.300 2363.595 2906.740 2363.765 ;
        RECT 2912.720 2363.595 2914.100 2363.765 ;
        RECT 5.605 2362.845 6.815 2363.595 ;
        RECT 2906.365 2362.870 2906.655 2363.595 ;
        RECT 2912.805 2362.845 2914.015 2363.595 ;
        RECT 5.605 2362.305 6.125 2362.845 ;
        RECT 2913.495 2362.305 2914.015 2362.845 ;
        RECT 5.605 2359.075 6.125 2359.615 ;
        RECT 2913.495 2359.075 2914.015 2359.615 ;
        RECT 5.605 2358.325 6.815 2359.075 ;
        RECT 2912.805 2358.325 2914.015 2359.075 ;
        RECT 5.520 2358.155 6.900 2358.325 ;
        RECT 2906.300 2358.155 2906.740 2358.325 ;
        RECT 2912.720 2358.155 2914.100 2358.325 ;
        RECT 5.605 2357.405 6.815 2358.155 ;
        RECT 2906.365 2357.430 2906.655 2358.155 ;
        RECT 2912.805 2357.405 2914.015 2358.155 ;
        RECT 5.605 2356.865 6.125 2357.405 ;
        RECT 2913.495 2356.865 2914.015 2357.405 ;
        RECT 5.605 2353.635 6.125 2354.175 ;
        RECT 2913.495 2353.635 2914.015 2354.175 ;
        RECT 5.605 2352.885 6.815 2353.635 ;
        RECT 2912.805 2352.885 2914.015 2353.635 ;
        RECT 5.520 2352.715 6.900 2352.885 ;
        RECT 2906.300 2352.715 2906.740 2352.885 ;
        RECT 2912.720 2352.715 2914.100 2352.885 ;
        RECT 5.605 2351.965 6.815 2352.715 ;
        RECT 2906.365 2351.990 2906.655 2352.715 ;
        RECT 2912.805 2351.965 2914.015 2352.715 ;
        RECT 5.605 2351.425 6.125 2351.965 ;
        RECT 2913.495 2351.425 2914.015 2351.965 ;
        RECT 5.605 2348.195 6.125 2348.735 ;
        RECT 2913.495 2348.195 2914.015 2348.735 ;
        RECT 5.605 2347.445 6.815 2348.195 ;
        RECT 2912.805 2347.445 2914.015 2348.195 ;
        RECT 5.520 2347.275 6.900 2347.445 ;
        RECT 2906.300 2347.275 2906.740 2347.445 ;
        RECT 2912.720 2347.275 2914.100 2347.445 ;
        RECT 5.605 2346.525 6.815 2347.275 ;
        RECT 2906.365 2346.550 2906.655 2347.275 ;
        RECT 2912.805 2346.525 2914.015 2347.275 ;
        RECT 5.605 2345.985 6.125 2346.525 ;
        RECT 2913.495 2345.985 2914.015 2346.525 ;
        RECT 5.605 2342.755 6.125 2343.295 ;
        RECT 2913.495 2342.755 2914.015 2343.295 ;
        RECT 5.605 2342.005 6.815 2342.755 ;
        RECT 2912.805 2342.005 2914.015 2342.755 ;
        RECT 5.520 2341.835 6.900 2342.005 ;
        RECT 2906.300 2341.835 2906.740 2342.005 ;
        RECT 2912.720 2341.835 2914.100 2342.005 ;
        RECT 5.605 2341.085 6.815 2341.835 ;
        RECT 2906.365 2341.110 2906.655 2341.835 ;
        RECT 2912.805 2341.085 2914.015 2341.835 ;
        RECT 5.605 2340.545 6.125 2341.085 ;
        RECT 2913.495 2340.545 2914.015 2341.085 ;
        RECT 5.605 2337.315 6.125 2337.855 ;
        RECT 2913.495 2337.315 2914.015 2337.855 ;
        RECT 5.605 2336.565 6.815 2337.315 ;
        RECT 2912.805 2336.565 2914.015 2337.315 ;
        RECT 5.520 2336.395 6.900 2336.565 ;
        RECT 2906.300 2336.395 2906.740 2336.565 ;
        RECT 2912.720 2336.395 2914.100 2336.565 ;
        RECT 5.605 2335.645 6.815 2336.395 ;
        RECT 2906.365 2335.670 2906.655 2336.395 ;
        RECT 2912.805 2335.645 2914.015 2336.395 ;
        RECT 5.605 2335.105 6.125 2335.645 ;
        RECT 2913.495 2335.105 2914.015 2335.645 ;
        RECT 5.605 2331.875 6.125 2332.415 ;
        RECT 2913.495 2331.875 2914.015 2332.415 ;
        RECT 5.605 2331.125 6.815 2331.875 ;
        RECT 2912.805 2331.125 2914.015 2331.875 ;
        RECT 5.520 2330.955 6.900 2331.125 ;
        RECT 2906.300 2330.955 2906.740 2331.125 ;
        RECT 2912.720 2330.955 2914.100 2331.125 ;
        RECT 5.605 2330.205 6.815 2330.955 ;
        RECT 2906.365 2330.230 2906.655 2330.955 ;
        RECT 2912.805 2330.205 2914.015 2330.955 ;
        RECT 5.605 2329.665 6.125 2330.205 ;
        RECT 2913.495 2329.665 2914.015 2330.205 ;
        RECT 5.605 2326.435 6.125 2326.975 ;
        RECT 2913.495 2326.435 2914.015 2326.975 ;
        RECT 5.605 2325.685 6.815 2326.435 ;
        RECT 2912.805 2325.685 2914.015 2326.435 ;
        RECT 5.520 2325.515 6.900 2325.685 ;
        RECT 2906.300 2325.515 2906.740 2325.685 ;
        RECT 2912.720 2325.515 2914.100 2325.685 ;
        RECT 5.605 2324.765 6.815 2325.515 ;
        RECT 2906.365 2324.790 2906.655 2325.515 ;
        RECT 2912.805 2324.765 2914.015 2325.515 ;
        RECT 5.605 2324.225 6.125 2324.765 ;
        RECT 2913.495 2324.225 2914.015 2324.765 ;
        RECT 5.605 2320.995 6.125 2321.535 ;
        RECT 2913.495 2320.995 2914.015 2321.535 ;
        RECT 5.605 2320.245 6.815 2320.995 ;
        RECT 2912.805 2320.245 2914.015 2320.995 ;
        RECT 5.520 2320.075 6.900 2320.245 ;
        RECT 2906.300 2320.075 2906.740 2320.245 ;
        RECT 2912.720 2320.075 2914.100 2320.245 ;
        RECT 5.605 2319.325 6.815 2320.075 ;
        RECT 2906.365 2319.350 2906.655 2320.075 ;
        RECT 2912.805 2319.325 2914.015 2320.075 ;
        RECT 5.605 2318.785 6.125 2319.325 ;
        RECT 2913.495 2318.785 2914.015 2319.325 ;
        RECT 5.605 2315.555 6.125 2316.095 ;
        RECT 2913.495 2315.555 2914.015 2316.095 ;
        RECT 5.605 2314.805 6.815 2315.555 ;
        RECT 2912.805 2314.805 2914.015 2315.555 ;
        RECT 5.520 2314.635 6.900 2314.805 ;
        RECT 2906.300 2314.635 2906.740 2314.805 ;
        RECT 2912.720 2314.635 2914.100 2314.805 ;
        RECT 5.605 2313.885 6.815 2314.635 ;
        RECT 2906.365 2313.910 2906.655 2314.635 ;
        RECT 2912.805 2313.885 2914.015 2314.635 ;
        RECT 5.605 2313.345 6.125 2313.885 ;
        RECT 2913.495 2313.345 2914.015 2313.885 ;
        RECT 5.605 2310.115 6.125 2310.655 ;
        RECT 2913.495 2310.115 2914.015 2310.655 ;
        RECT 5.605 2309.365 6.815 2310.115 ;
        RECT 2912.805 2309.365 2914.015 2310.115 ;
        RECT 5.520 2309.195 6.900 2309.365 ;
        RECT 2906.300 2309.195 2906.740 2309.365 ;
        RECT 2912.720 2309.195 2914.100 2309.365 ;
        RECT 5.605 2308.445 6.815 2309.195 ;
        RECT 2906.365 2308.470 2906.655 2309.195 ;
        RECT 2912.805 2308.445 2914.015 2309.195 ;
        RECT 5.605 2307.905 6.125 2308.445 ;
        RECT 2913.495 2307.905 2914.015 2308.445 ;
        RECT 5.605 2304.675 6.125 2305.215 ;
        RECT 2913.495 2304.675 2914.015 2305.215 ;
        RECT 5.605 2303.925 6.815 2304.675 ;
        RECT 2912.805 2303.925 2914.015 2304.675 ;
        RECT 5.520 2303.755 6.900 2303.925 ;
        RECT 2906.300 2303.755 2906.740 2303.925 ;
        RECT 2912.720 2303.755 2914.100 2303.925 ;
        RECT 5.605 2303.005 6.815 2303.755 ;
        RECT 2906.365 2303.030 2906.655 2303.755 ;
        RECT 2912.805 2303.005 2914.015 2303.755 ;
        RECT 5.605 2302.465 6.125 2303.005 ;
        RECT 2913.495 2302.465 2914.015 2303.005 ;
        RECT 5.605 2299.235 6.125 2299.775 ;
        RECT 2913.495 2299.235 2914.015 2299.775 ;
        RECT 5.605 2298.485 6.815 2299.235 ;
        RECT 2912.805 2298.485 2914.015 2299.235 ;
        RECT 5.520 2298.315 6.900 2298.485 ;
        RECT 2906.300 2298.315 2906.740 2298.485 ;
        RECT 2912.720 2298.315 2914.100 2298.485 ;
        RECT 5.605 2297.565 6.815 2298.315 ;
        RECT 2906.365 2297.590 2906.655 2298.315 ;
        RECT 2912.805 2297.565 2914.015 2298.315 ;
        RECT 5.605 2297.025 6.125 2297.565 ;
        RECT 2913.495 2297.025 2914.015 2297.565 ;
        RECT 5.605 2293.795 6.125 2294.335 ;
        RECT 2913.495 2293.795 2914.015 2294.335 ;
        RECT 5.605 2293.045 6.815 2293.795 ;
        RECT 2912.805 2293.045 2914.015 2293.795 ;
        RECT 5.520 2292.875 6.900 2293.045 ;
        RECT 2906.300 2292.875 2906.740 2293.045 ;
        RECT 2912.720 2292.875 2914.100 2293.045 ;
        RECT 5.605 2292.125 6.815 2292.875 ;
        RECT 2906.365 2292.150 2906.655 2292.875 ;
        RECT 2912.805 2292.125 2914.015 2292.875 ;
        RECT 5.605 2291.585 6.125 2292.125 ;
        RECT 2913.495 2291.585 2914.015 2292.125 ;
        RECT 5.605 2288.355 6.125 2288.895 ;
        RECT 2913.495 2288.355 2914.015 2288.895 ;
        RECT 5.605 2287.605 6.815 2288.355 ;
        RECT 2912.805 2287.605 2914.015 2288.355 ;
        RECT 5.520 2287.435 6.900 2287.605 ;
        RECT 2906.300 2287.435 2906.740 2287.605 ;
        RECT 2912.720 2287.435 2914.100 2287.605 ;
        RECT 5.605 2286.685 6.815 2287.435 ;
        RECT 2906.365 2286.710 2906.655 2287.435 ;
        RECT 2912.805 2286.685 2914.015 2287.435 ;
        RECT 5.605 2286.145 6.125 2286.685 ;
        RECT 2913.495 2286.145 2914.015 2286.685 ;
        RECT 5.605 2282.915 6.125 2283.455 ;
        RECT 2913.495 2282.915 2914.015 2283.455 ;
        RECT 5.605 2282.165 6.815 2282.915 ;
        RECT 2912.805 2282.165 2914.015 2282.915 ;
        RECT 5.520 2281.995 6.900 2282.165 ;
        RECT 2906.300 2281.995 2906.740 2282.165 ;
        RECT 2912.720 2281.995 2914.100 2282.165 ;
        RECT 5.605 2281.245 6.815 2281.995 ;
        RECT 2906.365 2281.270 2906.655 2281.995 ;
        RECT 2912.805 2281.245 2914.015 2281.995 ;
        RECT 5.605 2280.705 6.125 2281.245 ;
        RECT 2913.495 2280.705 2914.015 2281.245 ;
        RECT 5.605 2277.475 6.125 2278.015 ;
        RECT 2913.495 2277.475 2914.015 2278.015 ;
        RECT 5.605 2276.725 6.815 2277.475 ;
        RECT 2912.805 2276.725 2914.015 2277.475 ;
        RECT 5.520 2276.555 6.900 2276.725 ;
        RECT 2906.300 2276.555 2906.740 2276.725 ;
        RECT 2912.720 2276.555 2914.100 2276.725 ;
        RECT 5.605 2275.805 6.815 2276.555 ;
        RECT 2906.365 2275.830 2906.655 2276.555 ;
        RECT 2912.805 2275.805 2914.015 2276.555 ;
        RECT 5.605 2275.265 6.125 2275.805 ;
        RECT 2913.495 2275.265 2914.015 2275.805 ;
        RECT 5.605 2272.035 6.125 2272.575 ;
        RECT 2913.495 2272.035 2914.015 2272.575 ;
        RECT 5.605 2271.285 6.815 2272.035 ;
        RECT 2912.805 2271.285 2914.015 2272.035 ;
        RECT 5.520 2271.115 6.900 2271.285 ;
        RECT 2906.300 2271.115 2906.740 2271.285 ;
        RECT 2912.720 2271.115 2914.100 2271.285 ;
        RECT 5.605 2270.365 6.815 2271.115 ;
        RECT 2906.365 2270.390 2906.655 2271.115 ;
        RECT 2912.805 2270.365 2914.015 2271.115 ;
        RECT 5.605 2269.825 6.125 2270.365 ;
        RECT 2913.495 2269.825 2914.015 2270.365 ;
        RECT 5.605 2266.595 6.125 2267.135 ;
        RECT 2913.495 2266.595 2914.015 2267.135 ;
        RECT 5.605 2265.845 6.815 2266.595 ;
        RECT 2912.805 2265.845 2914.015 2266.595 ;
        RECT 5.520 2265.675 6.900 2265.845 ;
        RECT 2906.300 2265.675 2906.740 2265.845 ;
        RECT 2909.040 2265.675 2910.420 2265.845 ;
        RECT 2912.720 2265.675 2914.100 2265.845 ;
        RECT 5.605 2264.925 6.815 2265.675 ;
        RECT 2906.365 2264.950 2906.655 2265.675 ;
        RECT 2909.815 2265.015 2910.155 2265.675 ;
        RECT 2912.805 2264.925 2914.015 2265.675 ;
        RECT 5.605 2264.385 6.125 2264.925 ;
        RECT 2913.495 2264.385 2914.015 2264.925 ;
        RECT 5.605 2261.155 6.125 2261.695 ;
        RECT 2913.495 2261.155 2914.015 2261.695 ;
        RECT 5.605 2260.405 6.815 2261.155 ;
        RECT 2912.805 2260.405 2914.015 2261.155 ;
        RECT 5.520 2260.235 6.900 2260.405 ;
        RECT 2906.300 2260.235 2906.740 2260.405 ;
        RECT 2912.720 2260.235 2914.100 2260.405 ;
        RECT 5.605 2259.485 6.815 2260.235 ;
        RECT 2906.365 2259.510 2906.655 2260.235 ;
        RECT 2912.805 2259.485 2914.015 2260.235 ;
        RECT 5.605 2258.945 6.125 2259.485 ;
        RECT 2913.495 2258.945 2914.015 2259.485 ;
        RECT 5.605 2255.715 6.125 2256.255 ;
        RECT 2913.495 2255.715 2914.015 2256.255 ;
        RECT 5.605 2254.965 6.815 2255.715 ;
        RECT 2912.805 2254.965 2914.015 2255.715 ;
        RECT 5.520 2254.795 6.900 2254.965 ;
        RECT 2906.300 2254.795 2906.740 2254.965 ;
        RECT 2912.720 2254.795 2914.100 2254.965 ;
        RECT 5.605 2254.045 6.815 2254.795 ;
        RECT 2906.365 2254.070 2906.655 2254.795 ;
        RECT 2912.805 2254.045 2914.015 2254.795 ;
        RECT 5.605 2253.505 6.125 2254.045 ;
        RECT 2913.495 2253.505 2914.015 2254.045 ;
        RECT 5.605 2250.275 6.125 2250.815 ;
        RECT 2913.495 2250.275 2914.015 2250.815 ;
        RECT 5.605 2249.525 6.815 2250.275 ;
        RECT 2912.805 2249.525 2914.015 2250.275 ;
        RECT 5.520 2249.355 6.900 2249.525 ;
        RECT 2906.300 2249.355 2906.740 2249.525 ;
        RECT 2912.720 2249.355 2914.100 2249.525 ;
        RECT 5.605 2248.605 6.815 2249.355 ;
        RECT 2906.365 2248.630 2906.655 2249.355 ;
        RECT 2912.805 2248.605 2914.015 2249.355 ;
        RECT 5.605 2248.065 6.125 2248.605 ;
        RECT 2913.495 2248.065 2914.015 2248.605 ;
        RECT 5.605 2244.835 6.125 2245.375 ;
        RECT 2913.495 2244.835 2914.015 2245.375 ;
        RECT 5.605 2244.085 6.815 2244.835 ;
        RECT 2912.805 2244.085 2914.015 2244.835 ;
        RECT 5.520 2243.915 6.900 2244.085 ;
        RECT 2906.300 2243.915 2906.740 2244.085 ;
        RECT 2912.720 2243.915 2914.100 2244.085 ;
        RECT 5.605 2243.165 6.815 2243.915 ;
        RECT 2906.365 2243.190 2906.655 2243.915 ;
        RECT 2912.805 2243.165 2914.015 2243.915 ;
        RECT 5.605 2242.625 6.125 2243.165 ;
        RECT 2913.495 2242.625 2914.015 2243.165 ;
        RECT 5.605 2239.395 6.125 2239.935 ;
        RECT 2913.495 2239.395 2914.015 2239.935 ;
        RECT 5.605 2238.645 6.815 2239.395 ;
        RECT 2912.805 2238.645 2914.015 2239.395 ;
        RECT 5.520 2238.475 6.900 2238.645 ;
        RECT 2906.300 2238.475 2906.740 2238.645 ;
        RECT 2912.720 2238.475 2914.100 2238.645 ;
        RECT 5.605 2237.725 6.815 2238.475 ;
        RECT 2906.365 2237.750 2906.655 2238.475 ;
        RECT 2912.805 2237.725 2914.015 2238.475 ;
        RECT 5.605 2237.185 6.125 2237.725 ;
        RECT 2913.495 2237.185 2914.015 2237.725 ;
        RECT 5.605 2233.955 6.125 2234.495 ;
        RECT 2913.495 2233.955 2914.015 2234.495 ;
        RECT 5.605 2233.205 6.815 2233.955 ;
        RECT 2912.805 2233.205 2914.015 2233.955 ;
        RECT 5.520 2233.035 6.900 2233.205 ;
        RECT 2906.300 2233.035 2906.740 2233.205 ;
        RECT 2912.720 2233.035 2914.100 2233.205 ;
        RECT 5.605 2232.285 6.815 2233.035 ;
        RECT 2906.365 2232.310 2906.655 2233.035 ;
        RECT 2912.805 2232.285 2914.015 2233.035 ;
        RECT 5.605 2231.745 6.125 2232.285 ;
        RECT 2913.495 2231.745 2914.015 2232.285 ;
        RECT 5.605 2228.515 6.125 2229.055 ;
        RECT 2913.495 2228.515 2914.015 2229.055 ;
        RECT 5.605 2227.765 6.815 2228.515 ;
        RECT 2912.805 2227.765 2914.015 2228.515 ;
        RECT 5.520 2227.595 6.900 2227.765 ;
        RECT 2906.300 2227.595 2906.740 2227.765 ;
        RECT 2912.720 2227.595 2914.100 2227.765 ;
        RECT 5.605 2226.845 6.815 2227.595 ;
        RECT 2906.365 2226.870 2906.655 2227.595 ;
        RECT 2912.805 2226.845 2914.015 2227.595 ;
        RECT 5.605 2226.305 6.125 2226.845 ;
        RECT 2913.495 2226.305 2914.015 2226.845 ;
        RECT 5.605 2223.075 6.125 2223.615 ;
        RECT 2913.495 2223.075 2914.015 2223.615 ;
        RECT 5.605 2222.325 6.815 2223.075 ;
        RECT 2912.805 2222.325 2914.015 2223.075 ;
        RECT 5.520 2222.155 6.900 2222.325 ;
        RECT 2906.300 2222.155 2906.740 2222.325 ;
        RECT 2912.720 2222.155 2914.100 2222.325 ;
        RECT 5.605 2221.405 6.815 2222.155 ;
        RECT 2906.365 2221.430 2906.655 2222.155 ;
        RECT 2912.805 2221.405 2914.015 2222.155 ;
        RECT 5.605 2220.865 6.125 2221.405 ;
        RECT 2913.495 2220.865 2914.015 2221.405 ;
        RECT 5.605 2217.635 6.125 2218.175 ;
        RECT 2913.495 2217.635 2914.015 2218.175 ;
        RECT 5.605 2216.885 6.815 2217.635 ;
        RECT 2912.805 2216.885 2914.015 2217.635 ;
        RECT 5.520 2216.715 6.900 2216.885 ;
        RECT 2906.300 2216.715 2906.740 2216.885 ;
        RECT 2912.720 2216.715 2914.100 2216.885 ;
        RECT 5.605 2215.965 6.815 2216.715 ;
        RECT 2906.365 2215.990 2906.655 2216.715 ;
        RECT 2912.805 2215.965 2914.015 2216.715 ;
        RECT 5.605 2215.425 6.125 2215.965 ;
        RECT 2913.495 2215.425 2914.015 2215.965 ;
        RECT 5.605 2212.195 6.125 2212.735 ;
        RECT 2913.495 2212.195 2914.015 2212.735 ;
        RECT 5.605 2211.445 6.815 2212.195 ;
        RECT 2912.805 2211.445 2914.015 2212.195 ;
        RECT 5.520 2211.275 6.900 2211.445 ;
        RECT 2906.300 2211.275 2906.740 2211.445 ;
        RECT 2912.720 2211.275 2914.100 2211.445 ;
        RECT 5.605 2210.525 6.815 2211.275 ;
        RECT 2906.365 2210.550 2906.655 2211.275 ;
        RECT 2912.805 2210.525 2914.015 2211.275 ;
        RECT 5.605 2209.985 6.125 2210.525 ;
        RECT 2913.495 2209.985 2914.015 2210.525 ;
        RECT 5.605 2206.755 6.125 2207.295 ;
        RECT 2913.495 2206.755 2914.015 2207.295 ;
        RECT 5.605 2206.005 6.815 2206.755 ;
        RECT 2912.805 2206.005 2914.015 2206.755 ;
        RECT 5.520 2205.835 6.900 2206.005 ;
        RECT 2906.300 2205.835 2906.740 2206.005 ;
        RECT 2912.720 2205.835 2914.100 2206.005 ;
        RECT 5.605 2205.085 6.815 2205.835 ;
        RECT 2906.365 2205.110 2906.655 2205.835 ;
        RECT 2912.805 2205.085 2914.015 2205.835 ;
        RECT 5.605 2204.545 6.125 2205.085 ;
        RECT 2913.495 2204.545 2914.015 2205.085 ;
        RECT 5.605 2201.315 6.125 2201.855 ;
        RECT 2913.495 2201.315 2914.015 2201.855 ;
        RECT 5.605 2200.565 6.815 2201.315 ;
        RECT 2912.805 2200.565 2914.015 2201.315 ;
        RECT 5.520 2200.395 6.900 2200.565 ;
        RECT 2906.300 2200.395 2906.740 2200.565 ;
        RECT 2912.720 2200.395 2914.100 2200.565 ;
        RECT 5.605 2199.645 6.815 2200.395 ;
        RECT 2906.365 2199.670 2906.655 2200.395 ;
        RECT 2912.805 2199.645 2914.015 2200.395 ;
        RECT 5.605 2199.105 6.125 2199.645 ;
        RECT 2913.495 2199.105 2914.015 2199.645 ;
        RECT 5.605 2195.875 6.125 2196.415 ;
        RECT 2913.495 2195.875 2914.015 2196.415 ;
        RECT 5.605 2195.125 6.815 2195.875 ;
        RECT 2912.805 2195.125 2914.015 2195.875 ;
        RECT 5.520 2194.955 6.900 2195.125 ;
        RECT 2906.300 2194.955 2906.740 2195.125 ;
        RECT 2912.720 2194.955 2914.100 2195.125 ;
        RECT 5.605 2194.205 6.815 2194.955 ;
        RECT 2906.365 2194.230 2906.655 2194.955 ;
        RECT 2912.805 2194.205 2914.015 2194.955 ;
        RECT 5.605 2193.665 6.125 2194.205 ;
        RECT 2913.495 2193.665 2914.015 2194.205 ;
        RECT 5.605 2190.435 6.125 2190.975 ;
        RECT 2913.495 2190.435 2914.015 2190.975 ;
        RECT 5.605 2189.685 6.815 2190.435 ;
        RECT 2912.805 2189.685 2914.015 2190.435 ;
        RECT 5.520 2189.515 6.900 2189.685 ;
        RECT 2906.300 2189.515 2906.740 2189.685 ;
        RECT 2912.720 2189.515 2914.100 2189.685 ;
        RECT 5.605 2188.765 6.815 2189.515 ;
        RECT 2906.365 2188.790 2906.655 2189.515 ;
        RECT 2912.805 2188.765 2914.015 2189.515 ;
        RECT 5.605 2188.225 6.125 2188.765 ;
        RECT 2913.495 2188.225 2914.015 2188.765 ;
        RECT 5.605 2184.995 6.125 2185.535 ;
        RECT 2913.495 2184.995 2914.015 2185.535 ;
        RECT 5.605 2184.245 6.815 2184.995 ;
        RECT 2912.805 2184.245 2914.015 2184.995 ;
        RECT 5.520 2184.075 6.900 2184.245 ;
        RECT 2906.300 2184.075 2906.740 2184.245 ;
        RECT 2912.720 2184.075 2914.100 2184.245 ;
        RECT 5.605 2183.325 6.815 2184.075 ;
        RECT 2906.365 2183.350 2906.655 2184.075 ;
        RECT 2912.805 2183.325 2914.015 2184.075 ;
        RECT 5.605 2182.785 6.125 2183.325 ;
        RECT 2913.495 2182.785 2914.015 2183.325 ;
        RECT 5.605 2179.555 6.125 2180.095 ;
        RECT 2913.495 2179.555 2914.015 2180.095 ;
        RECT 5.605 2178.805 6.815 2179.555 ;
        RECT 2912.805 2178.805 2914.015 2179.555 ;
        RECT 5.520 2178.635 6.900 2178.805 ;
        RECT 2906.300 2178.635 2906.740 2178.805 ;
        RECT 2912.720 2178.635 2914.100 2178.805 ;
        RECT 5.605 2177.885 6.815 2178.635 ;
        RECT 2906.365 2177.910 2906.655 2178.635 ;
        RECT 2912.805 2177.885 2914.015 2178.635 ;
        RECT 5.605 2177.345 6.125 2177.885 ;
        RECT 2913.495 2177.345 2914.015 2177.885 ;
        RECT 5.605 2174.115 6.125 2174.655 ;
        RECT 2913.495 2174.115 2914.015 2174.655 ;
        RECT 5.605 2173.365 6.815 2174.115 ;
        RECT 2912.805 2173.365 2914.015 2174.115 ;
        RECT 5.520 2173.195 6.900 2173.365 ;
        RECT 2906.300 2173.195 2906.740 2173.365 ;
        RECT 2912.720 2173.195 2914.100 2173.365 ;
        RECT 5.605 2172.445 6.815 2173.195 ;
        RECT 2906.365 2172.470 2906.655 2173.195 ;
        RECT 2912.805 2172.445 2914.015 2173.195 ;
        RECT 5.605 2171.905 6.125 2172.445 ;
        RECT 2913.495 2171.905 2914.015 2172.445 ;
        RECT 5.605 2168.675 6.125 2169.215 ;
        RECT 2913.495 2168.675 2914.015 2169.215 ;
        RECT 5.605 2167.925 6.815 2168.675 ;
        RECT 2912.805 2167.925 2914.015 2168.675 ;
        RECT 5.520 2167.755 6.900 2167.925 ;
        RECT 2906.300 2167.755 2906.740 2167.925 ;
        RECT 2912.720 2167.755 2914.100 2167.925 ;
        RECT 5.605 2167.005 6.815 2167.755 ;
        RECT 2906.365 2167.030 2906.655 2167.755 ;
        RECT 2912.805 2167.005 2914.015 2167.755 ;
        RECT 5.605 2166.465 6.125 2167.005 ;
        RECT 2913.495 2166.465 2914.015 2167.005 ;
        RECT 5.605 2163.235 6.125 2163.775 ;
        RECT 2913.495 2163.235 2914.015 2163.775 ;
        RECT 5.605 2162.485 6.815 2163.235 ;
        RECT 2912.805 2162.485 2914.015 2163.235 ;
        RECT 5.520 2162.315 6.900 2162.485 ;
        RECT 2906.300 2162.315 2906.740 2162.485 ;
        RECT 2912.720 2162.315 2914.100 2162.485 ;
        RECT 5.605 2161.565 6.815 2162.315 ;
        RECT 2906.365 2161.590 2906.655 2162.315 ;
        RECT 2912.805 2161.565 2914.015 2162.315 ;
        RECT 5.605 2161.025 6.125 2161.565 ;
        RECT 2913.495 2161.025 2914.015 2161.565 ;
        RECT 5.605 2157.795 6.125 2158.335 ;
        RECT 2913.495 2157.795 2914.015 2158.335 ;
        RECT 5.605 2157.045 6.815 2157.795 ;
        RECT 2912.805 2157.045 2914.015 2157.795 ;
        RECT 5.520 2156.875 6.900 2157.045 ;
        RECT 2906.300 2156.875 2906.740 2157.045 ;
        RECT 2912.720 2156.875 2914.100 2157.045 ;
        RECT 5.605 2156.125 6.815 2156.875 ;
        RECT 2906.365 2156.150 2906.655 2156.875 ;
        RECT 2912.805 2156.125 2914.015 2156.875 ;
        RECT 5.605 2155.585 6.125 2156.125 ;
        RECT 2913.495 2155.585 2914.015 2156.125 ;
        RECT 5.605 2152.355 6.125 2152.895 ;
        RECT 2913.495 2152.355 2914.015 2152.895 ;
        RECT 5.605 2151.605 6.815 2152.355 ;
        RECT 2912.805 2151.605 2914.015 2152.355 ;
        RECT 5.520 2151.435 6.900 2151.605 ;
        RECT 2906.300 2151.435 2906.740 2151.605 ;
        RECT 2912.720 2151.435 2914.100 2151.605 ;
        RECT 5.605 2150.685 6.815 2151.435 ;
        RECT 2906.365 2150.710 2906.655 2151.435 ;
        RECT 2912.805 2150.685 2914.015 2151.435 ;
        RECT 5.605 2150.145 6.125 2150.685 ;
        RECT 2913.495 2150.145 2914.015 2150.685 ;
        RECT 5.605 2146.915 6.125 2147.455 ;
        RECT 2913.495 2146.915 2914.015 2147.455 ;
        RECT 5.605 2146.165 6.815 2146.915 ;
        RECT 2912.805 2146.165 2914.015 2146.915 ;
        RECT 5.520 2145.995 6.900 2146.165 ;
        RECT 2906.300 2145.995 2906.740 2146.165 ;
        RECT 2912.720 2145.995 2914.100 2146.165 ;
        RECT 5.605 2145.245 6.815 2145.995 ;
        RECT 2906.365 2145.270 2906.655 2145.995 ;
        RECT 2912.805 2145.245 2914.015 2145.995 ;
        RECT 5.605 2144.705 6.125 2145.245 ;
        RECT 2913.495 2144.705 2914.015 2145.245 ;
        RECT 5.605 2141.475 6.125 2142.015 ;
        RECT 2913.495 2141.475 2914.015 2142.015 ;
        RECT 5.605 2140.725 6.815 2141.475 ;
        RECT 2912.805 2140.725 2914.015 2141.475 ;
        RECT 5.520 2140.555 6.900 2140.725 ;
        RECT 2906.300 2140.555 2906.740 2140.725 ;
        RECT 2912.720 2140.555 2914.100 2140.725 ;
        RECT 5.605 2139.805 6.815 2140.555 ;
        RECT 2906.365 2139.830 2906.655 2140.555 ;
        RECT 2912.805 2139.805 2914.015 2140.555 ;
        RECT 5.605 2139.265 6.125 2139.805 ;
        RECT 2913.495 2139.265 2914.015 2139.805 ;
        RECT 5.605 2136.035 6.125 2136.575 ;
        RECT 2913.495 2136.035 2914.015 2136.575 ;
        RECT 5.605 2135.285 6.815 2136.035 ;
        RECT 2912.805 2135.285 2914.015 2136.035 ;
        RECT 5.520 2135.115 6.900 2135.285 ;
        RECT 2906.300 2135.115 2906.740 2135.285 ;
        RECT 2912.720 2135.115 2914.100 2135.285 ;
        RECT 5.605 2134.365 6.815 2135.115 ;
        RECT 2906.365 2134.390 2906.655 2135.115 ;
        RECT 2912.805 2134.365 2914.015 2135.115 ;
        RECT 5.605 2133.825 6.125 2134.365 ;
        RECT 2913.495 2133.825 2914.015 2134.365 ;
        RECT 5.605 2130.595 6.125 2131.135 ;
        RECT 2913.495 2130.595 2914.015 2131.135 ;
        RECT 5.605 2129.845 6.815 2130.595 ;
        RECT 2912.805 2129.845 2914.015 2130.595 ;
        RECT 5.520 2129.675 6.900 2129.845 ;
        RECT 2906.300 2129.675 2906.740 2129.845 ;
        RECT 2912.720 2129.675 2914.100 2129.845 ;
        RECT 5.605 2128.925 6.815 2129.675 ;
        RECT 2906.365 2128.950 2906.655 2129.675 ;
        RECT 2912.805 2128.925 2914.015 2129.675 ;
        RECT 5.605 2128.385 6.125 2128.925 ;
        RECT 2913.495 2128.385 2914.015 2128.925 ;
        RECT 5.605 2125.155 6.125 2125.695 ;
        RECT 2913.495 2125.155 2914.015 2125.695 ;
        RECT 5.605 2124.405 6.815 2125.155 ;
        RECT 2912.805 2124.405 2914.015 2125.155 ;
        RECT 5.520 2124.235 6.900 2124.405 ;
        RECT 2906.300 2124.235 2906.740 2124.405 ;
        RECT 2912.720 2124.235 2914.100 2124.405 ;
        RECT 5.605 2123.485 6.815 2124.235 ;
        RECT 2906.365 2123.510 2906.655 2124.235 ;
        RECT 2912.805 2123.485 2914.015 2124.235 ;
        RECT 5.605 2122.945 6.125 2123.485 ;
        RECT 2913.495 2122.945 2914.015 2123.485 ;
        RECT 5.605 2119.715 6.125 2120.255 ;
        RECT 2913.495 2119.715 2914.015 2120.255 ;
        RECT 5.605 2118.965 6.815 2119.715 ;
        RECT 2912.805 2118.965 2914.015 2119.715 ;
        RECT 5.520 2118.795 6.900 2118.965 ;
        RECT 2906.300 2118.795 2906.740 2118.965 ;
        RECT 2909.040 2118.795 2910.420 2118.965 ;
        RECT 2912.720 2118.795 2914.100 2118.965 ;
        RECT 5.605 2118.045 6.815 2118.795 ;
        RECT 2906.365 2118.070 2906.655 2118.795 ;
        RECT 2909.815 2118.135 2910.155 2118.795 ;
        RECT 2912.805 2118.045 2914.015 2118.795 ;
        RECT 5.605 2117.505 6.125 2118.045 ;
        RECT 2913.495 2117.505 2914.015 2118.045 ;
        RECT 5.605 2114.275 6.125 2114.815 ;
        RECT 2913.495 2114.275 2914.015 2114.815 ;
        RECT 5.605 2113.525 6.815 2114.275 ;
        RECT 2912.805 2113.525 2914.015 2114.275 ;
        RECT 5.520 2113.355 6.900 2113.525 ;
        RECT 2906.300 2113.355 2906.740 2113.525 ;
        RECT 2912.720 2113.355 2914.100 2113.525 ;
        RECT 5.605 2112.605 6.815 2113.355 ;
        RECT 2906.365 2112.630 2906.655 2113.355 ;
        RECT 2912.805 2112.605 2914.015 2113.355 ;
        RECT 5.605 2112.065 6.125 2112.605 ;
        RECT 2913.495 2112.065 2914.015 2112.605 ;
        RECT 5.605 2108.835 6.125 2109.375 ;
        RECT 2913.495 2108.835 2914.015 2109.375 ;
        RECT 5.605 2108.085 6.815 2108.835 ;
        RECT 2912.805 2108.085 2914.015 2108.835 ;
        RECT 5.520 2107.915 6.900 2108.085 ;
        RECT 2906.300 2107.915 2906.740 2108.085 ;
        RECT 2912.720 2107.915 2914.100 2108.085 ;
        RECT 5.605 2107.165 6.815 2107.915 ;
        RECT 2906.365 2107.190 2906.655 2107.915 ;
        RECT 2912.805 2107.165 2914.015 2107.915 ;
        RECT 5.605 2106.625 6.125 2107.165 ;
        RECT 2913.495 2106.625 2914.015 2107.165 ;
        RECT 5.605 2103.395 6.125 2103.935 ;
        RECT 2913.495 2103.395 2914.015 2103.935 ;
        RECT 5.605 2102.645 6.815 2103.395 ;
        RECT 2912.805 2102.645 2914.015 2103.395 ;
        RECT 5.520 2102.475 6.900 2102.645 ;
        RECT 2906.300 2102.475 2906.740 2102.645 ;
        RECT 2912.720 2102.475 2914.100 2102.645 ;
        RECT 5.605 2101.725 6.815 2102.475 ;
        RECT 2906.365 2101.750 2906.655 2102.475 ;
        RECT 2912.805 2101.725 2914.015 2102.475 ;
        RECT 5.605 2101.185 6.125 2101.725 ;
        RECT 2913.495 2101.185 2914.015 2101.725 ;
        RECT 5.605 2097.955 6.125 2098.495 ;
        RECT 2913.495 2097.955 2914.015 2098.495 ;
        RECT 5.605 2097.205 6.815 2097.955 ;
        RECT 2912.805 2097.205 2914.015 2097.955 ;
        RECT 5.520 2097.035 6.900 2097.205 ;
        RECT 2906.300 2097.035 2906.740 2097.205 ;
        RECT 2912.720 2097.035 2914.100 2097.205 ;
        RECT 5.605 2096.285 6.815 2097.035 ;
        RECT 2906.365 2096.310 2906.655 2097.035 ;
        RECT 2912.805 2096.285 2914.015 2097.035 ;
        RECT 5.605 2095.745 6.125 2096.285 ;
        RECT 2913.495 2095.745 2914.015 2096.285 ;
        RECT 5.605 2092.515 6.125 2093.055 ;
        RECT 2913.495 2092.515 2914.015 2093.055 ;
        RECT 5.605 2091.765 6.815 2092.515 ;
        RECT 2912.805 2091.765 2914.015 2092.515 ;
        RECT 5.520 2091.595 6.900 2091.765 ;
        RECT 2906.300 2091.595 2906.740 2091.765 ;
        RECT 2912.720 2091.595 2914.100 2091.765 ;
        RECT 5.605 2090.845 6.815 2091.595 ;
        RECT 2906.365 2090.870 2906.655 2091.595 ;
        RECT 2912.805 2090.845 2914.015 2091.595 ;
        RECT 5.605 2090.305 6.125 2090.845 ;
        RECT 2913.495 2090.305 2914.015 2090.845 ;
        RECT 5.605 2087.075 6.125 2087.615 ;
        RECT 2913.495 2087.075 2914.015 2087.615 ;
        RECT 5.605 2086.325 6.815 2087.075 ;
        RECT 2912.805 2086.325 2914.015 2087.075 ;
        RECT 5.520 2086.155 6.900 2086.325 ;
        RECT 2906.300 2086.155 2906.740 2086.325 ;
        RECT 2912.720 2086.155 2914.100 2086.325 ;
        RECT 5.605 2085.405 6.815 2086.155 ;
        RECT 2906.365 2085.430 2906.655 2086.155 ;
        RECT 2912.805 2085.405 2914.015 2086.155 ;
        RECT 5.605 2084.865 6.125 2085.405 ;
        RECT 2913.495 2084.865 2914.015 2085.405 ;
        RECT 5.605 2081.635 6.125 2082.175 ;
        RECT 2913.495 2081.635 2914.015 2082.175 ;
        RECT 5.605 2080.885 6.815 2081.635 ;
        RECT 2912.805 2080.885 2914.015 2081.635 ;
        RECT 5.520 2080.715 6.900 2080.885 ;
        RECT 2906.300 2080.715 2906.740 2080.885 ;
        RECT 2912.720 2080.715 2914.100 2080.885 ;
        RECT 5.605 2079.965 6.815 2080.715 ;
        RECT 2906.365 2079.990 2906.655 2080.715 ;
        RECT 2912.805 2079.965 2914.015 2080.715 ;
        RECT 5.605 2079.425 6.125 2079.965 ;
        RECT 2913.495 2079.425 2914.015 2079.965 ;
        RECT 5.605 2076.195 6.125 2076.735 ;
        RECT 2913.495 2076.195 2914.015 2076.735 ;
        RECT 5.605 2075.445 6.815 2076.195 ;
        RECT 2912.805 2075.445 2914.015 2076.195 ;
        RECT 5.520 2075.275 6.900 2075.445 ;
        RECT 2906.300 2075.275 2906.740 2075.445 ;
        RECT 2912.720 2075.275 2914.100 2075.445 ;
        RECT 5.605 2074.525 6.815 2075.275 ;
        RECT 2906.365 2074.550 2906.655 2075.275 ;
        RECT 2912.805 2074.525 2914.015 2075.275 ;
        RECT 5.605 2073.985 6.125 2074.525 ;
        RECT 2913.495 2073.985 2914.015 2074.525 ;
        RECT 5.605 2070.755 6.125 2071.295 ;
        RECT 2913.495 2070.755 2914.015 2071.295 ;
        RECT 5.605 2070.005 6.815 2070.755 ;
        RECT 2912.805 2070.005 2914.015 2070.755 ;
        RECT 5.520 2069.835 6.900 2070.005 ;
        RECT 2906.300 2069.835 2906.740 2070.005 ;
        RECT 2912.720 2069.835 2914.100 2070.005 ;
        RECT 5.605 2069.085 6.815 2069.835 ;
        RECT 2906.365 2069.110 2906.655 2069.835 ;
        RECT 2912.805 2069.085 2914.015 2069.835 ;
        RECT 5.605 2068.545 6.125 2069.085 ;
        RECT 2913.495 2068.545 2914.015 2069.085 ;
        RECT 5.605 2065.315 6.125 2065.855 ;
        RECT 2913.495 2065.315 2914.015 2065.855 ;
        RECT 5.605 2064.565 6.815 2065.315 ;
        RECT 2912.805 2064.565 2914.015 2065.315 ;
        RECT 5.520 2064.395 6.900 2064.565 ;
        RECT 2906.300 2064.395 2906.740 2064.565 ;
        RECT 2912.720 2064.395 2914.100 2064.565 ;
        RECT 5.605 2063.645 6.815 2064.395 ;
        RECT 2906.365 2063.670 2906.655 2064.395 ;
        RECT 2912.805 2063.645 2914.015 2064.395 ;
        RECT 5.605 2063.105 6.125 2063.645 ;
        RECT 2913.495 2063.105 2914.015 2063.645 ;
        RECT 5.605 2059.875 6.125 2060.415 ;
        RECT 2913.495 2059.875 2914.015 2060.415 ;
        RECT 5.605 2059.125 6.815 2059.875 ;
        RECT 2912.805 2059.125 2914.015 2059.875 ;
        RECT 5.520 2058.955 6.900 2059.125 ;
        RECT 2906.300 2058.955 2906.740 2059.125 ;
        RECT 2912.720 2058.955 2914.100 2059.125 ;
        RECT 5.605 2058.205 6.815 2058.955 ;
        RECT 2906.365 2058.230 2906.655 2058.955 ;
        RECT 2912.805 2058.205 2914.015 2058.955 ;
        RECT 5.605 2057.665 6.125 2058.205 ;
        RECT 2913.495 2057.665 2914.015 2058.205 ;
        RECT 5.605 2054.435 6.125 2054.975 ;
        RECT 2913.495 2054.435 2914.015 2054.975 ;
        RECT 5.605 2053.685 6.815 2054.435 ;
        RECT 2912.805 2053.685 2914.015 2054.435 ;
        RECT 5.520 2053.515 6.900 2053.685 ;
        RECT 2906.300 2053.515 2906.740 2053.685 ;
        RECT 2912.720 2053.515 2914.100 2053.685 ;
        RECT 5.605 2052.765 6.815 2053.515 ;
        RECT 2906.365 2052.790 2906.655 2053.515 ;
        RECT 2912.805 2052.765 2914.015 2053.515 ;
        RECT 5.605 2052.225 6.125 2052.765 ;
        RECT 2913.495 2052.225 2914.015 2052.765 ;
        RECT 5.605 2048.995 6.125 2049.535 ;
        RECT 2913.495 2048.995 2914.015 2049.535 ;
        RECT 5.605 2048.245 6.815 2048.995 ;
        RECT 2912.805 2048.245 2914.015 2048.995 ;
        RECT 5.520 2048.075 6.900 2048.245 ;
        RECT 2906.300 2048.075 2906.740 2048.245 ;
        RECT 2912.720 2048.075 2914.100 2048.245 ;
        RECT 5.605 2047.325 6.815 2048.075 ;
        RECT 2906.365 2047.350 2906.655 2048.075 ;
        RECT 2912.805 2047.325 2914.015 2048.075 ;
        RECT 5.605 2046.785 6.125 2047.325 ;
        RECT 2913.495 2046.785 2914.015 2047.325 ;
        RECT 5.605 2043.555 6.125 2044.095 ;
        RECT 2913.495 2043.555 2914.015 2044.095 ;
        RECT 5.605 2042.805 6.815 2043.555 ;
        RECT 2912.805 2042.805 2914.015 2043.555 ;
        RECT 5.520 2042.635 6.900 2042.805 ;
        RECT 2906.300 2042.635 2906.740 2042.805 ;
        RECT 2912.720 2042.635 2914.100 2042.805 ;
        RECT 5.605 2041.885 6.815 2042.635 ;
        RECT 2906.365 2041.910 2906.655 2042.635 ;
        RECT 2912.805 2041.885 2914.015 2042.635 ;
        RECT 5.605 2041.345 6.125 2041.885 ;
        RECT 2913.495 2041.345 2914.015 2041.885 ;
        RECT 5.605 2038.115 6.125 2038.655 ;
        RECT 2913.495 2038.115 2914.015 2038.655 ;
        RECT 5.605 2037.365 6.815 2038.115 ;
        RECT 2912.805 2037.365 2914.015 2038.115 ;
        RECT 5.520 2037.195 6.900 2037.365 ;
        RECT 2906.300 2037.195 2906.740 2037.365 ;
        RECT 2912.720 2037.195 2914.100 2037.365 ;
        RECT 5.605 2036.445 6.815 2037.195 ;
        RECT 2906.365 2036.470 2906.655 2037.195 ;
        RECT 2912.805 2036.445 2914.015 2037.195 ;
        RECT 5.605 2035.905 6.125 2036.445 ;
        RECT 2913.495 2035.905 2914.015 2036.445 ;
        RECT 5.605 2032.675 6.125 2033.215 ;
        RECT 2913.495 2032.675 2914.015 2033.215 ;
        RECT 5.605 2031.925 6.815 2032.675 ;
        RECT 2912.805 2031.925 2914.015 2032.675 ;
        RECT 5.520 2031.755 6.900 2031.925 ;
        RECT 2906.300 2031.755 2906.740 2031.925 ;
        RECT 2912.720 2031.755 2914.100 2031.925 ;
        RECT 5.605 2031.005 6.815 2031.755 ;
        RECT 2906.365 2031.030 2906.655 2031.755 ;
        RECT 2912.805 2031.005 2914.015 2031.755 ;
        RECT 5.605 2030.465 6.125 2031.005 ;
        RECT 2913.495 2030.465 2914.015 2031.005 ;
        RECT 5.605 2027.235 6.125 2027.775 ;
        RECT 2913.495 2027.235 2914.015 2027.775 ;
        RECT 5.605 2026.485 6.815 2027.235 ;
        RECT 2912.805 2026.485 2914.015 2027.235 ;
        RECT 5.520 2026.315 6.900 2026.485 ;
        RECT 2906.300 2026.315 2906.740 2026.485 ;
        RECT 2912.720 2026.315 2914.100 2026.485 ;
        RECT 5.605 2025.565 6.815 2026.315 ;
        RECT 2906.365 2025.590 2906.655 2026.315 ;
        RECT 2912.805 2025.565 2914.015 2026.315 ;
        RECT 5.605 2025.025 6.125 2025.565 ;
        RECT 2913.495 2025.025 2914.015 2025.565 ;
        RECT 5.605 2021.795 6.125 2022.335 ;
        RECT 2913.495 2021.795 2914.015 2022.335 ;
        RECT 5.605 2021.045 6.815 2021.795 ;
        RECT 2912.805 2021.045 2914.015 2021.795 ;
        RECT 5.520 2020.875 6.900 2021.045 ;
        RECT 2906.300 2020.875 2906.740 2021.045 ;
        RECT 2912.720 2020.875 2914.100 2021.045 ;
        RECT 5.605 2020.125 6.815 2020.875 ;
        RECT 2906.365 2020.150 2906.655 2020.875 ;
        RECT 2912.805 2020.125 2914.015 2020.875 ;
        RECT 5.605 2019.585 6.125 2020.125 ;
        RECT 2913.495 2019.585 2914.015 2020.125 ;
        RECT 5.605 2016.355 6.125 2016.895 ;
        RECT 2913.495 2016.355 2914.015 2016.895 ;
        RECT 5.605 2015.605 6.815 2016.355 ;
        RECT 2912.805 2015.605 2914.015 2016.355 ;
        RECT 5.520 2015.435 6.900 2015.605 ;
        RECT 2906.300 2015.435 2906.740 2015.605 ;
        RECT 2912.720 2015.435 2914.100 2015.605 ;
        RECT 5.605 2014.685 6.815 2015.435 ;
        RECT 2906.365 2014.710 2906.655 2015.435 ;
        RECT 2912.805 2014.685 2914.015 2015.435 ;
        RECT 5.605 2014.145 6.125 2014.685 ;
        RECT 2913.495 2014.145 2914.015 2014.685 ;
        RECT 5.605 2010.915 6.125 2011.455 ;
        RECT 2913.495 2010.915 2914.015 2011.455 ;
        RECT 5.605 2010.165 6.815 2010.915 ;
        RECT 2912.805 2010.165 2914.015 2010.915 ;
        RECT 5.520 2009.995 6.900 2010.165 ;
        RECT 2906.300 2009.995 2906.740 2010.165 ;
        RECT 2912.720 2009.995 2914.100 2010.165 ;
        RECT 5.605 2009.245 6.815 2009.995 ;
        RECT 2906.365 2009.270 2906.655 2009.995 ;
        RECT 2912.805 2009.245 2914.015 2009.995 ;
        RECT 5.605 2008.705 6.125 2009.245 ;
        RECT 2913.495 2008.705 2914.015 2009.245 ;
        RECT 5.605 2005.475 6.125 2006.015 ;
        RECT 2913.495 2005.475 2914.015 2006.015 ;
        RECT 5.605 2004.725 6.815 2005.475 ;
        RECT 2912.805 2004.725 2914.015 2005.475 ;
        RECT 5.520 2004.555 6.900 2004.725 ;
        RECT 2906.300 2004.555 2906.740 2004.725 ;
        RECT 2912.720 2004.555 2914.100 2004.725 ;
        RECT 5.605 2003.805 6.815 2004.555 ;
        RECT 2906.365 2003.830 2906.655 2004.555 ;
        RECT 2912.805 2003.805 2914.015 2004.555 ;
        RECT 5.605 2003.265 6.125 2003.805 ;
        RECT 2913.495 2003.265 2914.015 2003.805 ;
        RECT 5.605 2000.035 6.125 2000.575 ;
        RECT 2913.495 2000.035 2914.015 2000.575 ;
        RECT 5.605 1999.285 6.815 2000.035 ;
        RECT 2912.805 1999.285 2914.015 2000.035 ;
        RECT 5.520 1999.115 6.900 1999.285 ;
        RECT 2906.300 1999.115 2906.740 1999.285 ;
        RECT 2912.720 1999.115 2914.100 1999.285 ;
        RECT 5.605 1998.365 6.815 1999.115 ;
        RECT 2906.365 1998.390 2906.655 1999.115 ;
        RECT 2912.805 1998.365 2914.015 1999.115 ;
        RECT 5.605 1997.825 6.125 1998.365 ;
        RECT 2913.495 1997.825 2914.015 1998.365 ;
        RECT 5.605 1994.595 6.125 1995.135 ;
        RECT 2913.495 1994.595 2914.015 1995.135 ;
        RECT 5.605 1993.845 6.815 1994.595 ;
        RECT 2912.805 1993.845 2914.015 1994.595 ;
        RECT 5.520 1993.675 6.900 1993.845 ;
        RECT 2906.300 1993.675 2906.740 1993.845 ;
        RECT 2912.720 1993.675 2914.100 1993.845 ;
        RECT 5.605 1992.925 6.815 1993.675 ;
        RECT 2906.365 1992.950 2906.655 1993.675 ;
        RECT 2912.805 1992.925 2914.015 1993.675 ;
        RECT 5.605 1992.385 6.125 1992.925 ;
        RECT 2913.495 1992.385 2914.015 1992.925 ;
        RECT 5.605 1989.155 6.125 1989.695 ;
        RECT 2913.495 1989.155 2914.015 1989.695 ;
        RECT 5.605 1988.405 6.815 1989.155 ;
        RECT 2912.805 1988.405 2914.015 1989.155 ;
        RECT 5.520 1988.235 6.900 1988.405 ;
        RECT 2906.300 1988.235 2906.740 1988.405 ;
        RECT 2912.720 1988.235 2914.100 1988.405 ;
        RECT 5.605 1987.485 6.815 1988.235 ;
        RECT 2906.365 1987.510 2906.655 1988.235 ;
        RECT 2912.805 1987.485 2914.015 1988.235 ;
        RECT 5.605 1986.945 6.125 1987.485 ;
        RECT 2913.495 1986.945 2914.015 1987.485 ;
        RECT 5.605 1983.715 6.125 1984.255 ;
        RECT 2913.495 1983.715 2914.015 1984.255 ;
        RECT 5.605 1982.965 6.815 1983.715 ;
        RECT 9.515 1982.965 9.855 1983.625 ;
        RECT 2912.805 1982.965 2914.015 1983.715 ;
        RECT 5.520 1982.795 6.900 1982.965 ;
        RECT 8.740 1982.795 10.120 1982.965 ;
        RECT 2906.300 1982.795 2906.740 1982.965 ;
        RECT 2912.720 1982.795 2914.100 1982.965 ;
        RECT 5.605 1982.045 6.815 1982.795 ;
        RECT 2906.365 1982.070 2906.655 1982.795 ;
        RECT 2912.805 1982.045 2914.015 1982.795 ;
        RECT 5.605 1981.505 6.125 1982.045 ;
        RECT 2913.495 1981.505 2914.015 1982.045 ;
        RECT 5.605 1978.275 6.125 1978.815 ;
        RECT 2913.495 1978.275 2914.015 1978.815 ;
        RECT 5.605 1977.525 6.815 1978.275 ;
        RECT 2912.805 1977.525 2914.015 1978.275 ;
        RECT 5.520 1977.355 6.900 1977.525 ;
        RECT 2906.300 1977.355 2906.740 1977.525 ;
        RECT 2912.720 1977.355 2914.100 1977.525 ;
        RECT 5.605 1976.605 6.815 1977.355 ;
        RECT 2906.365 1976.630 2906.655 1977.355 ;
        RECT 2912.805 1976.605 2914.015 1977.355 ;
        RECT 5.605 1976.065 6.125 1976.605 ;
        RECT 2913.495 1976.065 2914.015 1976.605 ;
        RECT 5.605 1972.835 6.125 1973.375 ;
        RECT 2913.495 1972.835 2914.015 1973.375 ;
        RECT 5.605 1972.085 6.815 1972.835 ;
        RECT 2912.805 1972.085 2914.015 1972.835 ;
        RECT 5.520 1971.915 6.900 1972.085 ;
        RECT 2906.300 1971.915 2906.740 1972.085 ;
        RECT 2912.720 1971.915 2914.100 1972.085 ;
        RECT 5.605 1971.165 6.815 1971.915 ;
        RECT 2906.365 1971.190 2906.655 1971.915 ;
        RECT 2912.805 1971.165 2914.015 1971.915 ;
        RECT 5.605 1970.625 6.125 1971.165 ;
        RECT 2913.495 1970.625 2914.015 1971.165 ;
        RECT 5.605 1967.395 6.125 1967.935 ;
        RECT 2913.495 1967.395 2914.015 1967.935 ;
        RECT 5.605 1966.645 6.815 1967.395 ;
        RECT 2912.805 1966.645 2914.015 1967.395 ;
        RECT 5.520 1966.475 6.900 1966.645 ;
        RECT 2906.300 1966.475 2906.740 1966.645 ;
        RECT 2912.720 1966.475 2914.100 1966.645 ;
        RECT 5.605 1965.725 6.815 1966.475 ;
        RECT 2906.365 1965.750 2906.655 1966.475 ;
        RECT 2912.805 1965.725 2914.015 1966.475 ;
        RECT 5.605 1965.185 6.125 1965.725 ;
        RECT 2913.495 1965.185 2914.015 1965.725 ;
        RECT 5.605 1961.955 6.125 1962.495 ;
        RECT 2913.495 1961.955 2914.015 1962.495 ;
        RECT 5.605 1961.205 6.815 1961.955 ;
        RECT 2912.805 1961.205 2914.015 1961.955 ;
        RECT 5.520 1961.035 6.900 1961.205 ;
        RECT 2906.300 1961.035 2906.740 1961.205 ;
        RECT 2912.720 1961.035 2914.100 1961.205 ;
        RECT 5.605 1960.285 6.815 1961.035 ;
        RECT 2906.365 1960.310 2906.655 1961.035 ;
        RECT 2912.805 1960.285 2914.015 1961.035 ;
        RECT 5.605 1959.745 6.125 1960.285 ;
        RECT 2913.495 1959.745 2914.015 1960.285 ;
        RECT 5.605 1956.515 6.125 1957.055 ;
        RECT 2913.495 1956.515 2914.015 1957.055 ;
        RECT 5.605 1955.765 6.815 1956.515 ;
        RECT 2912.805 1955.765 2914.015 1956.515 ;
        RECT 5.520 1955.595 6.900 1955.765 ;
        RECT 8.740 1955.595 10.120 1955.765 ;
        RECT 2906.300 1955.595 2906.740 1955.765 ;
        RECT 2912.720 1955.595 2914.100 1955.765 ;
        RECT 5.605 1954.845 6.815 1955.595 ;
        RECT 9.515 1954.935 9.855 1955.595 ;
        RECT 2906.365 1954.870 2906.655 1955.595 ;
        RECT 2912.805 1954.845 2914.015 1955.595 ;
        RECT 5.605 1954.305 6.125 1954.845 ;
        RECT 2913.495 1954.305 2914.015 1954.845 ;
        RECT 5.605 1951.075 6.125 1951.615 ;
        RECT 2913.495 1951.075 2914.015 1951.615 ;
        RECT 5.605 1950.325 6.815 1951.075 ;
        RECT 2912.805 1950.325 2914.015 1951.075 ;
        RECT 5.520 1950.155 6.900 1950.325 ;
        RECT 2906.300 1950.155 2906.740 1950.325 ;
        RECT 2912.720 1950.155 2914.100 1950.325 ;
        RECT 5.605 1949.405 6.815 1950.155 ;
        RECT 2906.365 1949.430 2906.655 1950.155 ;
        RECT 2912.805 1949.405 2914.015 1950.155 ;
        RECT 5.605 1948.865 6.125 1949.405 ;
        RECT 2913.495 1948.865 2914.015 1949.405 ;
        RECT 5.605 1945.635 6.125 1946.175 ;
        RECT 2913.495 1945.635 2914.015 1946.175 ;
        RECT 5.605 1944.885 6.815 1945.635 ;
        RECT 2912.805 1944.885 2914.015 1945.635 ;
        RECT 5.520 1944.715 6.900 1944.885 ;
        RECT 2906.300 1944.715 2906.740 1944.885 ;
        RECT 2912.720 1944.715 2914.100 1944.885 ;
        RECT 5.605 1943.965 6.815 1944.715 ;
        RECT 2906.365 1943.990 2906.655 1944.715 ;
        RECT 2912.805 1943.965 2914.015 1944.715 ;
        RECT 5.605 1943.425 6.125 1943.965 ;
        RECT 2913.495 1943.425 2914.015 1943.965 ;
        RECT 5.605 1940.195 6.125 1940.735 ;
        RECT 2913.495 1940.195 2914.015 1940.735 ;
        RECT 5.605 1939.445 6.815 1940.195 ;
        RECT 2912.805 1939.445 2914.015 1940.195 ;
        RECT 5.520 1939.275 6.900 1939.445 ;
        RECT 2906.300 1939.275 2906.740 1939.445 ;
        RECT 2912.720 1939.275 2914.100 1939.445 ;
        RECT 5.605 1938.525 6.815 1939.275 ;
        RECT 2906.365 1938.550 2906.655 1939.275 ;
        RECT 2912.805 1938.525 2914.015 1939.275 ;
        RECT 5.605 1937.985 6.125 1938.525 ;
        RECT 2913.495 1937.985 2914.015 1938.525 ;
        RECT 5.605 1934.755 6.125 1935.295 ;
        RECT 2913.495 1934.755 2914.015 1935.295 ;
        RECT 5.605 1934.005 6.815 1934.755 ;
        RECT 2909.815 1934.005 2910.155 1934.665 ;
        RECT 2912.805 1934.005 2914.015 1934.755 ;
        RECT 5.520 1933.835 6.900 1934.005 ;
        RECT 2906.300 1933.835 2906.740 1934.005 ;
        RECT 2909.040 1933.835 2910.420 1934.005 ;
        RECT 2912.720 1933.835 2914.100 1934.005 ;
        RECT 5.605 1933.085 6.815 1933.835 ;
        RECT 2906.365 1933.110 2906.655 1933.835 ;
        RECT 2912.805 1933.085 2914.015 1933.835 ;
        RECT 5.605 1932.545 6.125 1933.085 ;
        RECT 2913.495 1932.545 2914.015 1933.085 ;
        RECT 5.605 1929.315 6.125 1929.855 ;
        RECT 2913.495 1929.315 2914.015 1929.855 ;
        RECT 5.605 1928.565 6.815 1929.315 ;
        RECT 2912.805 1928.565 2914.015 1929.315 ;
        RECT 5.520 1928.395 6.900 1928.565 ;
        RECT 2906.300 1928.395 2906.740 1928.565 ;
        RECT 2912.720 1928.395 2914.100 1928.565 ;
        RECT 5.605 1927.645 6.815 1928.395 ;
        RECT 2906.365 1927.670 2906.655 1928.395 ;
        RECT 2912.805 1927.645 2914.015 1928.395 ;
        RECT 5.605 1927.105 6.125 1927.645 ;
        RECT 2913.495 1927.105 2914.015 1927.645 ;
        RECT 5.605 1923.875 6.125 1924.415 ;
        RECT 2913.495 1923.875 2914.015 1924.415 ;
        RECT 5.605 1923.125 6.815 1923.875 ;
        RECT 2912.805 1923.125 2914.015 1923.875 ;
        RECT 5.520 1922.955 6.900 1923.125 ;
        RECT 2906.300 1922.955 2906.740 1923.125 ;
        RECT 2912.720 1922.955 2914.100 1923.125 ;
        RECT 5.605 1922.205 6.815 1922.955 ;
        RECT 2906.365 1922.230 2906.655 1922.955 ;
        RECT 2912.805 1922.205 2914.015 1922.955 ;
        RECT 5.605 1921.665 6.125 1922.205 ;
        RECT 2913.495 1921.665 2914.015 1922.205 ;
        RECT 5.605 1918.435 6.125 1918.975 ;
        RECT 2913.495 1918.435 2914.015 1918.975 ;
        RECT 5.605 1917.685 6.815 1918.435 ;
        RECT 2912.805 1917.685 2914.015 1918.435 ;
        RECT 5.520 1917.515 6.900 1917.685 ;
        RECT 2906.300 1917.515 2906.740 1917.685 ;
        RECT 2912.720 1917.515 2914.100 1917.685 ;
        RECT 5.605 1916.765 6.815 1917.515 ;
        RECT 2906.365 1916.790 2906.655 1917.515 ;
        RECT 2912.805 1916.765 2914.015 1917.515 ;
        RECT 5.605 1916.225 6.125 1916.765 ;
        RECT 2913.495 1916.225 2914.015 1916.765 ;
        RECT 5.605 1912.995 6.125 1913.535 ;
        RECT 2913.495 1912.995 2914.015 1913.535 ;
        RECT 5.605 1912.245 6.815 1912.995 ;
        RECT 2912.805 1912.245 2914.015 1912.995 ;
        RECT 5.520 1912.075 6.900 1912.245 ;
        RECT 2906.300 1912.075 2906.740 1912.245 ;
        RECT 2912.720 1912.075 2914.100 1912.245 ;
        RECT 5.605 1911.325 6.815 1912.075 ;
        RECT 2906.365 1911.350 2906.655 1912.075 ;
        RECT 2912.805 1911.325 2914.015 1912.075 ;
        RECT 5.605 1910.785 6.125 1911.325 ;
        RECT 2913.495 1910.785 2914.015 1911.325 ;
        RECT 5.605 1907.555 6.125 1908.095 ;
        RECT 2913.495 1907.555 2914.015 1908.095 ;
        RECT 5.605 1906.805 6.815 1907.555 ;
        RECT 2912.805 1906.805 2914.015 1907.555 ;
        RECT 5.520 1906.635 6.900 1906.805 ;
        RECT 2906.300 1906.635 2906.740 1906.805 ;
        RECT 2912.720 1906.635 2914.100 1906.805 ;
        RECT 5.605 1905.885 6.815 1906.635 ;
        RECT 2906.365 1905.910 2906.655 1906.635 ;
        RECT 2912.805 1905.885 2914.015 1906.635 ;
        RECT 5.605 1905.345 6.125 1905.885 ;
        RECT 2913.495 1905.345 2914.015 1905.885 ;
        RECT 5.605 1902.115 6.125 1902.655 ;
        RECT 2913.495 1902.115 2914.015 1902.655 ;
        RECT 5.605 1901.365 6.815 1902.115 ;
        RECT 2912.805 1901.365 2914.015 1902.115 ;
        RECT 5.520 1901.195 6.900 1901.365 ;
        RECT 2906.300 1901.195 2906.740 1901.365 ;
        RECT 2912.720 1901.195 2914.100 1901.365 ;
        RECT 5.605 1900.445 6.815 1901.195 ;
        RECT 2906.365 1900.470 2906.655 1901.195 ;
        RECT 2912.805 1900.445 2914.015 1901.195 ;
        RECT 5.605 1899.905 6.125 1900.445 ;
        RECT 2913.495 1899.905 2914.015 1900.445 ;
        RECT 5.605 1896.675 6.125 1897.215 ;
        RECT 2913.495 1896.675 2914.015 1897.215 ;
        RECT 5.605 1895.925 6.815 1896.675 ;
        RECT 2912.805 1895.925 2914.015 1896.675 ;
        RECT 5.520 1895.755 6.900 1895.925 ;
        RECT 2906.300 1895.755 2906.740 1895.925 ;
        RECT 2912.720 1895.755 2914.100 1895.925 ;
        RECT 5.605 1895.005 6.815 1895.755 ;
        RECT 2906.365 1895.030 2906.655 1895.755 ;
        RECT 2912.805 1895.005 2914.015 1895.755 ;
        RECT 5.605 1894.465 6.125 1895.005 ;
        RECT 2913.495 1894.465 2914.015 1895.005 ;
        RECT 5.605 1891.235 6.125 1891.775 ;
        RECT 2913.495 1891.235 2914.015 1891.775 ;
        RECT 5.605 1890.485 6.815 1891.235 ;
        RECT 2912.805 1890.485 2914.015 1891.235 ;
        RECT 5.520 1890.315 6.900 1890.485 ;
        RECT 2906.300 1890.315 2906.740 1890.485 ;
        RECT 2912.720 1890.315 2914.100 1890.485 ;
        RECT 5.605 1889.565 6.815 1890.315 ;
        RECT 2906.365 1889.590 2906.655 1890.315 ;
        RECT 2912.805 1889.565 2914.015 1890.315 ;
        RECT 5.605 1889.025 6.125 1889.565 ;
        RECT 2913.495 1889.025 2914.015 1889.565 ;
        RECT 5.605 1885.795 6.125 1886.335 ;
        RECT 2913.495 1885.795 2914.015 1886.335 ;
        RECT 5.605 1885.045 6.815 1885.795 ;
        RECT 2912.805 1885.045 2914.015 1885.795 ;
        RECT 5.520 1884.875 6.900 1885.045 ;
        RECT 2906.300 1884.875 2906.740 1885.045 ;
        RECT 2912.720 1884.875 2914.100 1885.045 ;
        RECT 5.605 1884.125 6.815 1884.875 ;
        RECT 2906.365 1884.150 2906.655 1884.875 ;
        RECT 2912.805 1884.125 2914.015 1884.875 ;
        RECT 5.605 1883.585 6.125 1884.125 ;
        RECT 2913.495 1883.585 2914.015 1884.125 ;
        RECT 5.605 1880.355 6.125 1880.895 ;
        RECT 2913.495 1880.355 2914.015 1880.895 ;
        RECT 5.605 1879.605 6.815 1880.355 ;
        RECT 2912.805 1879.605 2914.015 1880.355 ;
        RECT 5.520 1879.435 6.900 1879.605 ;
        RECT 2906.300 1879.435 2906.740 1879.605 ;
        RECT 2912.720 1879.435 2914.100 1879.605 ;
        RECT 5.605 1878.685 6.815 1879.435 ;
        RECT 2906.365 1878.710 2906.655 1879.435 ;
        RECT 2912.805 1878.685 2914.015 1879.435 ;
        RECT 5.605 1878.145 6.125 1878.685 ;
        RECT 2913.495 1878.145 2914.015 1878.685 ;
        RECT 5.605 1874.915 6.125 1875.455 ;
        RECT 2913.495 1874.915 2914.015 1875.455 ;
        RECT 5.605 1874.165 6.815 1874.915 ;
        RECT 2912.805 1874.165 2914.015 1874.915 ;
        RECT 5.520 1873.995 6.900 1874.165 ;
        RECT 2906.300 1873.995 2906.740 1874.165 ;
        RECT 2912.720 1873.995 2914.100 1874.165 ;
        RECT 5.605 1873.245 6.815 1873.995 ;
        RECT 2906.365 1873.270 2906.655 1873.995 ;
        RECT 2912.805 1873.245 2914.015 1873.995 ;
        RECT 5.605 1872.705 6.125 1873.245 ;
        RECT 2913.495 1872.705 2914.015 1873.245 ;
        RECT 5.605 1869.475 6.125 1870.015 ;
        RECT 2913.495 1869.475 2914.015 1870.015 ;
        RECT 5.605 1868.725 6.815 1869.475 ;
        RECT 2912.805 1868.725 2914.015 1869.475 ;
        RECT 5.520 1868.555 6.900 1868.725 ;
        RECT 2906.300 1868.555 2906.740 1868.725 ;
        RECT 2912.720 1868.555 2914.100 1868.725 ;
        RECT 5.605 1867.805 6.815 1868.555 ;
        RECT 2906.365 1867.830 2906.655 1868.555 ;
        RECT 2912.805 1867.805 2914.015 1868.555 ;
        RECT 5.605 1867.265 6.125 1867.805 ;
        RECT 2913.495 1867.265 2914.015 1867.805 ;
        RECT 5.605 1864.035 6.125 1864.575 ;
        RECT 2913.495 1864.035 2914.015 1864.575 ;
        RECT 5.605 1863.285 6.815 1864.035 ;
        RECT 2912.805 1863.285 2914.015 1864.035 ;
        RECT 5.520 1863.115 6.900 1863.285 ;
        RECT 2906.300 1863.115 2906.740 1863.285 ;
        RECT 2912.720 1863.115 2914.100 1863.285 ;
        RECT 5.605 1862.365 6.815 1863.115 ;
        RECT 2906.365 1862.390 2906.655 1863.115 ;
        RECT 2912.805 1862.365 2914.015 1863.115 ;
        RECT 5.605 1861.825 6.125 1862.365 ;
        RECT 2913.495 1861.825 2914.015 1862.365 ;
        RECT 5.605 1858.595 6.125 1859.135 ;
        RECT 2913.495 1858.595 2914.015 1859.135 ;
        RECT 5.605 1857.845 6.815 1858.595 ;
        RECT 2912.805 1857.845 2914.015 1858.595 ;
        RECT 5.520 1857.675 6.900 1857.845 ;
        RECT 2906.300 1857.675 2906.740 1857.845 ;
        RECT 2912.720 1857.675 2914.100 1857.845 ;
        RECT 5.605 1856.925 6.815 1857.675 ;
        RECT 2906.365 1856.950 2906.655 1857.675 ;
        RECT 2912.805 1856.925 2914.015 1857.675 ;
        RECT 5.605 1856.385 6.125 1856.925 ;
        RECT 2913.495 1856.385 2914.015 1856.925 ;
        RECT 5.605 1853.155 6.125 1853.695 ;
        RECT 2913.495 1853.155 2914.015 1853.695 ;
        RECT 5.605 1852.405 6.815 1853.155 ;
        RECT 2912.805 1852.405 2914.015 1853.155 ;
        RECT 5.520 1852.235 6.900 1852.405 ;
        RECT 2906.300 1852.235 2906.740 1852.405 ;
        RECT 2912.720 1852.235 2914.100 1852.405 ;
        RECT 5.605 1851.485 6.815 1852.235 ;
        RECT 2906.365 1851.510 2906.655 1852.235 ;
        RECT 2912.805 1851.485 2914.015 1852.235 ;
        RECT 5.605 1850.945 6.125 1851.485 ;
        RECT 2913.495 1850.945 2914.015 1851.485 ;
        RECT 5.605 1847.715 6.125 1848.255 ;
        RECT 2913.495 1847.715 2914.015 1848.255 ;
        RECT 5.605 1846.965 6.815 1847.715 ;
        RECT 2912.805 1846.965 2914.015 1847.715 ;
        RECT 5.520 1846.795 6.900 1846.965 ;
        RECT 2906.300 1846.795 2906.740 1846.965 ;
        RECT 2912.720 1846.795 2914.100 1846.965 ;
        RECT 5.605 1846.045 6.815 1846.795 ;
        RECT 2906.365 1846.070 2906.655 1846.795 ;
        RECT 2912.805 1846.045 2914.015 1846.795 ;
        RECT 5.605 1845.505 6.125 1846.045 ;
        RECT 2913.495 1845.505 2914.015 1846.045 ;
        RECT 5.605 1842.275 6.125 1842.815 ;
        RECT 2913.495 1842.275 2914.015 1842.815 ;
        RECT 5.605 1841.525 6.815 1842.275 ;
        RECT 2912.805 1841.525 2914.015 1842.275 ;
        RECT 5.520 1841.355 6.900 1841.525 ;
        RECT 2906.300 1841.355 2906.740 1841.525 ;
        RECT 2912.720 1841.355 2914.100 1841.525 ;
        RECT 5.605 1840.605 6.815 1841.355 ;
        RECT 2906.365 1840.630 2906.655 1841.355 ;
        RECT 2912.805 1840.605 2914.015 1841.355 ;
        RECT 5.605 1840.065 6.125 1840.605 ;
        RECT 2913.495 1840.065 2914.015 1840.605 ;
        RECT 5.605 1836.835 6.125 1837.375 ;
        RECT 2913.495 1836.835 2914.015 1837.375 ;
        RECT 5.605 1836.085 6.815 1836.835 ;
        RECT 2912.805 1836.085 2914.015 1836.835 ;
        RECT 5.520 1835.915 6.900 1836.085 ;
        RECT 2906.300 1835.915 2906.740 1836.085 ;
        RECT 2912.720 1835.915 2914.100 1836.085 ;
        RECT 5.605 1835.165 6.815 1835.915 ;
        RECT 2906.365 1835.190 2906.655 1835.915 ;
        RECT 2912.805 1835.165 2914.015 1835.915 ;
        RECT 5.605 1834.625 6.125 1835.165 ;
        RECT 2913.495 1834.625 2914.015 1835.165 ;
        RECT 5.605 1831.395 6.125 1831.935 ;
        RECT 2913.495 1831.395 2914.015 1831.935 ;
        RECT 5.605 1830.645 6.815 1831.395 ;
        RECT 2912.805 1830.645 2914.015 1831.395 ;
        RECT 5.520 1830.475 6.900 1830.645 ;
        RECT 2906.300 1830.475 2906.740 1830.645 ;
        RECT 2912.720 1830.475 2914.100 1830.645 ;
        RECT 5.605 1829.725 6.815 1830.475 ;
        RECT 2906.365 1829.750 2906.655 1830.475 ;
        RECT 2912.805 1829.725 2914.015 1830.475 ;
        RECT 5.605 1829.185 6.125 1829.725 ;
        RECT 2913.495 1829.185 2914.015 1829.725 ;
        RECT 5.605 1825.955 6.125 1826.495 ;
        RECT 2913.495 1825.955 2914.015 1826.495 ;
        RECT 5.605 1825.205 6.815 1825.955 ;
        RECT 2912.805 1825.205 2914.015 1825.955 ;
        RECT 5.520 1825.035 6.900 1825.205 ;
        RECT 2906.300 1825.035 2906.740 1825.205 ;
        RECT 2912.720 1825.035 2914.100 1825.205 ;
        RECT 5.605 1824.285 6.815 1825.035 ;
        RECT 2906.365 1824.310 2906.655 1825.035 ;
        RECT 2912.805 1824.285 2914.015 1825.035 ;
        RECT 5.605 1823.745 6.125 1824.285 ;
        RECT 2913.495 1823.745 2914.015 1824.285 ;
        RECT 5.605 1820.515 6.125 1821.055 ;
        RECT 2913.495 1820.515 2914.015 1821.055 ;
        RECT 5.605 1819.765 6.815 1820.515 ;
        RECT 2912.805 1819.765 2914.015 1820.515 ;
        RECT 5.520 1819.595 6.900 1819.765 ;
        RECT 2906.300 1819.595 2906.740 1819.765 ;
        RECT 2912.720 1819.595 2914.100 1819.765 ;
        RECT 5.605 1818.845 6.815 1819.595 ;
        RECT 2906.365 1818.870 2906.655 1819.595 ;
        RECT 2912.805 1818.845 2914.015 1819.595 ;
        RECT 5.605 1818.305 6.125 1818.845 ;
        RECT 2913.495 1818.305 2914.015 1818.845 ;
        RECT 5.605 1815.075 6.125 1815.615 ;
        RECT 2913.495 1815.075 2914.015 1815.615 ;
        RECT 5.605 1814.325 6.815 1815.075 ;
        RECT 2912.805 1814.325 2914.015 1815.075 ;
        RECT 5.520 1814.155 6.900 1814.325 ;
        RECT 2906.300 1814.155 2906.740 1814.325 ;
        RECT 2912.720 1814.155 2914.100 1814.325 ;
        RECT 5.605 1813.405 6.815 1814.155 ;
        RECT 2906.365 1813.430 2906.655 1814.155 ;
        RECT 2912.805 1813.405 2914.015 1814.155 ;
        RECT 5.605 1812.865 6.125 1813.405 ;
        RECT 2913.495 1812.865 2914.015 1813.405 ;
        RECT 5.605 1809.635 6.125 1810.175 ;
        RECT 2913.495 1809.635 2914.015 1810.175 ;
        RECT 5.605 1808.885 6.815 1809.635 ;
        RECT 2912.805 1808.885 2914.015 1809.635 ;
        RECT 5.520 1808.715 6.900 1808.885 ;
        RECT 2906.300 1808.715 2906.740 1808.885 ;
        RECT 2912.720 1808.715 2914.100 1808.885 ;
        RECT 5.605 1807.965 6.815 1808.715 ;
        RECT 2906.365 1807.990 2906.655 1808.715 ;
        RECT 2912.805 1807.965 2914.015 1808.715 ;
        RECT 5.605 1807.425 6.125 1807.965 ;
        RECT 2913.495 1807.425 2914.015 1807.965 ;
        RECT 5.605 1804.195 6.125 1804.735 ;
        RECT 2913.495 1804.195 2914.015 1804.735 ;
        RECT 5.605 1803.445 6.815 1804.195 ;
        RECT 2912.805 1803.445 2914.015 1804.195 ;
        RECT 5.520 1803.275 6.900 1803.445 ;
        RECT 2906.300 1803.275 2906.740 1803.445 ;
        RECT 2912.720 1803.275 2914.100 1803.445 ;
        RECT 5.605 1802.525 6.815 1803.275 ;
        RECT 2906.365 1802.550 2906.655 1803.275 ;
        RECT 2912.805 1802.525 2914.015 1803.275 ;
        RECT 5.605 1801.985 6.125 1802.525 ;
        RECT 2913.495 1801.985 2914.015 1802.525 ;
        RECT 5.605 1798.755 6.125 1799.295 ;
        RECT 2913.495 1798.755 2914.015 1799.295 ;
        RECT 5.605 1798.005 6.815 1798.755 ;
        RECT 2912.805 1798.005 2914.015 1798.755 ;
        RECT 5.520 1797.835 6.900 1798.005 ;
        RECT 2906.300 1797.835 2906.740 1798.005 ;
        RECT 2912.720 1797.835 2914.100 1798.005 ;
        RECT 5.605 1797.085 6.815 1797.835 ;
        RECT 2906.365 1797.110 2906.655 1797.835 ;
        RECT 2912.805 1797.085 2914.015 1797.835 ;
        RECT 5.605 1796.545 6.125 1797.085 ;
        RECT 2913.495 1796.545 2914.015 1797.085 ;
        RECT 5.605 1793.315 6.125 1793.855 ;
        RECT 2913.495 1793.315 2914.015 1793.855 ;
        RECT 5.605 1792.565 6.815 1793.315 ;
        RECT 2912.805 1792.565 2914.015 1793.315 ;
        RECT 5.520 1792.395 6.900 1792.565 ;
        RECT 2906.300 1792.395 2906.740 1792.565 ;
        RECT 2912.720 1792.395 2914.100 1792.565 ;
        RECT 5.605 1791.645 6.815 1792.395 ;
        RECT 2906.365 1791.670 2906.655 1792.395 ;
        RECT 2912.805 1791.645 2914.015 1792.395 ;
        RECT 5.605 1791.105 6.125 1791.645 ;
        RECT 2913.495 1791.105 2914.015 1791.645 ;
        RECT 5.605 1787.875 6.125 1788.415 ;
        RECT 2913.495 1787.875 2914.015 1788.415 ;
        RECT 5.605 1787.125 6.815 1787.875 ;
        RECT 2912.805 1787.125 2914.015 1787.875 ;
        RECT 5.520 1786.955 6.900 1787.125 ;
        RECT 2906.300 1786.955 2906.740 1787.125 ;
        RECT 2912.720 1786.955 2914.100 1787.125 ;
        RECT 5.605 1786.205 6.815 1786.955 ;
        RECT 2906.365 1786.230 2906.655 1786.955 ;
        RECT 2912.805 1786.205 2914.015 1786.955 ;
        RECT 5.605 1785.665 6.125 1786.205 ;
        RECT 2913.495 1785.665 2914.015 1786.205 ;
        RECT 5.605 1782.435 6.125 1782.975 ;
        RECT 2913.495 1782.435 2914.015 1782.975 ;
        RECT 5.605 1781.685 6.815 1782.435 ;
        RECT 2912.805 1781.685 2914.015 1782.435 ;
        RECT 5.520 1781.515 6.900 1781.685 ;
        RECT 2906.300 1781.515 2906.740 1781.685 ;
        RECT 2912.720 1781.515 2914.100 1781.685 ;
        RECT 5.605 1780.765 6.815 1781.515 ;
        RECT 2906.365 1780.790 2906.655 1781.515 ;
        RECT 2912.805 1780.765 2914.015 1781.515 ;
        RECT 5.605 1780.225 6.125 1780.765 ;
        RECT 2913.495 1780.225 2914.015 1780.765 ;
        RECT 5.605 1776.995 6.125 1777.535 ;
        RECT 2913.495 1776.995 2914.015 1777.535 ;
        RECT 5.605 1776.245 6.815 1776.995 ;
        RECT 9.515 1776.245 9.855 1776.905 ;
        RECT 2912.805 1776.245 2914.015 1776.995 ;
        RECT 5.520 1776.075 6.900 1776.245 ;
        RECT 8.740 1776.075 10.120 1776.245 ;
        RECT 2906.300 1776.075 2906.740 1776.245 ;
        RECT 2912.720 1776.075 2914.100 1776.245 ;
        RECT 5.605 1775.325 6.815 1776.075 ;
        RECT 2906.365 1775.350 2906.655 1776.075 ;
        RECT 2912.805 1775.325 2914.015 1776.075 ;
        RECT 5.605 1774.785 6.125 1775.325 ;
        RECT 2913.495 1774.785 2914.015 1775.325 ;
        RECT 5.605 1771.555 6.125 1772.095 ;
        RECT 2913.495 1771.555 2914.015 1772.095 ;
        RECT 5.605 1770.805 6.815 1771.555 ;
        RECT 2912.805 1770.805 2914.015 1771.555 ;
        RECT 5.520 1770.635 6.900 1770.805 ;
        RECT 2906.300 1770.635 2906.740 1770.805 ;
        RECT 2912.720 1770.635 2914.100 1770.805 ;
        RECT 5.605 1769.885 6.815 1770.635 ;
        RECT 2906.365 1769.910 2906.655 1770.635 ;
        RECT 2912.805 1769.885 2914.015 1770.635 ;
        RECT 5.605 1769.345 6.125 1769.885 ;
        RECT 2913.495 1769.345 2914.015 1769.885 ;
        RECT 5.605 1766.115 6.125 1766.655 ;
        RECT 2913.495 1766.115 2914.015 1766.655 ;
        RECT 5.605 1765.365 6.815 1766.115 ;
        RECT 2912.805 1765.365 2914.015 1766.115 ;
        RECT 5.520 1765.195 6.900 1765.365 ;
        RECT 2906.300 1765.195 2906.740 1765.365 ;
        RECT 2912.720 1765.195 2914.100 1765.365 ;
        RECT 5.605 1764.445 6.815 1765.195 ;
        RECT 2906.365 1764.470 2906.655 1765.195 ;
        RECT 2912.805 1764.445 2914.015 1765.195 ;
        RECT 5.605 1763.905 6.125 1764.445 ;
        RECT 2913.495 1763.905 2914.015 1764.445 ;
        RECT 5.605 1760.675 6.125 1761.215 ;
        RECT 2913.495 1760.675 2914.015 1761.215 ;
        RECT 5.605 1759.925 6.815 1760.675 ;
        RECT 2912.805 1759.925 2914.015 1760.675 ;
        RECT 5.520 1759.755 6.900 1759.925 ;
        RECT 2906.300 1759.755 2906.740 1759.925 ;
        RECT 2912.720 1759.755 2914.100 1759.925 ;
        RECT 5.605 1759.005 6.815 1759.755 ;
        RECT 2906.365 1759.030 2906.655 1759.755 ;
        RECT 2912.805 1759.005 2914.015 1759.755 ;
        RECT 5.605 1758.465 6.125 1759.005 ;
        RECT 2913.495 1758.465 2914.015 1759.005 ;
        RECT 5.605 1755.235 6.125 1755.775 ;
        RECT 2913.495 1755.235 2914.015 1755.775 ;
        RECT 5.605 1754.485 6.815 1755.235 ;
        RECT 2912.805 1754.485 2914.015 1755.235 ;
        RECT 5.520 1754.315 6.900 1754.485 ;
        RECT 2906.300 1754.315 2906.740 1754.485 ;
        RECT 2912.720 1754.315 2914.100 1754.485 ;
        RECT 5.605 1753.565 6.815 1754.315 ;
        RECT 2906.365 1753.590 2906.655 1754.315 ;
        RECT 2912.805 1753.565 2914.015 1754.315 ;
        RECT 5.605 1753.025 6.125 1753.565 ;
        RECT 2913.495 1753.025 2914.015 1753.565 ;
        RECT 5.605 1749.795 6.125 1750.335 ;
        RECT 2913.495 1749.795 2914.015 1750.335 ;
        RECT 5.605 1749.045 6.815 1749.795 ;
        RECT 2912.805 1749.045 2914.015 1749.795 ;
        RECT 5.520 1748.875 6.900 1749.045 ;
        RECT 2906.300 1748.875 2906.740 1749.045 ;
        RECT 2912.720 1748.875 2914.100 1749.045 ;
        RECT 5.605 1748.125 6.815 1748.875 ;
        RECT 2906.365 1748.150 2906.655 1748.875 ;
        RECT 2912.805 1748.125 2914.015 1748.875 ;
        RECT 5.605 1747.585 6.125 1748.125 ;
        RECT 2913.495 1747.585 2914.015 1748.125 ;
        RECT 5.605 1744.355 6.125 1744.895 ;
        RECT 2913.495 1744.355 2914.015 1744.895 ;
        RECT 5.605 1743.605 6.815 1744.355 ;
        RECT 2912.805 1743.605 2914.015 1744.355 ;
        RECT 5.520 1743.435 6.900 1743.605 ;
        RECT 2906.300 1743.435 2906.740 1743.605 ;
        RECT 2912.720 1743.435 2914.100 1743.605 ;
        RECT 5.605 1742.685 6.815 1743.435 ;
        RECT 2906.365 1742.710 2906.655 1743.435 ;
        RECT 2912.805 1742.685 2914.015 1743.435 ;
        RECT 5.605 1742.145 6.125 1742.685 ;
        RECT 2913.495 1742.145 2914.015 1742.685 ;
        RECT 5.605 1738.915 6.125 1739.455 ;
        RECT 2913.495 1738.915 2914.015 1739.455 ;
        RECT 5.605 1738.165 6.815 1738.915 ;
        RECT 2912.805 1738.165 2914.015 1738.915 ;
        RECT 5.520 1737.995 6.900 1738.165 ;
        RECT 2906.300 1737.995 2906.740 1738.165 ;
        RECT 2912.720 1737.995 2914.100 1738.165 ;
        RECT 5.605 1737.245 6.815 1737.995 ;
        RECT 2906.365 1737.270 2906.655 1737.995 ;
        RECT 2912.805 1737.245 2914.015 1737.995 ;
        RECT 5.605 1736.705 6.125 1737.245 ;
        RECT 2913.495 1736.705 2914.015 1737.245 ;
        RECT 5.605 1733.475 6.125 1734.015 ;
        RECT 2913.495 1733.475 2914.015 1734.015 ;
        RECT 5.605 1732.725 6.815 1733.475 ;
        RECT 2912.805 1732.725 2914.015 1733.475 ;
        RECT 5.520 1732.555 6.900 1732.725 ;
        RECT 2906.300 1732.555 2906.740 1732.725 ;
        RECT 2912.720 1732.555 2914.100 1732.725 ;
        RECT 5.605 1731.805 6.815 1732.555 ;
        RECT 2906.365 1731.830 2906.655 1732.555 ;
        RECT 2912.805 1731.805 2914.015 1732.555 ;
        RECT 5.605 1731.265 6.125 1731.805 ;
        RECT 2913.495 1731.265 2914.015 1731.805 ;
        RECT 5.605 1728.035 6.125 1728.575 ;
        RECT 2913.495 1728.035 2914.015 1728.575 ;
        RECT 5.605 1727.285 6.815 1728.035 ;
        RECT 2912.805 1727.285 2914.015 1728.035 ;
        RECT 5.520 1727.115 6.900 1727.285 ;
        RECT 2906.300 1727.115 2906.740 1727.285 ;
        RECT 2912.720 1727.115 2914.100 1727.285 ;
        RECT 5.605 1726.365 6.815 1727.115 ;
        RECT 2906.365 1726.390 2906.655 1727.115 ;
        RECT 2912.805 1726.365 2914.015 1727.115 ;
        RECT 5.605 1725.825 6.125 1726.365 ;
        RECT 2913.495 1725.825 2914.015 1726.365 ;
        RECT 5.605 1722.595 6.125 1723.135 ;
        RECT 2913.495 1722.595 2914.015 1723.135 ;
        RECT 5.605 1721.845 6.815 1722.595 ;
        RECT 2912.805 1721.845 2914.015 1722.595 ;
        RECT 5.520 1721.675 6.900 1721.845 ;
        RECT 2906.300 1721.675 2906.740 1721.845 ;
        RECT 2912.720 1721.675 2914.100 1721.845 ;
        RECT 5.605 1720.925 6.815 1721.675 ;
        RECT 2906.365 1720.950 2906.655 1721.675 ;
        RECT 2912.805 1720.925 2914.015 1721.675 ;
        RECT 5.605 1720.385 6.125 1720.925 ;
        RECT 2913.495 1720.385 2914.015 1720.925 ;
        RECT 5.605 1717.155 6.125 1717.695 ;
        RECT 2913.495 1717.155 2914.015 1717.695 ;
        RECT 5.605 1716.405 6.815 1717.155 ;
        RECT 2912.805 1716.405 2914.015 1717.155 ;
        RECT 5.520 1716.235 6.900 1716.405 ;
        RECT 2906.300 1716.235 2906.740 1716.405 ;
        RECT 2912.720 1716.235 2914.100 1716.405 ;
        RECT 5.605 1715.485 6.815 1716.235 ;
        RECT 2906.365 1715.510 2906.655 1716.235 ;
        RECT 2912.805 1715.485 2914.015 1716.235 ;
        RECT 5.605 1714.945 6.125 1715.485 ;
        RECT 2913.495 1714.945 2914.015 1715.485 ;
        RECT 5.605 1711.715 6.125 1712.255 ;
        RECT 2913.495 1711.715 2914.015 1712.255 ;
        RECT 5.605 1710.965 6.815 1711.715 ;
        RECT 2912.805 1710.965 2914.015 1711.715 ;
        RECT 5.520 1710.795 6.900 1710.965 ;
        RECT 2906.300 1710.795 2906.740 1710.965 ;
        RECT 2912.720 1710.795 2914.100 1710.965 ;
        RECT 5.605 1710.045 6.815 1710.795 ;
        RECT 2906.365 1710.070 2906.655 1710.795 ;
        RECT 2912.805 1710.045 2914.015 1710.795 ;
        RECT 5.605 1709.505 6.125 1710.045 ;
        RECT 2913.495 1709.505 2914.015 1710.045 ;
        RECT 5.605 1706.275 6.125 1706.815 ;
        RECT 2913.495 1706.275 2914.015 1706.815 ;
        RECT 5.605 1705.525 6.815 1706.275 ;
        RECT 9.515 1705.525 9.855 1706.185 ;
        RECT 2912.805 1705.525 2914.015 1706.275 ;
        RECT 5.520 1705.355 6.900 1705.525 ;
        RECT 8.740 1705.355 10.120 1705.525 ;
        RECT 2906.300 1705.355 2906.740 1705.525 ;
        RECT 2912.720 1705.355 2914.100 1705.525 ;
        RECT 5.605 1704.605 6.815 1705.355 ;
        RECT 2906.365 1704.630 2906.655 1705.355 ;
        RECT 2912.805 1704.605 2914.015 1705.355 ;
        RECT 5.605 1704.065 6.125 1704.605 ;
        RECT 2913.495 1704.065 2914.015 1704.605 ;
        RECT 5.605 1700.835 6.125 1701.375 ;
        RECT 2913.495 1700.835 2914.015 1701.375 ;
        RECT 5.605 1700.085 6.815 1700.835 ;
        RECT 2912.805 1700.085 2914.015 1700.835 ;
        RECT 5.520 1699.915 6.900 1700.085 ;
        RECT 2906.300 1699.915 2906.740 1700.085 ;
        RECT 2912.720 1699.915 2914.100 1700.085 ;
        RECT 5.605 1699.165 6.815 1699.915 ;
        RECT 2906.365 1699.190 2906.655 1699.915 ;
        RECT 2912.805 1699.165 2914.015 1699.915 ;
        RECT 5.605 1698.625 6.125 1699.165 ;
        RECT 2913.495 1698.625 2914.015 1699.165 ;
        RECT 5.605 1695.395 6.125 1695.935 ;
        RECT 2913.495 1695.395 2914.015 1695.935 ;
        RECT 5.605 1694.645 6.815 1695.395 ;
        RECT 2912.805 1694.645 2914.015 1695.395 ;
        RECT 5.520 1694.475 6.900 1694.645 ;
        RECT 2906.300 1694.475 2906.740 1694.645 ;
        RECT 2912.720 1694.475 2914.100 1694.645 ;
        RECT 5.605 1693.725 6.815 1694.475 ;
        RECT 2906.365 1693.750 2906.655 1694.475 ;
        RECT 2912.805 1693.725 2914.015 1694.475 ;
        RECT 5.605 1693.185 6.125 1693.725 ;
        RECT 2913.495 1693.185 2914.015 1693.725 ;
        RECT 5.605 1689.955 6.125 1690.495 ;
        RECT 2913.495 1689.955 2914.015 1690.495 ;
        RECT 5.605 1689.205 6.815 1689.955 ;
        RECT 2912.805 1689.205 2914.015 1689.955 ;
        RECT 5.520 1689.035 6.900 1689.205 ;
        RECT 2906.300 1689.035 2906.740 1689.205 ;
        RECT 2912.720 1689.035 2914.100 1689.205 ;
        RECT 5.605 1688.285 6.815 1689.035 ;
        RECT 2906.365 1688.310 2906.655 1689.035 ;
        RECT 2912.805 1688.285 2914.015 1689.035 ;
        RECT 5.605 1687.745 6.125 1688.285 ;
        RECT 2913.495 1687.745 2914.015 1688.285 ;
        RECT 5.605 1684.515 6.125 1685.055 ;
        RECT 2913.495 1684.515 2914.015 1685.055 ;
        RECT 5.605 1683.765 6.815 1684.515 ;
        RECT 2912.805 1683.765 2914.015 1684.515 ;
        RECT 5.520 1683.595 6.900 1683.765 ;
        RECT 2906.300 1683.595 2906.740 1683.765 ;
        RECT 2912.720 1683.595 2914.100 1683.765 ;
        RECT 5.605 1682.845 6.815 1683.595 ;
        RECT 2906.365 1682.870 2906.655 1683.595 ;
        RECT 2912.805 1682.845 2914.015 1683.595 ;
        RECT 5.605 1682.305 6.125 1682.845 ;
        RECT 2913.495 1682.305 2914.015 1682.845 ;
        RECT 5.605 1679.075 6.125 1679.615 ;
        RECT 2913.495 1679.075 2914.015 1679.615 ;
        RECT 5.605 1678.325 6.815 1679.075 ;
        RECT 2912.805 1678.325 2914.015 1679.075 ;
        RECT 5.520 1678.155 6.900 1678.325 ;
        RECT 2906.300 1678.155 2906.740 1678.325 ;
        RECT 2912.720 1678.155 2914.100 1678.325 ;
        RECT 5.605 1677.405 6.815 1678.155 ;
        RECT 2906.365 1677.430 2906.655 1678.155 ;
        RECT 2912.805 1677.405 2914.015 1678.155 ;
        RECT 5.605 1676.865 6.125 1677.405 ;
        RECT 2913.495 1676.865 2914.015 1677.405 ;
        RECT 5.605 1673.635 6.125 1674.175 ;
        RECT 2913.495 1673.635 2914.015 1674.175 ;
        RECT 5.605 1672.885 6.815 1673.635 ;
        RECT 2912.805 1672.885 2914.015 1673.635 ;
        RECT 5.520 1672.715 6.900 1672.885 ;
        RECT 2906.300 1672.715 2906.740 1672.885 ;
        RECT 2909.040 1672.715 2910.420 1672.885 ;
        RECT 2912.720 1672.715 2914.100 1672.885 ;
        RECT 5.605 1671.965 6.815 1672.715 ;
        RECT 2906.365 1671.990 2906.655 1672.715 ;
        RECT 2909.815 1672.055 2910.155 1672.715 ;
        RECT 2912.805 1671.965 2914.015 1672.715 ;
        RECT 5.605 1671.425 6.125 1671.965 ;
        RECT 2913.495 1671.425 2914.015 1671.965 ;
        RECT 5.605 1668.195 6.125 1668.735 ;
        RECT 2913.495 1668.195 2914.015 1668.735 ;
        RECT 5.605 1667.445 6.815 1668.195 ;
        RECT 2912.805 1667.445 2914.015 1668.195 ;
        RECT 5.520 1667.275 6.900 1667.445 ;
        RECT 2906.300 1667.275 2906.740 1667.445 ;
        RECT 2912.720 1667.275 2914.100 1667.445 ;
        RECT 5.605 1666.525 6.815 1667.275 ;
        RECT 2906.365 1666.550 2906.655 1667.275 ;
        RECT 2912.805 1666.525 2914.015 1667.275 ;
        RECT 5.605 1665.985 6.125 1666.525 ;
        RECT 2913.495 1665.985 2914.015 1666.525 ;
        RECT 5.605 1662.755 6.125 1663.295 ;
        RECT 2913.495 1662.755 2914.015 1663.295 ;
        RECT 5.605 1662.005 6.815 1662.755 ;
        RECT 2912.805 1662.005 2914.015 1662.755 ;
        RECT 5.520 1661.835 6.900 1662.005 ;
        RECT 2906.300 1661.835 2906.740 1662.005 ;
        RECT 2912.720 1661.835 2914.100 1662.005 ;
        RECT 5.605 1661.085 6.815 1661.835 ;
        RECT 2906.365 1661.110 2906.655 1661.835 ;
        RECT 2912.805 1661.085 2914.015 1661.835 ;
        RECT 5.605 1660.545 6.125 1661.085 ;
        RECT 2913.495 1660.545 2914.015 1661.085 ;
        RECT 5.605 1657.315 6.125 1657.855 ;
        RECT 2913.495 1657.315 2914.015 1657.855 ;
        RECT 5.605 1656.565 6.815 1657.315 ;
        RECT 2912.805 1656.565 2914.015 1657.315 ;
        RECT 5.520 1656.395 6.900 1656.565 ;
        RECT 2906.300 1656.395 2906.740 1656.565 ;
        RECT 2912.720 1656.395 2914.100 1656.565 ;
        RECT 5.605 1655.645 6.815 1656.395 ;
        RECT 2906.365 1655.670 2906.655 1656.395 ;
        RECT 2912.805 1655.645 2914.015 1656.395 ;
        RECT 5.605 1655.105 6.125 1655.645 ;
        RECT 2913.495 1655.105 2914.015 1655.645 ;
        RECT 5.605 1651.875 6.125 1652.415 ;
        RECT 2913.495 1651.875 2914.015 1652.415 ;
        RECT 5.605 1651.125 6.815 1651.875 ;
        RECT 2912.805 1651.125 2914.015 1651.875 ;
        RECT 5.520 1650.955 6.900 1651.125 ;
        RECT 2906.300 1650.955 2906.740 1651.125 ;
        RECT 2912.720 1650.955 2914.100 1651.125 ;
        RECT 5.605 1650.205 6.815 1650.955 ;
        RECT 2906.365 1650.230 2906.655 1650.955 ;
        RECT 2912.805 1650.205 2914.015 1650.955 ;
        RECT 5.605 1649.665 6.125 1650.205 ;
        RECT 2913.495 1649.665 2914.015 1650.205 ;
        RECT 5.605 1646.435 6.125 1646.975 ;
        RECT 2913.495 1646.435 2914.015 1646.975 ;
        RECT 5.605 1645.685 6.815 1646.435 ;
        RECT 2912.805 1645.685 2914.015 1646.435 ;
        RECT 5.520 1645.515 6.900 1645.685 ;
        RECT 2906.300 1645.515 2906.740 1645.685 ;
        RECT 2912.720 1645.515 2914.100 1645.685 ;
        RECT 5.605 1644.765 6.815 1645.515 ;
        RECT 2906.365 1644.790 2906.655 1645.515 ;
        RECT 2912.805 1644.765 2914.015 1645.515 ;
        RECT 5.605 1644.225 6.125 1644.765 ;
        RECT 2913.495 1644.225 2914.015 1644.765 ;
        RECT 5.605 1640.995 6.125 1641.535 ;
        RECT 2913.495 1640.995 2914.015 1641.535 ;
        RECT 5.605 1640.245 6.815 1640.995 ;
        RECT 2912.805 1640.245 2914.015 1640.995 ;
        RECT 5.520 1640.075 6.900 1640.245 ;
        RECT 2906.300 1640.075 2906.740 1640.245 ;
        RECT 2912.720 1640.075 2914.100 1640.245 ;
        RECT 5.605 1639.325 6.815 1640.075 ;
        RECT 2906.365 1639.350 2906.655 1640.075 ;
        RECT 2912.805 1639.325 2914.015 1640.075 ;
        RECT 5.605 1638.785 6.125 1639.325 ;
        RECT 2913.495 1638.785 2914.015 1639.325 ;
        RECT 5.605 1635.555 6.125 1636.095 ;
        RECT 2913.495 1635.555 2914.015 1636.095 ;
        RECT 5.605 1634.805 6.815 1635.555 ;
        RECT 2912.805 1634.805 2914.015 1635.555 ;
        RECT 5.520 1634.635 6.900 1634.805 ;
        RECT 2906.300 1634.635 2906.740 1634.805 ;
        RECT 2912.720 1634.635 2914.100 1634.805 ;
        RECT 5.605 1633.885 6.815 1634.635 ;
        RECT 2906.365 1633.910 2906.655 1634.635 ;
        RECT 2912.805 1633.885 2914.015 1634.635 ;
        RECT 5.605 1633.345 6.125 1633.885 ;
        RECT 2913.495 1633.345 2914.015 1633.885 ;
        RECT 5.605 1630.115 6.125 1630.655 ;
        RECT 2913.495 1630.115 2914.015 1630.655 ;
        RECT 5.605 1629.365 6.815 1630.115 ;
        RECT 2912.805 1629.365 2914.015 1630.115 ;
        RECT 5.520 1629.195 6.900 1629.365 ;
        RECT 2906.300 1629.195 2906.740 1629.365 ;
        RECT 2912.720 1629.195 2914.100 1629.365 ;
        RECT 5.605 1628.445 6.815 1629.195 ;
        RECT 2906.365 1628.470 2906.655 1629.195 ;
        RECT 2912.805 1628.445 2914.015 1629.195 ;
        RECT 5.605 1627.905 6.125 1628.445 ;
        RECT 2913.495 1627.905 2914.015 1628.445 ;
        RECT 5.605 1624.675 6.125 1625.215 ;
        RECT 2913.495 1624.675 2914.015 1625.215 ;
        RECT 5.605 1623.925 6.815 1624.675 ;
        RECT 2912.805 1623.925 2914.015 1624.675 ;
        RECT 5.520 1623.755 6.900 1623.925 ;
        RECT 2906.300 1623.755 2906.740 1623.925 ;
        RECT 2912.720 1623.755 2914.100 1623.925 ;
        RECT 5.605 1623.005 6.815 1623.755 ;
        RECT 2906.365 1623.030 2906.655 1623.755 ;
        RECT 2912.805 1623.005 2914.015 1623.755 ;
        RECT 5.605 1622.465 6.125 1623.005 ;
        RECT 2913.495 1622.465 2914.015 1623.005 ;
        RECT 5.605 1619.235 6.125 1619.775 ;
        RECT 2913.495 1619.235 2914.015 1619.775 ;
        RECT 5.605 1618.485 6.815 1619.235 ;
        RECT 2912.805 1618.485 2914.015 1619.235 ;
        RECT 5.520 1618.315 6.900 1618.485 ;
        RECT 2906.300 1618.315 2906.740 1618.485 ;
        RECT 2912.720 1618.315 2914.100 1618.485 ;
        RECT 5.605 1617.565 6.815 1618.315 ;
        RECT 2906.365 1617.590 2906.655 1618.315 ;
        RECT 2912.805 1617.565 2914.015 1618.315 ;
        RECT 5.605 1617.025 6.125 1617.565 ;
        RECT 2913.495 1617.025 2914.015 1617.565 ;
        RECT 5.605 1613.795 6.125 1614.335 ;
        RECT 2913.495 1613.795 2914.015 1614.335 ;
        RECT 5.605 1613.045 6.815 1613.795 ;
        RECT 2912.805 1613.045 2914.015 1613.795 ;
        RECT 5.520 1612.875 6.900 1613.045 ;
        RECT 2906.300 1612.875 2906.740 1613.045 ;
        RECT 2912.720 1612.875 2914.100 1613.045 ;
        RECT 5.605 1612.125 6.815 1612.875 ;
        RECT 2906.365 1612.150 2906.655 1612.875 ;
        RECT 2912.805 1612.125 2914.015 1612.875 ;
        RECT 5.605 1611.585 6.125 1612.125 ;
        RECT 2913.495 1611.585 2914.015 1612.125 ;
        RECT 5.605 1608.355 6.125 1608.895 ;
        RECT 2913.495 1608.355 2914.015 1608.895 ;
        RECT 5.605 1607.605 6.815 1608.355 ;
        RECT 2912.805 1607.605 2914.015 1608.355 ;
        RECT 5.520 1607.435 6.900 1607.605 ;
        RECT 2906.300 1607.435 2906.740 1607.605 ;
        RECT 2912.720 1607.435 2914.100 1607.605 ;
        RECT 5.605 1606.685 6.815 1607.435 ;
        RECT 2906.365 1606.710 2906.655 1607.435 ;
        RECT 2912.805 1606.685 2914.015 1607.435 ;
        RECT 5.605 1606.145 6.125 1606.685 ;
        RECT 2913.495 1606.145 2914.015 1606.685 ;
        RECT 5.605 1602.915 6.125 1603.455 ;
        RECT 2913.495 1602.915 2914.015 1603.455 ;
        RECT 5.605 1602.165 6.815 1602.915 ;
        RECT 2912.805 1602.165 2914.015 1602.915 ;
        RECT 5.520 1601.995 6.900 1602.165 ;
        RECT 2906.300 1601.995 2906.740 1602.165 ;
        RECT 2912.720 1601.995 2914.100 1602.165 ;
        RECT 5.605 1601.245 6.815 1601.995 ;
        RECT 2906.365 1601.270 2906.655 1601.995 ;
        RECT 2912.805 1601.245 2914.015 1601.995 ;
        RECT 5.605 1600.705 6.125 1601.245 ;
        RECT 2913.495 1600.705 2914.015 1601.245 ;
        RECT 5.605 1597.475 6.125 1598.015 ;
        RECT 2913.495 1597.475 2914.015 1598.015 ;
        RECT 5.605 1596.725 6.815 1597.475 ;
        RECT 2912.805 1596.725 2914.015 1597.475 ;
        RECT 5.520 1596.555 6.900 1596.725 ;
        RECT 2906.300 1596.555 2906.740 1596.725 ;
        RECT 2912.720 1596.555 2914.100 1596.725 ;
        RECT 5.605 1595.805 6.815 1596.555 ;
        RECT 2906.365 1595.830 2906.655 1596.555 ;
        RECT 2912.805 1595.805 2914.015 1596.555 ;
        RECT 5.605 1595.265 6.125 1595.805 ;
        RECT 2913.495 1595.265 2914.015 1595.805 ;
        RECT 5.605 1592.035 6.125 1592.575 ;
        RECT 2913.495 1592.035 2914.015 1592.575 ;
        RECT 5.605 1591.285 6.815 1592.035 ;
        RECT 2912.805 1591.285 2914.015 1592.035 ;
        RECT 5.520 1591.115 6.900 1591.285 ;
        RECT 2906.300 1591.115 2906.740 1591.285 ;
        RECT 2912.720 1591.115 2914.100 1591.285 ;
        RECT 5.605 1590.365 6.815 1591.115 ;
        RECT 2906.365 1590.390 2906.655 1591.115 ;
        RECT 2912.805 1590.365 2914.015 1591.115 ;
        RECT 5.605 1589.825 6.125 1590.365 ;
        RECT 2913.495 1589.825 2914.015 1590.365 ;
        RECT 5.605 1586.595 6.125 1587.135 ;
        RECT 2913.495 1586.595 2914.015 1587.135 ;
        RECT 5.605 1585.845 6.815 1586.595 ;
        RECT 2912.805 1585.845 2914.015 1586.595 ;
        RECT 5.520 1585.675 6.900 1585.845 ;
        RECT 2906.300 1585.675 2906.740 1585.845 ;
        RECT 2912.720 1585.675 2914.100 1585.845 ;
        RECT 5.605 1584.925 6.815 1585.675 ;
        RECT 2906.365 1584.950 2906.655 1585.675 ;
        RECT 2912.805 1584.925 2914.015 1585.675 ;
        RECT 5.605 1584.385 6.125 1584.925 ;
        RECT 2913.495 1584.385 2914.015 1584.925 ;
        RECT 5.605 1581.155 6.125 1581.695 ;
        RECT 2913.495 1581.155 2914.015 1581.695 ;
        RECT 5.605 1580.405 6.815 1581.155 ;
        RECT 9.515 1580.405 9.855 1581.065 ;
        RECT 2912.805 1580.405 2914.015 1581.155 ;
        RECT 5.520 1580.235 6.900 1580.405 ;
        RECT 8.740 1580.235 10.120 1580.405 ;
        RECT 2906.300 1580.235 2906.740 1580.405 ;
        RECT 2912.720 1580.235 2914.100 1580.405 ;
        RECT 5.605 1579.485 6.815 1580.235 ;
        RECT 2906.365 1579.510 2906.655 1580.235 ;
        RECT 2912.805 1579.485 2914.015 1580.235 ;
        RECT 5.605 1578.945 6.125 1579.485 ;
        RECT 2913.495 1578.945 2914.015 1579.485 ;
        RECT 5.605 1575.715 6.125 1576.255 ;
        RECT 2913.495 1575.715 2914.015 1576.255 ;
        RECT 5.605 1574.965 6.815 1575.715 ;
        RECT 2912.805 1574.965 2914.015 1575.715 ;
        RECT 5.520 1574.795 6.900 1574.965 ;
        RECT 2906.300 1574.795 2906.740 1574.965 ;
        RECT 2912.720 1574.795 2914.100 1574.965 ;
        RECT 5.605 1574.045 6.815 1574.795 ;
        RECT 2906.365 1574.070 2906.655 1574.795 ;
        RECT 2912.805 1574.045 2914.015 1574.795 ;
        RECT 5.605 1573.505 6.125 1574.045 ;
        RECT 2913.495 1573.505 2914.015 1574.045 ;
        RECT 5.605 1570.275 6.125 1570.815 ;
        RECT 2913.495 1570.275 2914.015 1570.815 ;
        RECT 5.605 1569.525 6.815 1570.275 ;
        RECT 2912.805 1569.525 2914.015 1570.275 ;
        RECT 5.520 1569.355 6.900 1569.525 ;
        RECT 2906.300 1569.355 2906.740 1569.525 ;
        RECT 2912.720 1569.355 2914.100 1569.525 ;
        RECT 5.605 1568.605 6.815 1569.355 ;
        RECT 2906.365 1568.630 2906.655 1569.355 ;
        RECT 2912.805 1568.605 2914.015 1569.355 ;
        RECT 5.605 1568.065 6.125 1568.605 ;
        RECT 2913.495 1568.065 2914.015 1568.605 ;
        RECT 5.605 1564.835 6.125 1565.375 ;
        RECT 2913.495 1564.835 2914.015 1565.375 ;
        RECT 5.605 1564.085 6.815 1564.835 ;
        RECT 2912.805 1564.085 2914.015 1564.835 ;
        RECT 5.520 1563.915 6.900 1564.085 ;
        RECT 2906.300 1563.915 2906.740 1564.085 ;
        RECT 2912.720 1563.915 2914.100 1564.085 ;
        RECT 5.605 1563.165 6.815 1563.915 ;
        RECT 2906.365 1563.190 2906.655 1563.915 ;
        RECT 2912.805 1563.165 2914.015 1563.915 ;
        RECT 5.605 1562.625 6.125 1563.165 ;
        RECT 2913.495 1562.625 2914.015 1563.165 ;
        RECT 5.605 1559.395 6.125 1559.935 ;
        RECT 2913.495 1559.395 2914.015 1559.935 ;
        RECT 5.605 1558.645 6.815 1559.395 ;
        RECT 2912.805 1558.645 2914.015 1559.395 ;
        RECT 5.520 1558.475 6.900 1558.645 ;
        RECT 2906.300 1558.475 2906.740 1558.645 ;
        RECT 2912.720 1558.475 2914.100 1558.645 ;
        RECT 5.605 1557.725 6.815 1558.475 ;
        RECT 2906.365 1557.750 2906.655 1558.475 ;
        RECT 2912.805 1557.725 2914.015 1558.475 ;
        RECT 5.605 1557.185 6.125 1557.725 ;
        RECT 2913.495 1557.185 2914.015 1557.725 ;
        RECT 5.605 1553.955 6.125 1554.495 ;
        RECT 2913.495 1553.955 2914.015 1554.495 ;
        RECT 5.605 1553.205 6.815 1553.955 ;
        RECT 2912.805 1553.205 2914.015 1553.955 ;
        RECT 5.520 1553.035 6.900 1553.205 ;
        RECT 2906.300 1553.035 2906.740 1553.205 ;
        RECT 2912.720 1553.035 2914.100 1553.205 ;
        RECT 5.605 1552.285 6.815 1553.035 ;
        RECT 2906.365 1552.310 2906.655 1553.035 ;
        RECT 2912.805 1552.285 2914.015 1553.035 ;
        RECT 5.605 1551.745 6.125 1552.285 ;
        RECT 2913.495 1551.745 2914.015 1552.285 ;
        RECT 5.605 1548.515 6.125 1549.055 ;
        RECT 2913.495 1548.515 2914.015 1549.055 ;
        RECT 5.605 1547.765 6.815 1548.515 ;
        RECT 2912.805 1547.765 2914.015 1548.515 ;
        RECT 5.520 1547.595 6.900 1547.765 ;
        RECT 2906.300 1547.595 2906.740 1547.765 ;
        RECT 2912.720 1547.595 2914.100 1547.765 ;
        RECT 5.605 1546.845 6.815 1547.595 ;
        RECT 2906.365 1546.870 2906.655 1547.595 ;
        RECT 2912.805 1546.845 2914.015 1547.595 ;
        RECT 5.605 1546.305 6.125 1546.845 ;
        RECT 2913.495 1546.305 2914.015 1546.845 ;
        RECT 5.605 1543.075 6.125 1543.615 ;
        RECT 2913.495 1543.075 2914.015 1543.615 ;
        RECT 5.605 1542.325 6.815 1543.075 ;
        RECT 2912.805 1542.325 2914.015 1543.075 ;
        RECT 5.520 1542.155 6.900 1542.325 ;
        RECT 2906.300 1542.155 2906.740 1542.325 ;
        RECT 2912.720 1542.155 2914.100 1542.325 ;
        RECT 5.605 1541.405 6.815 1542.155 ;
        RECT 2906.365 1541.430 2906.655 1542.155 ;
        RECT 2912.805 1541.405 2914.015 1542.155 ;
        RECT 5.605 1540.865 6.125 1541.405 ;
        RECT 2913.495 1540.865 2914.015 1541.405 ;
        RECT 5.605 1537.635 6.125 1538.175 ;
        RECT 2913.495 1537.635 2914.015 1538.175 ;
        RECT 5.605 1536.885 6.815 1537.635 ;
        RECT 2912.805 1536.885 2914.015 1537.635 ;
        RECT 5.520 1536.715 6.900 1536.885 ;
        RECT 2906.300 1536.715 2906.740 1536.885 ;
        RECT 2912.720 1536.715 2914.100 1536.885 ;
        RECT 5.605 1535.965 6.815 1536.715 ;
        RECT 2906.365 1535.990 2906.655 1536.715 ;
        RECT 2912.805 1535.965 2914.015 1536.715 ;
        RECT 5.605 1535.425 6.125 1535.965 ;
        RECT 2913.495 1535.425 2914.015 1535.965 ;
        RECT 5.605 1532.195 6.125 1532.735 ;
        RECT 2913.495 1532.195 2914.015 1532.735 ;
        RECT 5.605 1531.445 6.815 1532.195 ;
        RECT 2912.805 1531.445 2914.015 1532.195 ;
        RECT 5.520 1531.275 6.900 1531.445 ;
        RECT 2906.300 1531.275 2906.740 1531.445 ;
        RECT 2912.720 1531.275 2914.100 1531.445 ;
        RECT 5.605 1530.525 6.815 1531.275 ;
        RECT 2906.365 1530.550 2906.655 1531.275 ;
        RECT 2912.805 1530.525 2914.015 1531.275 ;
        RECT 5.605 1529.985 6.125 1530.525 ;
        RECT 2913.495 1529.985 2914.015 1530.525 ;
        RECT 5.605 1526.755 6.125 1527.295 ;
        RECT 2913.495 1526.755 2914.015 1527.295 ;
        RECT 5.605 1526.005 6.815 1526.755 ;
        RECT 2909.815 1526.005 2910.155 1526.665 ;
        RECT 2912.805 1526.005 2914.015 1526.755 ;
        RECT 5.520 1525.835 6.900 1526.005 ;
        RECT 2906.300 1525.835 2906.740 1526.005 ;
        RECT 2909.040 1525.835 2910.420 1526.005 ;
        RECT 2912.720 1525.835 2914.100 1526.005 ;
        RECT 5.605 1525.085 6.815 1525.835 ;
        RECT 2906.365 1525.110 2906.655 1525.835 ;
        RECT 2912.805 1525.085 2914.015 1525.835 ;
        RECT 5.605 1524.545 6.125 1525.085 ;
        RECT 2913.495 1524.545 2914.015 1525.085 ;
        RECT 5.605 1521.315 6.125 1521.855 ;
        RECT 2913.495 1521.315 2914.015 1521.855 ;
        RECT 5.605 1520.565 6.815 1521.315 ;
        RECT 2912.805 1520.565 2914.015 1521.315 ;
        RECT 5.520 1520.395 6.900 1520.565 ;
        RECT 2906.300 1520.395 2906.740 1520.565 ;
        RECT 2912.720 1520.395 2914.100 1520.565 ;
        RECT 5.605 1519.645 6.815 1520.395 ;
        RECT 2906.365 1519.670 2906.655 1520.395 ;
        RECT 2912.805 1519.645 2914.015 1520.395 ;
        RECT 5.605 1519.105 6.125 1519.645 ;
        RECT 2913.495 1519.105 2914.015 1519.645 ;
        RECT 5.605 1515.875 6.125 1516.415 ;
        RECT 2913.495 1515.875 2914.015 1516.415 ;
        RECT 5.605 1515.125 6.815 1515.875 ;
        RECT 2909.815 1515.125 2910.155 1515.785 ;
        RECT 2912.805 1515.125 2914.015 1515.875 ;
        RECT 5.520 1514.955 6.900 1515.125 ;
        RECT 2906.300 1514.955 2906.740 1515.125 ;
        RECT 2909.040 1514.955 2910.420 1515.125 ;
        RECT 2912.720 1514.955 2914.100 1515.125 ;
        RECT 5.605 1514.205 6.815 1514.955 ;
        RECT 2906.365 1514.230 2906.655 1514.955 ;
        RECT 2912.805 1514.205 2914.015 1514.955 ;
        RECT 5.605 1513.665 6.125 1514.205 ;
        RECT 2913.495 1513.665 2914.015 1514.205 ;
        RECT 5.605 1510.435 6.125 1510.975 ;
        RECT 2913.495 1510.435 2914.015 1510.975 ;
        RECT 5.605 1509.685 6.815 1510.435 ;
        RECT 2912.805 1509.685 2914.015 1510.435 ;
        RECT 5.520 1509.515 6.900 1509.685 ;
        RECT 2906.300 1509.515 2906.740 1509.685 ;
        RECT 2912.720 1509.515 2914.100 1509.685 ;
        RECT 5.605 1508.765 6.815 1509.515 ;
        RECT 2906.365 1508.790 2906.655 1509.515 ;
        RECT 2912.805 1508.765 2914.015 1509.515 ;
        RECT 5.605 1508.225 6.125 1508.765 ;
        RECT 2913.495 1508.225 2914.015 1508.765 ;
        RECT 5.605 1504.995 6.125 1505.535 ;
        RECT 2913.495 1504.995 2914.015 1505.535 ;
        RECT 5.605 1504.245 6.815 1504.995 ;
        RECT 2912.805 1504.245 2914.015 1504.995 ;
        RECT 5.520 1504.075 6.900 1504.245 ;
        RECT 2906.300 1504.075 2906.740 1504.245 ;
        RECT 2912.720 1504.075 2914.100 1504.245 ;
        RECT 5.605 1503.325 6.815 1504.075 ;
        RECT 2906.365 1503.350 2906.655 1504.075 ;
        RECT 2912.805 1503.325 2914.015 1504.075 ;
        RECT 5.605 1502.785 6.125 1503.325 ;
        RECT 2913.495 1502.785 2914.015 1503.325 ;
        RECT 5.605 1499.555 6.125 1500.095 ;
        RECT 2913.495 1499.555 2914.015 1500.095 ;
        RECT 5.605 1498.805 6.815 1499.555 ;
        RECT 2912.805 1498.805 2914.015 1499.555 ;
        RECT 5.520 1498.635 6.900 1498.805 ;
        RECT 2906.300 1498.635 2906.740 1498.805 ;
        RECT 2912.720 1498.635 2914.100 1498.805 ;
        RECT 5.605 1497.885 6.815 1498.635 ;
        RECT 2906.365 1497.910 2906.655 1498.635 ;
        RECT 2912.805 1497.885 2914.015 1498.635 ;
        RECT 5.605 1497.345 6.125 1497.885 ;
        RECT 2913.495 1497.345 2914.015 1497.885 ;
        RECT 5.605 1494.115 6.125 1494.655 ;
        RECT 2913.495 1494.115 2914.015 1494.655 ;
        RECT 5.605 1493.365 6.815 1494.115 ;
        RECT 2912.805 1493.365 2914.015 1494.115 ;
        RECT 5.520 1493.195 6.900 1493.365 ;
        RECT 2906.300 1493.195 2906.740 1493.365 ;
        RECT 2912.720 1493.195 2914.100 1493.365 ;
        RECT 5.605 1492.445 6.815 1493.195 ;
        RECT 2906.365 1492.470 2906.655 1493.195 ;
        RECT 2912.805 1492.445 2914.015 1493.195 ;
        RECT 5.605 1491.905 6.125 1492.445 ;
        RECT 2913.495 1491.905 2914.015 1492.445 ;
        RECT 5.605 1488.675 6.125 1489.215 ;
        RECT 2913.495 1488.675 2914.015 1489.215 ;
        RECT 5.605 1487.925 6.815 1488.675 ;
        RECT 2912.805 1487.925 2914.015 1488.675 ;
        RECT 5.520 1487.755 6.900 1487.925 ;
        RECT 2906.300 1487.755 2906.740 1487.925 ;
        RECT 2912.720 1487.755 2914.100 1487.925 ;
        RECT 5.605 1487.005 6.815 1487.755 ;
        RECT 2906.365 1487.030 2906.655 1487.755 ;
        RECT 2912.805 1487.005 2914.015 1487.755 ;
        RECT 5.605 1486.465 6.125 1487.005 ;
        RECT 2913.495 1486.465 2914.015 1487.005 ;
        RECT 5.605 1483.235 6.125 1483.775 ;
        RECT 2913.495 1483.235 2914.015 1483.775 ;
        RECT 5.605 1482.485 6.815 1483.235 ;
        RECT 2912.805 1482.485 2914.015 1483.235 ;
        RECT 5.520 1482.315 6.900 1482.485 ;
        RECT 2906.300 1482.315 2906.740 1482.485 ;
        RECT 2912.720 1482.315 2914.100 1482.485 ;
        RECT 5.605 1481.565 6.815 1482.315 ;
        RECT 2906.365 1481.590 2906.655 1482.315 ;
        RECT 2912.805 1481.565 2914.015 1482.315 ;
        RECT 5.605 1481.025 6.125 1481.565 ;
        RECT 2913.495 1481.025 2914.015 1481.565 ;
        RECT 5.605 1477.795 6.125 1478.335 ;
        RECT 2913.495 1477.795 2914.015 1478.335 ;
        RECT 5.605 1477.045 6.815 1477.795 ;
        RECT 2912.805 1477.045 2914.015 1477.795 ;
        RECT 5.520 1476.875 6.900 1477.045 ;
        RECT 2906.300 1476.875 2906.740 1477.045 ;
        RECT 2912.720 1476.875 2914.100 1477.045 ;
        RECT 5.605 1476.125 6.815 1476.875 ;
        RECT 2906.365 1476.150 2906.655 1476.875 ;
        RECT 2912.805 1476.125 2914.015 1476.875 ;
        RECT 5.605 1475.585 6.125 1476.125 ;
        RECT 2913.495 1475.585 2914.015 1476.125 ;
        RECT 5.605 1472.355 6.125 1472.895 ;
        RECT 2913.495 1472.355 2914.015 1472.895 ;
        RECT 5.605 1471.605 6.815 1472.355 ;
        RECT 2909.815 1471.605 2910.155 1472.265 ;
        RECT 2912.805 1471.605 2914.015 1472.355 ;
        RECT 5.520 1471.435 6.900 1471.605 ;
        RECT 2906.300 1471.435 2906.740 1471.605 ;
        RECT 2909.040 1471.435 2910.420 1471.605 ;
        RECT 2912.720 1471.435 2914.100 1471.605 ;
        RECT 5.605 1470.685 6.815 1471.435 ;
        RECT 2906.365 1470.710 2906.655 1471.435 ;
        RECT 2912.805 1470.685 2914.015 1471.435 ;
        RECT 5.605 1470.145 6.125 1470.685 ;
        RECT 2913.495 1470.145 2914.015 1470.685 ;
        RECT 5.605 1466.915 6.125 1467.455 ;
        RECT 2913.495 1466.915 2914.015 1467.455 ;
        RECT 5.605 1466.165 6.815 1466.915 ;
        RECT 2912.805 1466.165 2914.015 1466.915 ;
        RECT 5.520 1465.995 6.900 1466.165 ;
        RECT 2906.300 1465.995 2906.740 1466.165 ;
        RECT 2912.720 1465.995 2914.100 1466.165 ;
        RECT 5.605 1465.245 6.815 1465.995 ;
        RECT 2906.365 1465.270 2906.655 1465.995 ;
        RECT 2912.805 1465.245 2914.015 1465.995 ;
        RECT 5.605 1464.705 6.125 1465.245 ;
        RECT 2913.495 1464.705 2914.015 1465.245 ;
        RECT 5.605 1461.475 6.125 1462.015 ;
        RECT 2913.495 1461.475 2914.015 1462.015 ;
        RECT 5.605 1460.725 6.815 1461.475 ;
        RECT 2912.805 1460.725 2914.015 1461.475 ;
        RECT 5.520 1460.555 6.900 1460.725 ;
        RECT 2906.300 1460.555 2906.740 1460.725 ;
        RECT 2912.720 1460.555 2914.100 1460.725 ;
        RECT 5.605 1459.805 6.815 1460.555 ;
        RECT 2906.365 1459.830 2906.655 1460.555 ;
        RECT 2912.805 1459.805 2914.015 1460.555 ;
        RECT 5.605 1459.265 6.125 1459.805 ;
        RECT 2913.495 1459.265 2914.015 1459.805 ;
        RECT 5.605 1456.035 6.125 1456.575 ;
        RECT 2913.495 1456.035 2914.015 1456.575 ;
        RECT 5.605 1455.285 6.815 1456.035 ;
        RECT 2912.805 1455.285 2914.015 1456.035 ;
        RECT 5.520 1455.115 6.900 1455.285 ;
        RECT 2906.300 1455.115 2906.740 1455.285 ;
        RECT 2912.720 1455.115 2914.100 1455.285 ;
        RECT 5.605 1454.365 6.815 1455.115 ;
        RECT 2906.365 1454.390 2906.655 1455.115 ;
        RECT 2912.805 1454.365 2914.015 1455.115 ;
        RECT 5.605 1453.825 6.125 1454.365 ;
        RECT 2913.495 1453.825 2914.015 1454.365 ;
        RECT 5.605 1450.595 6.125 1451.135 ;
        RECT 2913.495 1450.595 2914.015 1451.135 ;
        RECT 5.605 1449.845 6.815 1450.595 ;
        RECT 2912.805 1449.845 2914.015 1450.595 ;
        RECT 5.520 1449.675 6.900 1449.845 ;
        RECT 2906.300 1449.675 2906.740 1449.845 ;
        RECT 2912.720 1449.675 2914.100 1449.845 ;
        RECT 5.605 1448.925 6.815 1449.675 ;
        RECT 2906.365 1448.950 2906.655 1449.675 ;
        RECT 2912.805 1448.925 2914.015 1449.675 ;
        RECT 5.605 1448.385 6.125 1448.925 ;
        RECT 2913.495 1448.385 2914.015 1448.925 ;
        RECT 5.605 1445.155 6.125 1445.695 ;
        RECT 2913.495 1445.155 2914.015 1445.695 ;
        RECT 5.605 1444.405 6.815 1445.155 ;
        RECT 2912.805 1444.405 2914.015 1445.155 ;
        RECT 5.520 1444.235 6.900 1444.405 ;
        RECT 2906.300 1444.235 2906.740 1444.405 ;
        RECT 2912.720 1444.235 2914.100 1444.405 ;
        RECT 5.605 1443.485 6.815 1444.235 ;
        RECT 2906.365 1443.510 2906.655 1444.235 ;
        RECT 2912.805 1443.485 2914.015 1444.235 ;
        RECT 5.605 1442.945 6.125 1443.485 ;
        RECT 2913.495 1442.945 2914.015 1443.485 ;
        RECT 5.605 1439.715 6.125 1440.255 ;
        RECT 2913.495 1439.715 2914.015 1440.255 ;
        RECT 5.605 1438.965 6.815 1439.715 ;
        RECT 2912.805 1438.965 2914.015 1439.715 ;
        RECT 5.520 1438.795 6.900 1438.965 ;
        RECT 2906.300 1438.795 2906.740 1438.965 ;
        RECT 2912.720 1438.795 2914.100 1438.965 ;
        RECT 5.605 1438.045 6.815 1438.795 ;
        RECT 2906.365 1438.070 2906.655 1438.795 ;
        RECT 2912.805 1438.045 2914.015 1438.795 ;
        RECT 5.605 1437.505 6.125 1438.045 ;
        RECT 2913.495 1437.505 2914.015 1438.045 ;
        RECT 5.605 1434.275 6.125 1434.815 ;
        RECT 2913.495 1434.275 2914.015 1434.815 ;
        RECT 5.605 1433.525 6.815 1434.275 ;
        RECT 2912.805 1433.525 2914.015 1434.275 ;
        RECT 5.520 1433.355 6.900 1433.525 ;
        RECT 2906.300 1433.355 2906.740 1433.525 ;
        RECT 2912.720 1433.355 2914.100 1433.525 ;
        RECT 5.605 1432.605 6.815 1433.355 ;
        RECT 2906.365 1432.630 2906.655 1433.355 ;
        RECT 2912.805 1432.605 2914.015 1433.355 ;
        RECT 5.605 1432.065 6.125 1432.605 ;
        RECT 2913.495 1432.065 2914.015 1432.605 ;
        RECT 5.605 1428.835 6.125 1429.375 ;
        RECT 2913.495 1428.835 2914.015 1429.375 ;
        RECT 5.605 1428.085 6.815 1428.835 ;
        RECT 2912.805 1428.085 2914.015 1428.835 ;
        RECT 5.520 1427.915 6.900 1428.085 ;
        RECT 2906.300 1427.915 2906.740 1428.085 ;
        RECT 2912.720 1427.915 2914.100 1428.085 ;
        RECT 5.605 1427.165 6.815 1427.915 ;
        RECT 2906.365 1427.190 2906.655 1427.915 ;
        RECT 2912.805 1427.165 2914.015 1427.915 ;
        RECT 5.605 1426.625 6.125 1427.165 ;
        RECT 2913.495 1426.625 2914.015 1427.165 ;
        RECT 5.605 1423.395 6.125 1423.935 ;
        RECT 2913.495 1423.395 2914.015 1423.935 ;
        RECT 5.605 1422.645 6.815 1423.395 ;
        RECT 2912.805 1422.645 2914.015 1423.395 ;
        RECT 5.520 1422.475 6.900 1422.645 ;
        RECT 2906.300 1422.475 2906.740 1422.645 ;
        RECT 2912.720 1422.475 2914.100 1422.645 ;
        RECT 5.605 1421.725 6.815 1422.475 ;
        RECT 2906.365 1421.750 2906.655 1422.475 ;
        RECT 2912.805 1421.725 2914.015 1422.475 ;
        RECT 5.605 1421.185 6.125 1421.725 ;
        RECT 2913.495 1421.185 2914.015 1421.725 ;
        RECT 5.605 1417.955 6.125 1418.495 ;
        RECT 2913.495 1417.955 2914.015 1418.495 ;
        RECT 5.605 1417.205 6.815 1417.955 ;
        RECT 2912.805 1417.205 2914.015 1417.955 ;
        RECT 5.520 1417.035 6.900 1417.205 ;
        RECT 2906.300 1417.035 2906.740 1417.205 ;
        RECT 2912.720 1417.035 2914.100 1417.205 ;
        RECT 5.605 1416.285 6.815 1417.035 ;
        RECT 2906.365 1416.310 2906.655 1417.035 ;
        RECT 2912.805 1416.285 2914.015 1417.035 ;
        RECT 5.605 1415.745 6.125 1416.285 ;
        RECT 2913.495 1415.745 2914.015 1416.285 ;
        RECT 5.605 1412.515 6.125 1413.055 ;
        RECT 2913.495 1412.515 2914.015 1413.055 ;
        RECT 5.605 1411.765 6.815 1412.515 ;
        RECT 2912.805 1411.765 2914.015 1412.515 ;
        RECT 5.520 1411.595 6.900 1411.765 ;
        RECT 2906.300 1411.595 2906.740 1411.765 ;
        RECT 2912.720 1411.595 2914.100 1411.765 ;
        RECT 5.605 1410.845 6.815 1411.595 ;
        RECT 2906.365 1410.870 2906.655 1411.595 ;
        RECT 2912.805 1410.845 2914.015 1411.595 ;
        RECT 5.605 1410.305 6.125 1410.845 ;
        RECT 2913.495 1410.305 2914.015 1410.845 ;
        RECT 5.605 1407.075 6.125 1407.615 ;
        RECT 2913.495 1407.075 2914.015 1407.615 ;
        RECT 5.605 1406.325 6.815 1407.075 ;
        RECT 2912.805 1406.325 2914.015 1407.075 ;
        RECT 5.520 1406.155 6.900 1406.325 ;
        RECT 2906.300 1406.155 2906.740 1406.325 ;
        RECT 2912.720 1406.155 2914.100 1406.325 ;
        RECT 5.605 1405.405 6.815 1406.155 ;
        RECT 2906.365 1405.430 2906.655 1406.155 ;
        RECT 2912.805 1405.405 2914.015 1406.155 ;
        RECT 5.605 1404.865 6.125 1405.405 ;
        RECT 2913.495 1404.865 2914.015 1405.405 ;
        RECT 5.605 1401.635 6.125 1402.175 ;
        RECT 2913.495 1401.635 2914.015 1402.175 ;
        RECT 5.605 1400.885 6.815 1401.635 ;
        RECT 2912.805 1400.885 2914.015 1401.635 ;
        RECT 5.520 1400.715 6.900 1400.885 ;
        RECT 2906.300 1400.715 2906.740 1400.885 ;
        RECT 2912.720 1400.715 2914.100 1400.885 ;
        RECT 5.605 1399.965 6.815 1400.715 ;
        RECT 2906.365 1399.990 2906.655 1400.715 ;
        RECT 2912.805 1399.965 2914.015 1400.715 ;
        RECT 5.605 1399.425 6.125 1399.965 ;
        RECT 2913.495 1399.425 2914.015 1399.965 ;
        RECT 5.605 1396.195 6.125 1396.735 ;
        RECT 2913.495 1396.195 2914.015 1396.735 ;
        RECT 5.605 1395.445 6.815 1396.195 ;
        RECT 2912.805 1395.445 2914.015 1396.195 ;
        RECT 5.520 1395.275 6.900 1395.445 ;
        RECT 2906.300 1395.275 2906.740 1395.445 ;
        RECT 2912.720 1395.275 2914.100 1395.445 ;
        RECT 5.605 1394.525 6.815 1395.275 ;
        RECT 2906.365 1394.550 2906.655 1395.275 ;
        RECT 2912.805 1394.525 2914.015 1395.275 ;
        RECT 5.605 1393.985 6.125 1394.525 ;
        RECT 2913.495 1393.985 2914.015 1394.525 ;
        RECT 5.605 1390.755 6.125 1391.295 ;
        RECT 2913.495 1390.755 2914.015 1391.295 ;
        RECT 5.605 1390.005 6.815 1390.755 ;
        RECT 2912.805 1390.005 2914.015 1390.755 ;
        RECT 5.520 1389.835 6.900 1390.005 ;
        RECT 2906.300 1389.835 2906.740 1390.005 ;
        RECT 2912.720 1389.835 2914.100 1390.005 ;
        RECT 5.605 1389.085 6.815 1389.835 ;
        RECT 2906.365 1389.110 2906.655 1389.835 ;
        RECT 2912.805 1389.085 2914.015 1389.835 ;
        RECT 5.605 1388.545 6.125 1389.085 ;
        RECT 2913.495 1388.545 2914.015 1389.085 ;
        RECT 5.605 1385.315 6.125 1385.855 ;
        RECT 2913.495 1385.315 2914.015 1385.855 ;
        RECT 5.605 1384.565 6.815 1385.315 ;
        RECT 2912.805 1384.565 2914.015 1385.315 ;
        RECT 5.520 1384.395 6.900 1384.565 ;
        RECT 2906.300 1384.395 2906.740 1384.565 ;
        RECT 2912.720 1384.395 2914.100 1384.565 ;
        RECT 5.605 1383.645 6.815 1384.395 ;
        RECT 2906.365 1383.670 2906.655 1384.395 ;
        RECT 2912.805 1383.645 2914.015 1384.395 ;
        RECT 5.605 1383.105 6.125 1383.645 ;
        RECT 2913.495 1383.105 2914.015 1383.645 ;
        RECT 5.605 1379.875 6.125 1380.415 ;
        RECT 2913.495 1379.875 2914.015 1380.415 ;
        RECT 5.605 1379.125 6.815 1379.875 ;
        RECT 2912.805 1379.125 2914.015 1379.875 ;
        RECT 5.520 1378.955 6.900 1379.125 ;
        RECT 2906.300 1378.955 2906.740 1379.125 ;
        RECT 2912.720 1378.955 2914.100 1379.125 ;
        RECT 5.605 1378.205 6.815 1378.955 ;
        RECT 2906.365 1378.230 2906.655 1378.955 ;
        RECT 2912.805 1378.205 2914.015 1378.955 ;
        RECT 5.605 1377.665 6.125 1378.205 ;
        RECT 2913.495 1377.665 2914.015 1378.205 ;
        RECT 5.605 1374.435 6.125 1374.975 ;
        RECT 2913.495 1374.435 2914.015 1374.975 ;
        RECT 5.605 1373.685 6.815 1374.435 ;
        RECT 2912.805 1373.685 2914.015 1374.435 ;
        RECT 5.520 1373.515 6.900 1373.685 ;
        RECT 2906.300 1373.515 2906.740 1373.685 ;
        RECT 2912.720 1373.515 2914.100 1373.685 ;
        RECT 5.605 1372.765 6.815 1373.515 ;
        RECT 2906.365 1372.790 2906.655 1373.515 ;
        RECT 2912.805 1372.765 2914.015 1373.515 ;
        RECT 5.605 1372.225 6.125 1372.765 ;
        RECT 2913.495 1372.225 2914.015 1372.765 ;
        RECT 5.605 1368.995 6.125 1369.535 ;
        RECT 2913.495 1368.995 2914.015 1369.535 ;
        RECT 5.605 1368.245 6.815 1368.995 ;
        RECT 2912.805 1368.245 2914.015 1368.995 ;
        RECT 5.520 1368.075 6.900 1368.245 ;
        RECT 2906.300 1368.075 2906.740 1368.245 ;
        RECT 2912.720 1368.075 2914.100 1368.245 ;
        RECT 5.605 1367.325 6.815 1368.075 ;
        RECT 2906.365 1367.350 2906.655 1368.075 ;
        RECT 2912.805 1367.325 2914.015 1368.075 ;
        RECT 5.605 1366.785 6.125 1367.325 ;
        RECT 2913.495 1366.785 2914.015 1367.325 ;
        RECT 5.605 1363.555 6.125 1364.095 ;
        RECT 2913.495 1363.555 2914.015 1364.095 ;
        RECT 5.605 1362.805 6.815 1363.555 ;
        RECT 2912.805 1362.805 2914.015 1363.555 ;
        RECT 5.520 1362.635 6.900 1362.805 ;
        RECT 2906.300 1362.635 2906.740 1362.805 ;
        RECT 2912.720 1362.635 2914.100 1362.805 ;
        RECT 5.605 1361.885 6.815 1362.635 ;
        RECT 2906.365 1361.910 2906.655 1362.635 ;
        RECT 2912.805 1361.885 2914.015 1362.635 ;
        RECT 5.605 1361.345 6.125 1361.885 ;
        RECT 2913.495 1361.345 2914.015 1361.885 ;
        RECT 5.605 1358.115 6.125 1358.655 ;
        RECT 2913.495 1358.115 2914.015 1358.655 ;
        RECT 5.605 1357.365 6.815 1358.115 ;
        RECT 2912.805 1357.365 2914.015 1358.115 ;
        RECT 5.520 1357.195 6.900 1357.365 ;
        RECT 2906.300 1357.195 2906.740 1357.365 ;
        RECT 2912.720 1357.195 2914.100 1357.365 ;
        RECT 5.605 1356.445 6.815 1357.195 ;
        RECT 2906.365 1356.470 2906.655 1357.195 ;
        RECT 2912.805 1356.445 2914.015 1357.195 ;
        RECT 5.605 1355.905 6.125 1356.445 ;
        RECT 2913.495 1355.905 2914.015 1356.445 ;
        RECT 5.605 1352.675 6.125 1353.215 ;
        RECT 2913.495 1352.675 2914.015 1353.215 ;
        RECT 5.605 1351.925 6.815 1352.675 ;
        RECT 2912.805 1351.925 2914.015 1352.675 ;
        RECT 5.520 1351.755 6.900 1351.925 ;
        RECT 2906.300 1351.755 2906.740 1351.925 ;
        RECT 2912.720 1351.755 2914.100 1351.925 ;
        RECT 5.605 1351.005 6.815 1351.755 ;
        RECT 2906.365 1351.030 2906.655 1351.755 ;
        RECT 2912.805 1351.005 2914.015 1351.755 ;
        RECT 5.605 1350.465 6.125 1351.005 ;
        RECT 2913.495 1350.465 2914.015 1351.005 ;
        RECT 5.605 1347.235 6.125 1347.775 ;
        RECT 2913.495 1347.235 2914.015 1347.775 ;
        RECT 5.605 1346.485 6.815 1347.235 ;
        RECT 2912.805 1346.485 2914.015 1347.235 ;
        RECT 5.520 1346.315 6.900 1346.485 ;
        RECT 2906.300 1346.315 2906.740 1346.485 ;
        RECT 2912.720 1346.315 2914.100 1346.485 ;
        RECT 5.605 1345.565 6.815 1346.315 ;
        RECT 2906.365 1345.590 2906.655 1346.315 ;
        RECT 2912.805 1345.565 2914.015 1346.315 ;
        RECT 5.605 1345.025 6.125 1345.565 ;
        RECT 2913.495 1345.025 2914.015 1345.565 ;
        RECT 5.605 1341.795 6.125 1342.335 ;
        RECT 2913.495 1341.795 2914.015 1342.335 ;
        RECT 5.605 1341.045 6.815 1341.795 ;
        RECT 2912.805 1341.045 2914.015 1341.795 ;
        RECT 5.520 1340.875 6.900 1341.045 ;
        RECT 2906.300 1340.875 2906.740 1341.045 ;
        RECT 2912.720 1340.875 2914.100 1341.045 ;
        RECT 5.605 1340.125 6.815 1340.875 ;
        RECT 2906.365 1340.150 2906.655 1340.875 ;
        RECT 2912.805 1340.125 2914.015 1340.875 ;
        RECT 5.605 1339.585 6.125 1340.125 ;
        RECT 2913.495 1339.585 2914.015 1340.125 ;
        RECT 5.605 1336.355 6.125 1336.895 ;
        RECT 2913.495 1336.355 2914.015 1336.895 ;
        RECT 5.605 1335.605 6.815 1336.355 ;
        RECT 2912.805 1335.605 2914.015 1336.355 ;
        RECT 5.520 1335.435 6.900 1335.605 ;
        RECT 2906.300 1335.435 2906.740 1335.605 ;
        RECT 2912.720 1335.435 2914.100 1335.605 ;
        RECT 5.605 1334.685 6.815 1335.435 ;
        RECT 2906.365 1334.710 2906.655 1335.435 ;
        RECT 2912.805 1334.685 2914.015 1335.435 ;
        RECT 5.605 1334.145 6.125 1334.685 ;
        RECT 2913.495 1334.145 2914.015 1334.685 ;
        RECT 5.605 1330.915 6.125 1331.455 ;
        RECT 2913.495 1330.915 2914.015 1331.455 ;
        RECT 5.605 1330.165 6.815 1330.915 ;
        RECT 2912.805 1330.165 2914.015 1330.915 ;
        RECT 5.520 1329.995 6.900 1330.165 ;
        RECT 8.740 1329.995 10.120 1330.165 ;
        RECT 2906.300 1329.995 2906.740 1330.165 ;
        RECT 2912.720 1329.995 2914.100 1330.165 ;
        RECT 5.605 1329.245 6.815 1329.995 ;
        RECT 9.515 1329.335 9.855 1329.995 ;
        RECT 2906.365 1329.270 2906.655 1329.995 ;
        RECT 2912.805 1329.245 2914.015 1329.995 ;
        RECT 5.605 1328.705 6.125 1329.245 ;
        RECT 2913.495 1328.705 2914.015 1329.245 ;
        RECT 5.605 1325.475 6.125 1326.015 ;
        RECT 2913.495 1325.475 2914.015 1326.015 ;
        RECT 5.605 1324.725 6.815 1325.475 ;
        RECT 2912.805 1324.725 2914.015 1325.475 ;
        RECT 5.520 1324.555 6.900 1324.725 ;
        RECT 2906.300 1324.555 2906.740 1324.725 ;
        RECT 2912.720 1324.555 2914.100 1324.725 ;
        RECT 5.605 1323.805 6.815 1324.555 ;
        RECT 2906.365 1323.830 2906.655 1324.555 ;
        RECT 2912.805 1323.805 2914.015 1324.555 ;
        RECT 5.605 1323.265 6.125 1323.805 ;
        RECT 2913.495 1323.265 2914.015 1323.805 ;
        RECT 5.605 1320.035 6.125 1320.575 ;
        RECT 2913.495 1320.035 2914.015 1320.575 ;
        RECT 5.605 1319.285 6.815 1320.035 ;
        RECT 2912.805 1319.285 2914.015 1320.035 ;
        RECT 5.520 1319.115 6.900 1319.285 ;
        RECT 2906.300 1319.115 2906.740 1319.285 ;
        RECT 2912.720 1319.115 2914.100 1319.285 ;
        RECT 5.605 1318.365 6.815 1319.115 ;
        RECT 2906.365 1318.390 2906.655 1319.115 ;
        RECT 2912.805 1318.365 2914.015 1319.115 ;
        RECT 5.605 1317.825 6.125 1318.365 ;
        RECT 2913.495 1317.825 2914.015 1318.365 ;
        RECT 5.605 1314.595 6.125 1315.135 ;
        RECT 2913.495 1314.595 2914.015 1315.135 ;
        RECT 5.605 1313.845 6.815 1314.595 ;
        RECT 2912.805 1313.845 2914.015 1314.595 ;
        RECT 5.520 1313.675 6.900 1313.845 ;
        RECT 2906.300 1313.675 2906.740 1313.845 ;
        RECT 2912.720 1313.675 2914.100 1313.845 ;
        RECT 5.605 1312.925 6.815 1313.675 ;
        RECT 2906.365 1312.950 2906.655 1313.675 ;
        RECT 2912.805 1312.925 2914.015 1313.675 ;
        RECT 5.605 1312.385 6.125 1312.925 ;
        RECT 2913.495 1312.385 2914.015 1312.925 ;
        RECT 5.605 1309.155 6.125 1309.695 ;
        RECT 2913.495 1309.155 2914.015 1309.695 ;
        RECT 5.605 1308.405 6.815 1309.155 ;
        RECT 2912.805 1308.405 2914.015 1309.155 ;
        RECT 5.520 1308.235 6.900 1308.405 ;
        RECT 2906.300 1308.235 2906.740 1308.405 ;
        RECT 2912.720 1308.235 2914.100 1308.405 ;
        RECT 5.605 1307.485 6.815 1308.235 ;
        RECT 2906.365 1307.510 2906.655 1308.235 ;
        RECT 2912.805 1307.485 2914.015 1308.235 ;
        RECT 5.605 1306.945 6.125 1307.485 ;
        RECT 2913.495 1306.945 2914.015 1307.485 ;
        RECT 5.605 1303.715 6.125 1304.255 ;
        RECT 2913.495 1303.715 2914.015 1304.255 ;
        RECT 5.605 1302.965 6.815 1303.715 ;
        RECT 2912.805 1302.965 2914.015 1303.715 ;
        RECT 5.520 1302.795 6.900 1302.965 ;
        RECT 2906.300 1302.795 2906.740 1302.965 ;
        RECT 2909.040 1302.795 2910.420 1302.965 ;
        RECT 2912.720 1302.795 2914.100 1302.965 ;
        RECT 5.605 1302.045 6.815 1302.795 ;
        RECT 2906.365 1302.070 2906.655 1302.795 ;
        RECT 2909.815 1302.135 2910.155 1302.795 ;
        RECT 2912.805 1302.045 2914.015 1302.795 ;
        RECT 5.605 1301.505 6.125 1302.045 ;
        RECT 2913.495 1301.505 2914.015 1302.045 ;
        RECT 5.605 1298.275 6.125 1298.815 ;
        RECT 2913.495 1298.275 2914.015 1298.815 ;
        RECT 5.605 1297.525 6.815 1298.275 ;
        RECT 2912.805 1297.525 2914.015 1298.275 ;
        RECT 5.520 1297.355 6.900 1297.525 ;
        RECT 2906.300 1297.355 2906.740 1297.525 ;
        RECT 2912.720 1297.355 2914.100 1297.525 ;
        RECT 5.605 1296.605 6.815 1297.355 ;
        RECT 2906.365 1296.630 2906.655 1297.355 ;
        RECT 2912.805 1296.605 2914.015 1297.355 ;
        RECT 5.605 1296.065 6.125 1296.605 ;
        RECT 2913.495 1296.065 2914.015 1296.605 ;
        RECT 5.605 1292.835 6.125 1293.375 ;
        RECT 2913.495 1292.835 2914.015 1293.375 ;
        RECT 5.605 1292.085 6.815 1292.835 ;
        RECT 2912.805 1292.085 2914.015 1292.835 ;
        RECT 5.520 1291.915 6.900 1292.085 ;
        RECT 2906.300 1291.915 2906.740 1292.085 ;
        RECT 2912.720 1291.915 2914.100 1292.085 ;
        RECT 5.605 1291.165 6.815 1291.915 ;
        RECT 2906.365 1291.190 2906.655 1291.915 ;
        RECT 2912.805 1291.165 2914.015 1291.915 ;
        RECT 5.605 1290.625 6.125 1291.165 ;
        RECT 2913.495 1290.625 2914.015 1291.165 ;
        RECT 5.605 1287.395 6.125 1287.935 ;
        RECT 2913.495 1287.395 2914.015 1287.935 ;
        RECT 5.605 1286.645 6.815 1287.395 ;
        RECT 2912.805 1286.645 2914.015 1287.395 ;
        RECT 5.520 1286.475 6.900 1286.645 ;
        RECT 8.740 1286.475 10.120 1286.645 ;
        RECT 2906.300 1286.475 2906.740 1286.645 ;
        RECT 2912.720 1286.475 2914.100 1286.645 ;
        RECT 5.605 1285.725 6.815 1286.475 ;
        RECT 9.515 1285.815 9.855 1286.475 ;
        RECT 2906.365 1285.750 2906.655 1286.475 ;
        RECT 2912.805 1285.725 2914.015 1286.475 ;
        RECT 5.605 1285.185 6.125 1285.725 ;
        RECT 2913.495 1285.185 2914.015 1285.725 ;
        RECT 5.605 1281.955 6.125 1282.495 ;
        RECT 2913.495 1281.955 2914.015 1282.495 ;
        RECT 5.605 1281.205 6.815 1281.955 ;
        RECT 2912.805 1281.205 2914.015 1281.955 ;
        RECT 5.520 1281.035 6.900 1281.205 ;
        RECT 2906.300 1281.035 2906.740 1281.205 ;
        RECT 2912.720 1281.035 2914.100 1281.205 ;
        RECT 5.605 1280.285 6.815 1281.035 ;
        RECT 2906.365 1280.310 2906.655 1281.035 ;
        RECT 2912.805 1280.285 2914.015 1281.035 ;
        RECT 5.605 1279.745 6.125 1280.285 ;
        RECT 2913.495 1279.745 2914.015 1280.285 ;
        RECT 5.605 1276.515 6.125 1277.055 ;
        RECT 2913.495 1276.515 2914.015 1277.055 ;
        RECT 5.605 1275.765 6.815 1276.515 ;
        RECT 2912.805 1275.765 2914.015 1276.515 ;
        RECT 5.520 1275.595 6.900 1275.765 ;
        RECT 8.740 1275.595 10.120 1275.765 ;
        RECT 2906.300 1275.595 2906.740 1275.765 ;
        RECT 2912.720 1275.595 2914.100 1275.765 ;
        RECT 5.605 1274.845 6.815 1275.595 ;
        RECT 9.515 1274.935 9.855 1275.595 ;
        RECT 2906.365 1274.870 2906.655 1275.595 ;
        RECT 2912.805 1274.845 2914.015 1275.595 ;
        RECT 5.605 1274.305 6.125 1274.845 ;
        RECT 2913.495 1274.305 2914.015 1274.845 ;
        RECT 5.605 1271.075 6.125 1271.615 ;
        RECT 2913.495 1271.075 2914.015 1271.615 ;
        RECT 5.605 1270.325 6.815 1271.075 ;
        RECT 2912.805 1270.325 2914.015 1271.075 ;
        RECT 5.520 1270.155 6.900 1270.325 ;
        RECT 2906.300 1270.155 2906.740 1270.325 ;
        RECT 2912.720 1270.155 2914.100 1270.325 ;
        RECT 5.605 1269.405 6.815 1270.155 ;
        RECT 2906.365 1269.430 2906.655 1270.155 ;
        RECT 2912.805 1269.405 2914.015 1270.155 ;
        RECT 5.605 1268.865 6.125 1269.405 ;
        RECT 2913.495 1268.865 2914.015 1269.405 ;
        RECT 5.605 1265.635 6.125 1266.175 ;
        RECT 2913.495 1265.635 2914.015 1266.175 ;
        RECT 5.605 1264.885 6.815 1265.635 ;
        RECT 2909.815 1264.885 2910.155 1265.545 ;
        RECT 2912.805 1264.885 2914.015 1265.635 ;
        RECT 5.520 1264.715 6.900 1264.885 ;
        RECT 2906.300 1264.715 2906.740 1264.885 ;
        RECT 2909.040 1264.715 2910.420 1264.885 ;
        RECT 2912.720 1264.715 2914.100 1264.885 ;
        RECT 5.605 1263.965 6.815 1264.715 ;
        RECT 2906.365 1263.990 2906.655 1264.715 ;
        RECT 2912.805 1263.965 2914.015 1264.715 ;
        RECT 5.605 1263.425 6.125 1263.965 ;
        RECT 2913.495 1263.425 2914.015 1263.965 ;
        RECT 5.605 1260.195 6.125 1260.735 ;
        RECT 2913.495 1260.195 2914.015 1260.735 ;
        RECT 5.605 1259.445 6.815 1260.195 ;
        RECT 2912.805 1259.445 2914.015 1260.195 ;
        RECT 5.520 1259.275 6.900 1259.445 ;
        RECT 2906.300 1259.275 2906.740 1259.445 ;
        RECT 2912.720 1259.275 2914.100 1259.445 ;
        RECT 5.605 1258.525 6.815 1259.275 ;
        RECT 2906.365 1258.550 2906.655 1259.275 ;
        RECT 2912.805 1258.525 2914.015 1259.275 ;
        RECT 5.605 1257.985 6.125 1258.525 ;
        RECT 2913.495 1257.985 2914.015 1258.525 ;
        RECT 5.605 1254.755 6.125 1255.295 ;
        RECT 2913.495 1254.755 2914.015 1255.295 ;
        RECT 5.605 1254.005 6.815 1254.755 ;
        RECT 2912.805 1254.005 2914.015 1254.755 ;
        RECT 5.520 1253.835 6.900 1254.005 ;
        RECT 2906.300 1253.835 2906.740 1254.005 ;
        RECT 2912.720 1253.835 2914.100 1254.005 ;
        RECT 5.605 1253.085 6.815 1253.835 ;
        RECT 2906.365 1253.110 2906.655 1253.835 ;
        RECT 2912.805 1253.085 2914.015 1253.835 ;
        RECT 5.605 1252.545 6.125 1253.085 ;
        RECT 2913.495 1252.545 2914.015 1253.085 ;
        RECT 5.605 1249.315 6.125 1249.855 ;
        RECT 2913.495 1249.315 2914.015 1249.855 ;
        RECT 5.605 1248.565 6.815 1249.315 ;
        RECT 2912.805 1248.565 2914.015 1249.315 ;
        RECT 5.520 1248.395 6.900 1248.565 ;
        RECT 2906.300 1248.395 2906.740 1248.565 ;
        RECT 2912.720 1248.395 2914.100 1248.565 ;
        RECT 5.605 1247.645 6.815 1248.395 ;
        RECT 2906.365 1247.670 2906.655 1248.395 ;
        RECT 2912.805 1247.645 2914.015 1248.395 ;
        RECT 5.605 1247.105 6.125 1247.645 ;
        RECT 2913.495 1247.105 2914.015 1247.645 ;
        RECT 5.605 1243.875 6.125 1244.415 ;
        RECT 2913.495 1243.875 2914.015 1244.415 ;
        RECT 5.605 1243.125 6.815 1243.875 ;
        RECT 2912.805 1243.125 2914.015 1243.875 ;
        RECT 5.520 1242.955 6.900 1243.125 ;
        RECT 2912.720 1242.955 2914.100 1243.125 ;
        RECT 5.605 1242.205 6.815 1242.955 ;
        RECT 2912.805 1242.205 2914.015 1242.955 ;
        RECT 5.605 1241.665 6.125 1242.205 ;
        RECT 2913.495 1241.665 2914.015 1242.205 ;
        RECT 5.605 1238.435 6.125 1238.975 ;
        RECT 2913.495 1238.435 2914.015 1238.975 ;
        RECT 5.605 1237.685 6.815 1238.435 ;
        RECT 2910.045 1237.685 2910.335 1238.410 ;
        RECT 2912.805 1237.685 2914.015 1238.435 ;
        RECT 5.520 1237.515 6.900 1237.685 ;
        RECT 2909.960 1237.515 2910.420 1237.685 ;
        RECT 2912.720 1237.515 2914.100 1237.685 ;
        RECT 5.605 1236.765 6.815 1237.515 ;
        RECT 2912.805 1236.765 2914.015 1237.515 ;
        RECT 5.605 1236.225 6.125 1236.765 ;
        RECT 2913.495 1236.225 2914.015 1236.765 ;
        RECT 5.605 1232.995 6.125 1233.535 ;
        RECT 2913.495 1232.995 2914.015 1233.535 ;
        RECT 5.605 1232.245 6.815 1232.995 ;
        RECT 2910.045 1232.245 2910.335 1232.970 ;
        RECT 2912.805 1232.245 2914.015 1232.995 ;
        RECT 5.520 1232.075 6.900 1232.245 ;
        RECT 2909.960 1232.075 2910.420 1232.245 ;
        RECT 2912.720 1232.075 2914.100 1232.245 ;
        RECT 5.605 1231.325 6.815 1232.075 ;
        RECT 2912.805 1231.325 2914.015 1232.075 ;
        RECT 5.605 1230.785 6.125 1231.325 ;
        RECT 2913.495 1230.785 2914.015 1231.325 ;
        RECT 5.605 1227.555 6.125 1228.095 ;
        RECT 2913.495 1227.555 2914.015 1228.095 ;
        RECT 5.605 1226.805 6.815 1227.555 ;
        RECT 2910.045 1226.805 2910.335 1227.530 ;
        RECT 2912.805 1226.805 2914.015 1227.555 ;
        RECT 5.520 1226.635 6.900 1226.805 ;
        RECT 2909.960 1226.635 2910.420 1226.805 ;
        RECT 2912.720 1226.635 2914.100 1226.805 ;
        RECT 5.605 1225.885 6.815 1226.635 ;
        RECT 2912.805 1225.885 2914.015 1226.635 ;
        RECT 5.605 1225.345 6.125 1225.885 ;
        RECT 2913.495 1225.345 2914.015 1225.885 ;
        RECT 5.605 1222.115 6.125 1222.655 ;
        RECT 2913.495 1222.115 2914.015 1222.655 ;
        RECT 5.605 1221.365 6.815 1222.115 ;
        RECT 2910.045 1221.365 2910.335 1222.090 ;
        RECT 2912.805 1221.365 2914.015 1222.115 ;
        RECT 5.520 1221.195 6.900 1221.365 ;
        RECT 2909.960 1221.195 2910.420 1221.365 ;
        RECT 2912.720 1221.195 2914.100 1221.365 ;
        RECT 5.605 1220.445 6.815 1221.195 ;
        RECT 2912.805 1220.445 2914.015 1221.195 ;
        RECT 5.605 1219.905 6.125 1220.445 ;
        RECT 2913.495 1219.905 2914.015 1220.445 ;
        RECT 5.605 1216.675 6.125 1217.215 ;
        RECT 2913.495 1216.675 2914.015 1217.215 ;
        RECT 5.605 1215.925 6.815 1216.675 ;
        RECT 9.515 1215.925 9.855 1216.585 ;
        RECT 2910.045 1215.925 2910.335 1216.650 ;
        RECT 2912.805 1215.925 2914.015 1216.675 ;
        RECT 5.520 1215.755 6.900 1215.925 ;
        RECT 8.740 1215.755 10.120 1215.925 ;
        RECT 2909.960 1215.755 2910.420 1215.925 ;
        RECT 2912.720 1215.755 2914.100 1215.925 ;
        RECT 5.605 1215.005 6.815 1215.755 ;
        RECT 2912.805 1215.005 2914.015 1215.755 ;
        RECT 5.605 1214.465 6.125 1215.005 ;
        RECT 2913.495 1214.465 2914.015 1215.005 ;
        RECT 5.605 1211.235 6.125 1211.775 ;
        RECT 2913.495 1211.235 2914.015 1211.775 ;
        RECT 5.605 1210.485 6.815 1211.235 ;
        RECT 2910.045 1210.485 2910.335 1211.210 ;
        RECT 2912.805 1210.485 2914.015 1211.235 ;
        RECT 5.520 1210.315 6.900 1210.485 ;
        RECT 2909.960 1210.315 2910.420 1210.485 ;
        RECT 2912.720 1210.315 2914.100 1210.485 ;
        RECT 5.605 1209.565 6.815 1210.315 ;
        RECT 2912.805 1209.565 2914.015 1210.315 ;
        RECT 5.605 1209.025 6.125 1209.565 ;
        RECT 2913.495 1209.025 2914.015 1209.565 ;
        RECT 5.605 1205.795 6.125 1206.335 ;
        RECT 2913.495 1205.795 2914.015 1206.335 ;
        RECT 5.605 1205.045 6.815 1205.795 ;
        RECT 2910.045 1205.045 2910.335 1205.770 ;
        RECT 2912.805 1205.045 2914.015 1205.795 ;
        RECT 5.520 1204.875 6.900 1205.045 ;
        RECT 2909.960 1204.875 2910.420 1205.045 ;
        RECT 2912.720 1204.875 2914.100 1205.045 ;
        RECT 5.605 1204.125 6.815 1204.875 ;
        RECT 2912.805 1204.125 2914.015 1204.875 ;
        RECT 5.605 1203.585 6.125 1204.125 ;
        RECT 2913.495 1203.585 2914.015 1204.125 ;
        RECT 5.605 1200.355 6.125 1200.895 ;
        RECT 2913.495 1200.355 2914.015 1200.895 ;
        RECT 5.605 1199.605 6.815 1200.355 ;
        RECT 2910.045 1199.605 2910.335 1200.330 ;
        RECT 2912.805 1199.605 2914.015 1200.355 ;
        RECT 5.520 1199.435 6.900 1199.605 ;
        RECT 2909.960 1199.435 2910.420 1199.605 ;
        RECT 2912.720 1199.435 2914.100 1199.605 ;
        RECT 5.605 1198.685 6.815 1199.435 ;
        RECT 2912.805 1198.685 2914.015 1199.435 ;
        RECT 5.605 1198.145 6.125 1198.685 ;
        RECT 2913.495 1198.145 2914.015 1198.685 ;
        RECT 5.605 1194.915 6.125 1195.455 ;
        RECT 2913.495 1194.915 2914.015 1195.455 ;
        RECT 5.605 1194.165 6.815 1194.915 ;
        RECT 2910.045 1194.165 2910.335 1194.890 ;
        RECT 2912.805 1194.165 2914.015 1194.915 ;
        RECT 5.520 1193.995 6.900 1194.165 ;
        RECT 2909.960 1193.995 2910.420 1194.165 ;
        RECT 2912.720 1193.995 2914.100 1194.165 ;
        RECT 5.605 1193.245 6.815 1193.995 ;
        RECT 2912.805 1193.245 2914.015 1193.995 ;
        RECT 5.605 1192.705 6.125 1193.245 ;
        RECT 2913.495 1192.705 2914.015 1193.245 ;
        RECT 5.605 1189.475 6.125 1190.015 ;
        RECT 2913.495 1189.475 2914.015 1190.015 ;
        RECT 5.605 1188.725 6.815 1189.475 ;
        RECT 2910.045 1188.725 2910.335 1189.450 ;
        RECT 2912.805 1188.725 2914.015 1189.475 ;
        RECT 5.520 1188.555 6.900 1188.725 ;
        RECT 2909.960 1188.555 2910.420 1188.725 ;
        RECT 2912.720 1188.555 2914.100 1188.725 ;
        RECT 5.605 1187.805 6.815 1188.555 ;
        RECT 2912.805 1187.805 2914.015 1188.555 ;
        RECT 5.605 1187.265 6.125 1187.805 ;
        RECT 2913.495 1187.265 2914.015 1187.805 ;
        RECT 5.605 1184.035 6.125 1184.575 ;
        RECT 2913.495 1184.035 2914.015 1184.575 ;
        RECT 5.605 1183.285 6.815 1184.035 ;
        RECT 2910.045 1183.285 2910.335 1184.010 ;
        RECT 2912.805 1183.285 2914.015 1184.035 ;
        RECT 5.520 1183.115 6.900 1183.285 ;
        RECT 2909.960 1183.115 2910.420 1183.285 ;
        RECT 2912.720 1183.115 2914.100 1183.285 ;
        RECT 5.605 1182.365 6.815 1183.115 ;
        RECT 2912.805 1182.365 2914.015 1183.115 ;
        RECT 5.605 1181.825 6.125 1182.365 ;
        RECT 2913.495 1181.825 2914.015 1182.365 ;
        RECT 5.605 1178.595 6.125 1179.135 ;
        RECT 2913.495 1178.595 2914.015 1179.135 ;
        RECT 5.605 1177.845 6.815 1178.595 ;
        RECT 2910.045 1177.845 2910.335 1178.570 ;
        RECT 2912.805 1177.845 2914.015 1178.595 ;
        RECT 5.520 1177.675 6.900 1177.845 ;
        RECT 2909.960 1177.675 2910.420 1177.845 ;
        RECT 2912.720 1177.675 2914.100 1177.845 ;
        RECT 5.605 1176.925 6.815 1177.675 ;
        RECT 2912.805 1176.925 2914.015 1177.675 ;
        RECT 5.605 1176.385 6.125 1176.925 ;
        RECT 2913.495 1176.385 2914.015 1176.925 ;
        RECT 5.605 1173.155 6.125 1173.695 ;
        RECT 2913.495 1173.155 2914.015 1173.695 ;
        RECT 5.605 1172.405 6.815 1173.155 ;
        RECT 2910.045 1172.405 2910.335 1173.130 ;
        RECT 2912.805 1172.405 2914.015 1173.155 ;
        RECT 5.520 1172.235 6.900 1172.405 ;
        RECT 2909.960 1172.235 2910.420 1172.405 ;
        RECT 2912.720 1172.235 2914.100 1172.405 ;
        RECT 5.605 1171.485 6.815 1172.235 ;
        RECT 2912.805 1171.485 2914.015 1172.235 ;
        RECT 5.605 1170.945 6.125 1171.485 ;
        RECT 2913.495 1170.945 2914.015 1171.485 ;
        RECT 5.605 1167.715 6.125 1168.255 ;
        RECT 2913.495 1167.715 2914.015 1168.255 ;
        RECT 5.605 1166.965 6.815 1167.715 ;
        RECT 2910.045 1166.965 2910.335 1167.690 ;
        RECT 2912.805 1166.965 2914.015 1167.715 ;
        RECT 5.520 1166.795 6.900 1166.965 ;
        RECT 2909.960 1166.795 2910.420 1166.965 ;
        RECT 2912.720 1166.795 2914.100 1166.965 ;
        RECT 5.605 1166.045 6.815 1166.795 ;
        RECT 2912.805 1166.045 2914.015 1166.795 ;
        RECT 5.605 1165.505 6.125 1166.045 ;
        RECT 2913.495 1165.505 2914.015 1166.045 ;
        RECT 5.605 1162.275 6.125 1162.815 ;
        RECT 2913.495 1162.275 2914.015 1162.815 ;
        RECT 5.605 1161.525 6.815 1162.275 ;
        RECT 2910.045 1161.525 2910.335 1162.250 ;
        RECT 2912.805 1161.525 2914.015 1162.275 ;
        RECT 5.520 1161.355 6.900 1161.525 ;
        RECT 2909.960 1161.355 2910.420 1161.525 ;
        RECT 2912.720 1161.355 2914.100 1161.525 ;
        RECT 5.605 1160.605 6.815 1161.355 ;
        RECT 2912.805 1160.605 2914.015 1161.355 ;
        RECT 5.605 1160.065 6.125 1160.605 ;
        RECT 2913.495 1160.065 2914.015 1160.605 ;
        RECT 5.605 1156.835 6.125 1157.375 ;
        RECT 2913.495 1156.835 2914.015 1157.375 ;
        RECT 5.605 1156.085 6.815 1156.835 ;
        RECT 2910.045 1156.085 2910.335 1156.810 ;
        RECT 2912.805 1156.085 2914.015 1156.835 ;
        RECT 5.520 1155.915 6.900 1156.085 ;
        RECT 2909.960 1155.915 2910.420 1156.085 ;
        RECT 2912.720 1155.915 2914.100 1156.085 ;
        RECT 5.605 1155.165 6.815 1155.915 ;
        RECT 2912.805 1155.165 2914.015 1155.915 ;
        RECT 5.605 1154.625 6.125 1155.165 ;
        RECT 2913.495 1154.625 2914.015 1155.165 ;
        RECT 5.605 1151.395 6.125 1151.935 ;
        RECT 2913.495 1151.395 2914.015 1151.935 ;
        RECT 5.605 1150.645 6.815 1151.395 ;
        RECT 2910.045 1150.645 2910.335 1151.370 ;
        RECT 2912.805 1150.645 2914.015 1151.395 ;
        RECT 5.520 1150.475 6.900 1150.645 ;
        RECT 2909.960 1150.475 2910.420 1150.645 ;
        RECT 2912.720 1150.475 2914.100 1150.645 ;
        RECT 5.605 1149.725 6.815 1150.475 ;
        RECT 2912.805 1149.725 2914.015 1150.475 ;
        RECT 5.605 1149.185 6.125 1149.725 ;
        RECT 2913.495 1149.185 2914.015 1149.725 ;
        RECT 5.605 1145.955 6.125 1146.495 ;
        RECT 2913.495 1145.955 2914.015 1146.495 ;
        RECT 5.605 1145.205 6.815 1145.955 ;
        RECT 2910.045 1145.205 2910.335 1145.930 ;
        RECT 2912.805 1145.205 2914.015 1145.955 ;
        RECT 5.520 1145.035 6.900 1145.205 ;
        RECT 2909.960 1145.035 2910.420 1145.205 ;
        RECT 2912.720 1145.035 2914.100 1145.205 ;
        RECT 5.605 1144.285 6.815 1145.035 ;
        RECT 2912.805 1144.285 2914.015 1145.035 ;
        RECT 5.605 1143.745 6.125 1144.285 ;
        RECT 2913.495 1143.745 2914.015 1144.285 ;
        RECT 5.605 1140.515 6.125 1141.055 ;
        RECT 2913.495 1140.515 2914.015 1141.055 ;
        RECT 5.605 1139.765 6.815 1140.515 ;
        RECT 2910.045 1139.765 2910.335 1140.490 ;
        RECT 2912.805 1139.765 2914.015 1140.515 ;
        RECT 5.520 1139.595 6.900 1139.765 ;
        RECT 2909.960 1139.595 2910.420 1139.765 ;
        RECT 2912.720 1139.595 2914.100 1139.765 ;
        RECT 5.605 1138.845 6.815 1139.595 ;
        RECT 2912.805 1138.845 2914.015 1139.595 ;
        RECT 5.605 1138.305 6.125 1138.845 ;
        RECT 2913.495 1138.305 2914.015 1138.845 ;
        RECT 5.605 1135.075 6.125 1135.615 ;
        RECT 2913.495 1135.075 2914.015 1135.615 ;
        RECT 5.605 1134.325 6.815 1135.075 ;
        RECT 2910.045 1134.325 2910.335 1135.050 ;
        RECT 2912.805 1134.325 2914.015 1135.075 ;
        RECT 5.520 1134.155 6.900 1134.325 ;
        RECT 2909.960 1134.155 2910.420 1134.325 ;
        RECT 2912.720 1134.155 2914.100 1134.325 ;
        RECT 5.605 1133.405 6.815 1134.155 ;
        RECT 2912.805 1133.405 2914.015 1134.155 ;
        RECT 5.605 1132.865 6.125 1133.405 ;
        RECT 2913.495 1132.865 2914.015 1133.405 ;
        RECT 5.605 1129.635 6.125 1130.175 ;
        RECT 2913.495 1129.635 2914.015 1130.175 ;
        RECT 5.605 1128.885 6.815 1129.635 ;
        RECT 2910.045 1128.885 2910.335 1129.610 ;
        RECT 2912.805 1128.885 2914.015 1129.635 ;
        RECT 5.520 1128.715 6.900 1128.885 ;
        RECT 2909.960 1128.715 2910.420 1128.885 ;
        RECT 2912.720 1128.715 2914.100 1128.885 ;
        RECT 5.605 1127.965 6.815 1128.715 ;
        RECT 2912.805 1127.965 2914.015 1128.715 ;
        RECT 5.605 1127.425 6.125 1127.965 ;
        RECT 2913.495 1127.425 2914.015 1127.965 ;
        RECT 5.605 1124.195 6.125 1124.735 ;
        RECT 2913.495 1124.195 2914.015 1124.735 ;
        RECT 5.605 1123.445 6.815 1124.195 ;
        RECT 2910.045 1123.445 2910.335 1124.170 ;
        RECT 2912.805 1123.445 2914.015 1124.195 ;
        RECT 5.520 1123.275 6.900 1123.445 ;
        RECT 2909.960 1123.275 2910.420 1123.445 ;
        RECT 2912.720 1123.275 2914.100 1123.445 ;
        RECT 5.605 1122.525 6.815 1123.275 ;
        RECT 2912.805 1122.525 2914.015 1123.275 ;
        RECT 5.605 1121.985 6.125 1122.525 ;
        RECT 2913.495 1121.985 2914.015 1122.525 ;
        RECT 5.605 1118.755 6.125 1119.295 ;
        RECT 2913.495 1118.755 2914.015 1119.295 ;
        RECT 5.605 1118.005 6.815 1118.755 ;
        RECT 2910.045 1118.005 2910.335 1118.730 ;
        RECT 2912.805 1118.005 2914.015 1118.755 ;
        RECT 5.520 1117.835 6.900 1118.005 ;
        RECT 2909.960 1117.835 2910.420 1118.005 ;
        RECT 2912.720 1117.835 2914.100 1118.005 ;
        RECT 5.605 1117.085 6.815 1117.835 ;
        RECT 2912.805 1117.085 2914.015 1117.835 ;
        RECT 5.605 1116.545 6.125 1117.085 ;
        RECT 2913.495 1116.545 2914.015 1117.085 ;
        RECT 5.605 1113.315 6.125 1113.855 ;
        RECT 2913.495 1113.315 2914.015 1113.855 ;
        RECT 5.605 1112.565 6.815 1113.315 ;
        RECT 2910.045 1112.565 2910.335 1113.290 ;
        RECT 2912.805 1112.565 2914.015 1113.315 ;
        RECT 5.520 1112.395 6.900 1112.565 ;
        RECT 8.740 1112.395 10.120 1112.565 ;
        RECT 2909.960 1112.395 2910.420 1112.565 ;
        RECT 2912.720 1112.395 2914.100 1112.565 ;
        RECT 5.605 1111.645 6.815 1112.395 ;
        RECT 9.515 1111.735 9.855 1112.395 ;
        RECT 2912.805 1111.645 2914.015 1112.395 ;
        RECT 5.605 1111.105 6.125 1111.645 ;
        RECT 2913.495 1111.105 2914.015 1111.645 ;
        RECT 5.605 1107.875 6.125 1108.415 ;
        RECT 2913.495 1107.875 2914.015 1108.415 ;
        RECT 5.605 1107.125 6.815 1107.875 ;
        RECT 2910.045 1107.125 2910.335 1107.850 ;
        RECT 2912.805 1107.125 2914.015 1107.875 ;
        RECT 5.520 1106.955 6.900 1107.125 ;
        RECT 2909.960 1106.955 2910.420 1107.125 ;
        RECT 2912.720 1106.955 2914.100 1107.125 ;
        RECT 5.605 1106.205 6.815 1106.955 ;
        RECT 2912.805 1106.205 2914.015 1106.955 ;
        RECT 5.605 1105.665 6.125 1106.205 ;
        RECT 2913.495 1105.665 2914.015 1106.205 ;
        RECT 5.605 1102.435 6.125 1102.975 ;
        RECT 2913.495 1102.435 2914.015 1102.975 ;
        RECT 5.605 1101.685 6.815 1102.435 ;
        RECT 2910.045 1101.685 2910.335 1102.410 ;
        RECT 2912.805 1101.685 2914.015 1102.435 ;
        RECT 5.520 1101.515 6.900 1101.685 ;
        RECT 2909.960 1101.515 2910.420 1101.685 ;
        RECT 2912.720 1101.515 2914.100 1101.685 ;
        RECT 5.605 1100.765 6.815 1101.515 ;
        RECT 2912.805 1100.765 2914.015 1101.515 ;
        RECT 5.605 1100.225 6.125 1100.765 ;
        RECT 2913.495 1100.225 2914.015 1100.765 ;
        RECT 5.605 1096.995 6.125 1097.535 ;
        RECT 2913.495 1096.995 2914.015 1097.535 ;
        RECT 5.605 1096.245 6.815 1096.995 ;
        RECT 2910.045 1096.245 2910.335 1096.970 ;
        RECT 2912.805 1096.245 2914.015 1096.995 ;
        RECT 5.520 1096.075 6.900 1096.245 ;
        RECT 2909.960 1096.075 2910.420 1096.245 ;
        RECT 2912.720 1096.075 2914.100 1096.245 ;
        RECT 5.605 1095.325 6.815 1096.075 ;
        RECT 2912.805 1095.325 2914.015 1096.075 ;
        RECT 5.605 1094.785 6.125 1095.325 ;
        RECT 2913.495 1094.785 2914.015 1095.325 ;
        RECT 5.605 1091.555 6.125 1092.095 ;
        RECT 2913.495 1091.555 2914.015 1092.095 ;
        RECT 5.605 1090.805 6.815 1091.555 ;
        RECT 2910.045 1090.805 2910.335 1091.530 ;
        RECT 2912.805 1090.805 2914.015 1091.555 ;
        RECT 5.520 1090.635 6.900 1090.805 ;
        RECT 2909.960 1090.635 2910.420 1090.805 ;
        RECT 2912.720 1090.635 2914.100 1090.805 ;
        RECT 5.605 1089.885 6.815 1090.635 ;
        RECT 2912.805 1089.885 2914.015 1090.635 ;
        RECT 5.605 1089.345 6.125 1089.885 ;
        RECT 2913.495 1089.345 2914.015 1089.885 ;
        RECT 5.605 1086.115 6.125 1086.655 ;
        RECT 2913.495 1086.115 2914.015 1086.655 ;
        RECT 5.605 1085.365 6.815 1086.115 ;
        RECT 2910.045 1085.365 2910.335 1086.090 ;
        RECT 2912.805 1085.365 2914.015 1086.115 ;
        RECT 5.520 1085.195 6.900 1085.365 ;
        RECT 2909.960 1085.195 2910.420 1085.365 ;
        RECT 2912.720 1085.195 2914.100 1085.365 ;
        RECT 5.605 1084.445 6.815 1085.195 ;
        RECT 2912.805 1084.445 2914.015 1085.195 ;
        RECT 5.605 1083.905 6.125 1084.445 ;
        RECT 2913.495 1083.905 2914.015 1084.445 ;
        RECT 5.605 1080.675 6.125 1081.215 ;
        RECT 2913.495 1080.675 2914.015 1081.215 ;
        RECT 5.605 1079.925 6.815 1080.675 ;
        RECT 2910.045 1079.925 2910.335 1080.650 ;
        RECT 2912.805 1079.925 2914.015 1080.675 ;
        RECT 5.520 1079.755 6.900 1079.925 ;
        RECT 2909.960 1079.755 2910.420 1079.925 ;
        RECT 2912.720 1079.755 2914.100 1079.925 ;
        RECT 5.605 1079.005 6.815 1079.755 ;
        RECT 2912.805 1079.005 2914.015 1079.755 ;
        RECT 5.605 1078.465 6.125 1079.005 ;
        RECT 2913.495 1078.465 2914.015 1079.005 ;
        RECT 5.605 1075.235 6.125 1075.775 ;
        RECT 2913.495 1075.235 2914.015 1075.775 ;
        RECT 5.605 1074.485 6.815 1075.235 ;
        RECT 2910.045 1074.485 2910.335 1075.210 ;
        RECT 2912.805 1074.485 2914.015 1075.235 ;
        RECT 5.520 1074.315 6.900 1074.485 ;
        RECT 2909.960 1074.315 2910.420 1074.485 ;
        RECT 2912.720 1074.315 2914.100 1074.485 ;
        RECT 5.605 1073.565 6.815 1074.315 ;
        RECT 2912.805 1073.565 2914.015 1074.315 ;
        RECT 5.605 1073.025 6.125 1073.565 ;
        RECT 2913.495 1073.025 2914.015 1073.565 ;
        RECT 5.605 1069.795 6.125 1070.335 ;
        RECT 2913.495 1069.795 2914.015 1070.335 ;
        RECT 5.605 1069.045 6.815 1069.795 ;
        RECT 2910.045 1069.045 2910.335 1069.770 ;
        RECT 2912.805 1069.045 2914.015 1069.795 ;
        RECT 5.520 1068.875 6.900 1069.045 ;
        RECT 2909.960 1068.875 2910.420 1069.045 ;
        RECT 2912.720 1068.875 2914.100 1069.045 ;
        RECT 5.605 1068.125 6.815 1068.875 ;
        RECT 2912.805 1068.125 2914.015 1068.875 ;
        RECT 5.605 1067.585 6.125 1068.125 ;
        RECT 2913.495 1067.585 2914.015 1068.125 ;
        RECT 5.605 1064.355 6.125 1064.895 ;
        RECT 2913.495 1064.355 2914.015 1064.895 ;
        RECT 5.605 1063.605 6.815 1064.355 ;
        RECT 2910.045 1063.605 2910.335 1064.330 ;
        RECT 2912.805 1063.605 2914.015 1064.355 ;
        RECT 5.520 1063.435 6.900 1063.605 ;
        RECT 2909.960 1063.435 2910.420 1063.605 ;
        RECT 2912.720 1063.435 2914.100 1063.605 ;
        RECT 5.605 1062.685 6.815 1063.435 ;
        RECT 2912.805 1062.685 2914.015 1063.435 ;
        RECT 5.605 1062.145 6.125 1062.685 ;
        RECT 2913.495 1062.145 2914.015 1062.685 ;
        RECT 5.605 1058.915 6.125 1059.455 ;
        RECT 2913.495 1058.915 2914.015 1059.455 ;
        RECT 5.605 1058.165 6.815 1058.915 ;
        RECT 2910.045 1058.165 2910.335 1058.890 ;
        RECT 2912.805 1058.165 2914.015 1058.915 ;
        RECT 5.520 1057.995 6.900 1058.165 ;
        RECT 2909.960 1057.995 2910.420 1058.165 ;
        RECT 2912.720 1057.995 2914.100 1058.165 ;
        RECT 5.605 1057.245 6.815 1057.995 ;
        RECT 2912.805 1057.245 2914.015 1057.995 ;
        RECT 5.605 1056.705 6.125 1057.245 ;
        RECT 2913.495 1056.705 2914.015 1057.245 ;
        RECT 5.605 1053.475 6.125 1054.015 ;
        RECT 2913.495 1053.475 2914.015 1054.015 ;
        RECT 5.605 1052.725 6.815 1053.475 ;
        RECT 2910.045 1052.725 2910.335 1053.450 ;
        RECT 2912.805 1052.725 2914.015 1053.475 ;
        RECT 5.520 1052.555 6.900 1052.725 ;
        RECT 2909.960 1052.555 2910.420 1052.725 ;
        RECT 2912.720 1052.555 2914.100 1052.725 ;
        RECT 5.605 1051.805 6.815 1052.555 ;
        RECT 2912.805 1051.805 2914.015 1052.555 ;
        RECT 5.605 1051.265 6.125 1051.805 ;
        RECT 2913.495 1051.265 2914.015 1051.805 ;
        RECT 5.605 1048.035 6.125 1048.575 ;
        RECT 2913.495 1048.035 2914.015 1048.575 ;
        RECT 5.605 1047.285 6.815 1048.035 ;
        RECT 2910.045 1047.285 2910.335 1048.010 ;
        RECT 2912.805 1047.285 2914.015 1048.035 ;
        RECT 5.520 1047.115 6.900 1047.285 ;
        RECT 2909.960 1047.115 2910.420 1047.285 ;
        RECT 2912.720 1047.115 2914.100 1047.285 ;
        RECT 5.605 1046.365 6.815 1047.115 ;
        RECT 2912.805 1046.365 2914.015 1047.115 ;
        RECT 5.605 1045.825 6.125 1046.365 ;
        RECT 2913.495 1045.825 2914.015 1046.365 ;
        RECT 5.605 1042.595 6.125 1043.135 ;
        RECT 2913.495 1042.595 2914.015 1043.135 ;
        RECT 5.605 1041.845 6.815 1042.595 ;
        RECT 2910.045 1041.845 2910.335 1042.570 ;
        RECT 2912.805 1041.845 2914.015 1042.595 ;
        RECT 5.520 1041.675 6.900 1041.845 ;
        RECT 2909.960 1041.675 2910.420 1041.845 ;
        RECT 2912.720 1041.675 2914.100 1041.845 ;
        RECT 5.605 1040.925 6.815 1041.675 ;
        RECT 2912.805 1040.925 2914.015 1041.675 ;
        RECT 5.605 1040.385 6.125 1040.925 ;
        RECT 2913.495 1040.385 2914.015 1040.925 ;
        RECT 5.605 1037.155 6.125 1037.695 ;
        RECT 2913.495 1037.155 2914.015 1037.695 ;
        RECT 5.605 1036.405 6.815 1037.155 ;
        RECT 2910.045 1036.405 2910.335 1037.130 ;
        RECT 2912.805 1036.405 2914.015 1037.155 ;
        RECT 5.520 1036.235 6.900 1036.405 ;
        RECT 8.740 1036.235 10.120 1036.405 ;
        RECT 2909.960 1036.235 2910.420 1036.405 ;
        RECT 2912.720 1036.235 2914.100 1036.405 ;
        RECT 5.605 1035.485 6.815 1036.235 ;
        RECT 9.515 1035.575 9.855 1036.235 ;
        RECT 2912.805 1035.485 2914.015 1036.235 ;
        RECT 5.605 1034.945 6.125 1035.485 ;
        RECT 2913.495 1034.945 2914.015 1035.485 ;
        RECT 5.605 1031.715 6.125 1032.255 ;
        RECT 2913.495 1031.715 2914.015 1032.255 ;
        RECT 5.605 1030.965 6.815 1031.715 ;
        RECT 2910.045 1030.965 2910.335 1031.690 ;
        RECT 2912.805 1030.965 2914.015 1031.715 ;
        RECT 5.520 1030.795 6.900 1030.965 ;
        RECT 2909.960 1030.795 2910.420 1030.965 ;
        RECT 2912.720 1030.795 2914.100 1030.965 ;
        RECT 5.605 1030.045 6.815 1030.795 ;
        RECT 2912.805 1030.045 2914.015 1030.795 ;
        RECT 5.605 1029.505 6.125 1030.045 ;
        RECT 2913.495 1029.505 2914.015 1030.045 ;
        RECT 5.605 1026.275 6.125 1026.815 ;
        RECT 2913.495 1026.275 2914.015 1026.815 ;
        RECT 5.605 1025.525 6.815 1026.275 ;
        RECT 2910.045 1025.525 2910.335 1026.250 ;
        RECT 2912.805 1025.525 2914.015 1026.275 ;
        RECT 5.520 1025.355 6.900 1025.525 ;
        RECT 2909.960 1025.355 2910.420 1025.525 ;
        RECT 2912.720 1025.355 2914.100 1025.525 ;
        RECT 5.605 1024.605 6.815 1025.355 ;
        RECT 2912.805 1024.605 2914.015 1025.355 ;
        RECT 5.605 1024.065 6.125 1024.605 ;
        RECT 2913.495 1024.065 2914.015 1024.605 ;
        RECT 5.605 1020.835 6.125 1021.375 ;
        RECT 2913.495 1020.835 2914.015 1021.375 ;
        RECT 5.605 1020.085 6.815 1020.835 ;
        RECT 2910.045 1020.085 2910.335 1020.810 ;
        RECT 2912.805 1020.085 2914.015 1020.835 ;
        RECT 5.520 1019.915 6.900 1020.085 ;
        RECT 2909.960 1019.915 2910.420 1020.085 ;
        RECT 2912.720 1019.915 2914.100 1020.085 ;
        RECT 5.605 1019.165 6.815 1019.915 ;
        RECT 2912.805 1019.165 2914.015 1019.915 ;
        RECT 5.605 1018.625 6.125 1019.165 ;
        RECT 2913.495 1018.625 2914.015 1019.165 ;
        RECT 5.605 1015.395 6.125 1015.935 ;
        RECT 2913.495 1015.395 2914.015 1015.935 ;
        RECT 5.605 1014.645 6.815 1015.395 ;
        RECT 2910.045 1014.645 2910.335 1015.370 ;
        RECT 2912.805 1014.645 2914.015 1015.395 ;
        RECT 5.520 1014.475 6.900 1014.645 ;
        RECT 2909.960 1014.475 2910.420 1014.645 ;
        RECT 2912.720 1014.475 2914.100 1014.645 ;
        RECT 5.605 1013.725 6.815 1014.475 ;
        RECT 2912.805 1013.725 2914.015 1014.475 ;
        RECT 5.605 1013.185 6.125 1013.725 ;
        RECT 2913.495 1013.185 2914.015 1013.725 ;
        RECT 5.605 1009.955 6.125 1010.495 ;
        RECT 2913.495 1009.955 2914.015 1010.495 ;
        RECT 5.605 1009.205 6.815 1009.955 ;
        RECT 2910.045 1009.205 2910.335 1009.930 ;
        RECT 2912.805 1009.205 2914.015 1009.955 ;
        RECT 5.520 1009.035 6.900 1009.205 ;
        RECT 2909.040 1009.035 2910.420 1009.205 ;
        RECT 2912.720 1009.035 2914.100 1009.205 ;
        RECT 5.605 1008.285 6.815 1009.035 ;
        RECT 2909.815 1008.375 2910.155 1009.035 ;
        RECT 2912.805 1008.285 2914.015 1009.035 ;
        RECT 5.605 1007.745 6.125 1008.285 ;
        RECT 2913.495 1007.745 2914.015 1008.285 ;
        RECT 5.605 1004.515 6.125 1005.055 ;
        RECT 2913.495 1004.515 2914.015 1005.055 ;
        RECT 5.605 1003.765 6.815 1004.515 ;
        RECT 2910.045 1003.765 2910.335 1004.490 ;
        RECT 2912.805 1003.765 2914.015 1004.515 ;
        RECT 5.520 1003.595 6.900 1003.765 ;
        RECT 2909.960 1003.595 2910.420 1003.765 ;
        RECT 2912.720 1003.595 2914.100 1003.765 ;
        RECT 5.605 1002.845 6.815 1003.595 ;
        RECT 2912.805 1002.845 2914.015 1003.595 ;
        RECT 5.605 1002.305 6.125 1002.845 ;
        RECT 2913.495 1002.305 2914.015 1002.845 ;
        RECT 5.605 999.075 6.125 999.615 ;
        RECT 2913.495 999.075 2914.015 999.615 ;
        RECT 5.605 998.325 6.815 999.075 ;
        RECT 2910.045 998.325 2910.335 999.050 ;
        RECT 2912.805 998.325 2914.015 999.075 ;
        RECT 5.520 998.155 6.900 998.325 ;
        RECT 2909.040 998.155 2910.420 998.325 ;
        RECT 2912.720 998.155 2914.100 998.325 ;
        RECT 5.605 997.405 6.815 998.155 ;
        RECT 2909.815 997.495 2910.155 998.155 ;
        RECT 2912.805 997.405 2914.015 998.155 ;
        RECT 5.605 996.865 6.125 997.405 ;
        RECT 2913.495 996.865 2914.015 997.405 ;
        RECT 5.605 993.635 6.125 994.175 ;
        RECT 2913.495 993.635 2914.015 994.175 ;
        RECT 5.605 992.885 6.815 993.635 ;
        RECT 2910.045 992.885 2910.335 993.610 ;
        RECT 2912.805 992.885 2914.015 993.635 ;
        RECT 5.520 992.715 6.900 992.885 ;
        RECT 2909.960 992.715 2910.420 992.885 ;
        RECT 2912.720 992.715 2914.100 992.885 ;
        RECT 5.605 991.965 6.815 992.715 ;
        RECT 2912.805 991.965 2914.015 992.715 ;
        RECT 5.605 991.425 6.125 991.965 ;
        RECT 2913.495 991.425 2914.015 991.965 ;
        RECT 5.605 988.195 6.125 988.735 ;
        RECT 2913.495 988.195 2914.015 988.735 ;
        RECT 5.605 987.445 6.815 988.195 ;
        RECT 2910.045 987.445 2910.335 988.170 ;
        RECT 2912.805 987.445 2914.015 988.195 ;
        RECT 5.520 987.275 6.900 987.445 ;
        RECT 2909.960 987.275 2910.420 987.445 ;
        RECT 2912.720 987.275 2914.100 987.445 ;
        RECT 5.605 986.525 6.815 987.275 ;
        RECT 2912.805 986.525 2914.015 987.275 ;
        RECT 5.605 985.985 6.125 986.525 ;
        RECT 2913.495 985.985 2914.015 986.525 ;
        RECT 5.605 982.755 6.125 983.295 ;
        RECT 2913.495 982.755 2914.015 983.295 ;
        RECT 5.605 982.005 6.815 982.755 ;
        RECT 2910.045 982.005 2910.335 982.730 ;
        RECT 2912.805 982.005 2914.015 982.755 ;
        RECT 5.520 981.835 6.900 982.005 ;
        RECT 2909.960 981.835 2910.420 982.005 ;
        RECT 2912.720 981.835 2914.100 982.005 ;
        RECT 5.605 981.085 6.815 981.835 ;
        RECT 2912.805 981.085 2914.015 981.835 ;
        RECT 5.605 980.545 6.125 981.085 ;
        RECT 2913.495 980.545 2914.015 981.085 ;
        RECT 5.605 977.315 6.125 977.855 ;
        RECT 2913.495 977.315 2914.015 977.855 ;
        RECT 5.605 976.565 6.815 977.315 ;
        RECT 2910.045 976.565 2910.335 977.290 ;
        RECT 2912.805 976.565 2914.015 977.315 ;
        RECT 5.520 976.395 6.900 976.565 ;
        RECT 2909.960 976.395 2910.420 976.565 ;
        RECT 2912.720 976.395 2914.100 976.565 ;
        RECT 5.605 975.645 6.815 976.395 ;
        RECT 2912.805 975.645 2914.015 976.395 ;
        RECT 5.605 975.105 6.125 975.645 ;
        RECT 2913.495 975.105 2914.015 975.645 ;
        RECT 5.605 971.875 6.125 972.415 ;
        RECT 2913.495 971.875 2914.015 972.415 ;
        RECT 5.605 971.125 6.815 971.875 ;
        RECT 2910.045 971.125 2910.335 971.850 ;
        RECT 2912.805 971.125 2914.015 971.875 ;
        RECT 5.520 970.955 6.900 971.125 ;
        RECT 2909.960 970.955 2910.420 971.125 ;
        RECT 2912.720 970.955 2914.100 971.125 ;
        RECT 5.605 970.205 6.815 970.955 ;
        RECT 2912.805 970.205 2914.015 970.955 ;
        RECT 5.605 969.665 6.125 970.205 ;
        RECT 2913.495 969.665 2914.015 970.205 ;
        RECT 5.605 966.435 6.125 966.975 ;
        RECT 2913.495 966.435 2914.015 966.975 ;
        RECT 5.605 965.685 6.815 966.435 ;
        RECT 2910.045 965.685 2910.335 966.410 ;
        RECT 2912.805 965.685 2914.015 966.435 ;
        RECT 5.520 965.515 6.900 965.685 ;
        RECT 2909.960 965.515 2910.420 965.685 ;
        RECT 2912.720 965.515 2914.100 965.685 ;
        RECT 5.605 964.765 6.815 965.515 ;
        RECT 2912.805 964.765 2914.015 965.515 ;
        RECT 5.605 964.225 6.125 964.765 ;
        RECT 2913.495 964.225 2914.015 964.765 ;
        RECT 5.605 960.995 6.125 961.535 ;
        RECT 2913.495 960.995 2914.015 961.535 ;
        RECT 5.605 960.245 6.815 960.995 ;
        RECT 2910.045 960.245 2910.335 960.970 ;
        RECT 2912.805 960.245 2914.015 960.995 ;
        RECT 5.520 960.075 6.900 960.245 ;
        RECT 2909.960 960.075 2910.420 960.245 ;
        RECT 2912.720 960.075 2914.100 960.245 ;
        RECT 5.605 959.325 6.815 960.075 ;
        RECT 2912.805 959.325 2914.015 960.075 ;
        RECT 5.605 958.785 6.125 959.325 ;
        RECT 2913.495 958.785 2914.015 959.325 ;
        RECT 5.605 955.555 6.125 956.095 ;
        RECT 2913.495 955.555 2914.015 956.095 ;
        RECT 5.605 954.805 6.815 955.555 ;
        RECT 2910.045 954.805 2910.335 955.530 ;
        RECT 2912.805 954.805 2914.015 955.555 ;
        RECT 5.520 954.635 6.900 954.805 ;
        RECT 2909.960 954.635 2910.420 954.805 ;
        RECT 2912.720 954.635 2914.100 954.805 ;
        RECT 5.605 953.885 6.815 954.635 ;
        RECT 2912.805 953.885 2914.015 954.635 ;
        RECT 5.605 953.345 6.125 953.885 ;
        RECT 2913.495 953.345 2914.015 953.885 ;
        RECT 5.605 950.115 6.125 950.655 ;
        RECT 2913.495 950.115 2914.015 950.655 ;
        RECT 5.605 949.365 6.815 950.115 ;
        RECT 2910.045 949.365 2910.335 950.090 ;
        RECT 2912.805 949.365 2914.015 950.115 ;
        RECT 5.520 949.195 6.900 949.365 ;
        RECT 2909.960 949.195 2910.420 949.365 ;
        RECT 2912.720 949.195 2914.100 949.365 ;
        RECT 5.605 948.445 6.815 949.195 ;
        RECT 2912.805 948.445 2914.015 949.195 ;
        RECT 5.605 947.905 6.125 948.445 ;
        RECT 2913.495 947.905 2914.015 948.445 ;
        RECT 5.605 944.675 6.125 945.215 ;
        RECT 2913.495 944.675 2914.015 945.215 ;
        RECT 5.605 943.925 6.815 944.675 ;
        RECT 2910.045 943.925 2910.335 944.650 ;
        RECT 2912.805 943.925 2914.015 944.675 ;
        RECT 5.520 943.755 6.900 943.925 ;
        RECT 2909.960 943.755 2910.420 943.925 ;
        RECT 2912.720 943.755 2914.100 943.925 ;
        RECT 5.605 943.005 6.815 943.755 ;
        RECT 2912.805 943.005 2914.015 943.755 ;
        RECT 5.605 942.465 6.125 943.005 ;
        RECT 2913.495 942.465 2914.015 943.005 ;
        RECT 5.605 939.235 6.125 939.775 ;
        RECT 2913.495 939.235 2914.015 939.775 ;
        RECT 5.605 938.485 6.815 939.235 ;
        RECT 2910.045 938.485 2910.335 939.210 ;
        RECT 2912.805 938.485 2914.015 939.235 ;
        RECT 5.520 938.315 6.900 938.485 ;
        RECT 2909.960 938.315 2910.420 938.485 ;
        RECT 2912.720 938.315 2914.100 938.485 ;
        RECT 5.605 937.565 6.815 938.315 ;
        RECT 2912.805 937.565 2914.015 938.315 ;
        RECT 5.605 937.025 6.125 937.565 ;
        RECT 2913.495 937.025 2914.015 937.565 ;
        RECT 5.605 933.795 6.125 934.335 ;
        RECT 2913.495 933.795 2914.015 934.335 ;
        RECT 5.605 933.045 6.815 933.795 ;
        RECT 2910.045 933.045 2910.335 933.770 ;
        RECT 2912.805 933.045 2914.015 933.795 ;
        RECT 5.520 932.875 6.900 933.045 ;
        RECT 2909.960 932.875 2910.420 933.045 ;
        RECT 2912.720 932.875 2914.100 933.045 ;
        RECT 5.605 932.125 6.815 932.875 ;
        RECT 2912.805 932.125 2914.015 932.875 ;
        RECT 5.605 931.585 6.125 932.125 ;
        RECT 2913.495 931.585 2914.015 932.125 ;
        RECT 5.605 928.355 6.125 928.895 ;
        RECT 2913.495 928.355 2914.015 928.895 ;
        RECT 5.605 927.605 6.815 928.355 ;
        RECT 2910.045 927.605 2910.335 928.330 ;
        RECT 2912.805 927.605 2914.015 928.355 ;
        RECT 5.520 927.435 6.900 927.605 ;
        RECT 2909.960 927.435 2910.420 927.605 ;
        RECT 2912.720 927.435 2914.100 927.605 ;
        RECT 5.605 926.685 6.815 927.435 ;
        RECT 2912.805 926.685 2914.015 927.435 ;
        RECT 5.605 926.145 6.125 926.685 ;
        RECT 2913.495 926.145 2914.015 926.685 ;
        RECT 5.605 922.915 6.125 923.455 ;
        RECT 2913.495 922.915 2914.015 923.455 ;
        RECT 5.605 922.165 6.815 922.915 ;
        RECT 2910.045 922.165 2910.335 922.890 ;
        RECT 2912.805 922.165 2914.015 922.915 ;
        RECT 5.520 921.995 6.900 922.165 ;
        RECT 2909.960 921.995 2910.420 922.165 ;
        RECT 2912.720 921.995 2914.100 922.165 ;
        RECT 5.605 921.245 6.815 921.995 ;
        RECT 2912.805 921.245 2914.015 921.995 ;
        RECT 5.605 920.705 6.125 921.245 ;
        RECT 2913.495 920.705 2914.015 921.245 ;
        RECT 5.605 917.475 6.125 918.015 ;
        RECT 2913.495 917.475 2914.015 918.015 ;
        RECT 5.605 916.725 6.815 917.475 ;
        RECT 2910.045 916.725 2910.335 917.450 ;
        RECT 2912.805 916.725 2914.015 917.475 ;
        RECT 5.520 916.555 6.900 916.725 ;
        RECT 2909.960 916.555 2910.420 916.725 ;
        RECT 2912.720 916.555 2914.100 916.725 ;
        RECT 5.605 915.805 6.815 916.555 ;
        RECT 2912.805 915.805 2914.015 916.555 ;
        RECT 5.605 915.265 6.125 915.805 ;
        RECT 2913.495 915.265 2914.015 915.805 ;
        RECT 5.605 912.035 6.125 912.575 ;
        RECT 2913.495 912.035 2914.015 912.575 ;
        RECT 5.605 911.285 6.815 912.035 ;
        RECT 2910.045 911.285 2910.335 912.010 ;
        RECT 2912.805 911.285 2914.015 912.035 ;
        RECT 5.520 911.115 6.900 911.285 ;
        RECT 2909.960 911.115 2910.420 911.285 ;
        RECT 2912.720 911.115 2914.100 911.285 ;
        RECT 5.605 910.365 6.815 911.115 ;
        RECT 2912.805 910.365 2914.015 911.115 ;
        RECT 5.605 909.825 6.125 910.365 ;
        RECT 2913.495 909.825 2914.015 910.365 ;
        RECT 5.605 906.595 6.125 907.135 ;
        RECT 2913.495 906.595 2914.015 907.135 ;
        RECT 5.605 905.845 6.815 906.595 ;
        RECT 2910.045 905.845 2910.335 906.570 ;
        RECT 2912.805 905.845 2914.015 906.595 ;
        RECT 5.520 905.675 6.900 905.845 ;
        RECT 2909.960 905.675 2910.420 905.845 ;
        RECT 2912.720 905.675 2914.100 905.845 ;
        RECT 5.605 904.925 6.815 905.675 ;
        RECT 2912.805 904.925 2914.015 905.675 ;
        RECT 5.605 904.385 6.125 904.925 ;
        RECT 2913.495 904.385 2914.015 904.925 ;
        RECT 5.605 901.155 6.125 901.695 ;
        RECT 2913.495 901.155 2914.015 901.695 ;
        RECT 5.605 900.405 6.815 901.155 ;
        RECT 2910.045 900.405 2910.335 901.130 ;
        RECT 2912.805 900.405 2914.015 901.155 ;
        RECT 5.520 900.235 6.900 900.405 ;
        RECT 2909.960 900.235 2910.420 900.405 ;
        RECT 2912.720 900.235 2914.100 900.405 ;
        RECT 5.605 899.485 6.815 900.235 ;
        RECT 2912.805 899.485 2914.015 900.235 ;
        RECT 5.605 898.945 6.125 899.485 ;
        RECT 2913.495 898.945 2914.015 899.485 ;
        RECT 5.605 895.715 6.125 896.255 ;
        RECT 2913.495 895.715 2914.015 896.255 ;
        RECT 5.605 894.965 6.815 895.715 ;
        RECT 2910.045 894.965 2910.335 895.690 ;
        RECT 2912.805 894.965 2914.015 895.715 ;
        RECT 5.520 894.795 6.900 894.965 ;
        RECT 2909.960 894.795 2910.420 894.965 ;
        RECT 2912.720 894.795 2914.100 894.965 ;
        RECT 5.605 894.045 6.815 894.795 ;
        RECT 2912.805 894.045 2914.015 894.795 ;
        RECT 5.605 893.505 6.125 894.045 ;
        RECT 2913.495 893.505 2914.015 894.045 ;
        RECT 5.605 890.275 6.125 890.815 ;
        RECT 2913.495 890.275 2914.015 890.815 ;
        RECT 5.605 889.525 6.815 890.275 ;
        RECT 2910.045 889.525 2910.335 890.250 ;
        RECT 2912.805 889.525 2914.015 890.275 ;
        RECT 5.520 889.355 6.900 889.525 ;
        RECT 2909.960 889.355 2910.420 889.525 ;
        RECT 2912.720 889.355 2914.100 889.525 ;
        RECT 5.605 888.605 6.815 889.355 ;
        RECT 2912.805 888.605 2914.015 889.355 ;
        RECT 5.605 888.065 6.125 888.605 ;
        RECT 2913.495 888.065 2914.015 888.605 ;
        RECT 5.605 884.835 6.125 885.375 ;
        RECT 2913.495 884.835 2914.015 885.375 ;
        RECT 5.605 884.085 6.815 884.835 ;
        RECT 2910.045 884.085 2910.335 884.810 ;
        RECT 2912.805 884.085 2914.015 884.835 ;
        RECT 5.520 883.915 6.900 884.085 ;
        RECT 2909.960 883.915 2910.420 884.085 ;
        RECT 2912.720 883.915 2914.100 884.085 ;
        RECT 5.605 883.165 6.815 883.915 ;
        RECT 2912.805 883.165 2914.015 883.915 ;
        RECT 5.605 882.625 6.125 883.165 ;
        RECT 2913.495 882.625 2914.015 883.165 ;
        RECT 5.605 879.395 6.125 879.935 ;
        RECT 2913.495 879.395 2914.015 879.935 ;
        RECT 5.605 878.645 6.815 879.395 ;
        RECT 2910.045 878.645 2910.335 879.370 ;
        RECT 2912.805 878.645 2914.015 879.395 ;
        RECT 5.520 878.475 6.900 878.645 ;
        RECT 2909.960 878.475 2910.420 878.645 ;
        RECT 2912.720 878.475 2914.100 878.645 ;
        RECT 5.605 877.725 6.815 878.475 ;
        RECT 2912.805 877.725 2914.015 878.475 ;
        RECT 5.605 877.185 6.125 877.725 ;
        RECT 2913.495 877.185 2914.015 877.725 ;
        RECT 5.605 873.955 6.125 874.495 ;
        RECT 2913.495 873.955 2914.015 874.495 ;
        RECT 5.605 873.205 6.815 873.955 ;
        RECT 2910.045 873.205 2910.335 873.930 ;
        RECT 2912.805 873.205 2914.015 873.955 ;
        RECT 5.520 873.035 6.900 873.205 ;
        RECT 2909.960 873.035 2910.420 873.205 ;
        RECT 2912.720 873.035 2914.100 873.205 ;
        RECT 5.605 872.285 6.815 873.035 ;
        RECT 2912.805 872.285 2914.015 873.035 ;
        RECT 5.605 871.745 6.125 872.285 ;
        RECT 2913.495 871.745 2914.015 872.285 ;
        RECT 5.605 868.515 6.125 869.055 ;
        RECT 2913.495 868.515 2914.015 869.055 ;
        RECT 5.605 867.765 6.815 868.515 ;
        RECT 2910.045 867.765 2910.335 868.490 ;
        RECT 2912.805 867.765 2914.015 868.515 ;
        RECT 5.520 867.595 6.900 867.765 ;
        RECT 2909.960 867.595 2910.420 867.765 ;
        RECT 2912.720 867.595 2914.100 867.765 ;
        RECT 5.605 866.845 6.815 867.595 ;
        RECT 2912.805 866.845 2914.015 867.595 ;
        RECT 5.605 866.305 6.125 866.845 ;
        RECT 2913.495 866.305 2914.015 866.845 ;
        RECT 5.605 863.075 6.125 863.615 ;
        RECT 2913.495 863.075 2914.015 863.615 ;
        RECT 5.605 862.325 6.815 863.075 ;
        RECT 2910.045 862.325 2910.335 863.050 ;
        RECT 2912.805 862.325 2914.015 863.075 ;
        RECT 5.520 862.155 6.900 862.325 ;
        RECT 2909.960 862.155 2910.420 862.325 ;
        RECT 2912.720 862.155 2914.100 862.325 ;
        RECT 5.605 861.405 6.815 862.155 ;
        RECT 2912.805 861.405 2914.015 862.155 ;
        RECT 5.605 860.865 6.125 861.405 ;
        RECT 2913.495 860.865 2914.015 861.405 ;
        RECT 5.605 857.635 6.125 858.175 ;
        RECT 2913.495 857.635 2914.015 858.175 ;
        RECT 5.605 856.885 6.815 857.635 ;
        RECT 2910.045 856.885 2910.335 857.610 ;
        RECT 2912.805 856.885 2914.015 857.635 ;
        RECT 5.520 856.715 6.900 856.885 ;
        RECT 2909.960 856.715 2910.420 856.885 ;
        RECT 2912.720 856.715 2914.100 856.885 ;
        RECT 5.605 855.965 6.815 856.715 ;
        RECT 2912.805 855.965 2914.015 856.715 ;
        RECT 5.605 855.425 6.125 855.965 ;
        RECT 2913.495 855.425 2914.015 855.965 ;
        RECT 5.605 852.195 6.125 852.735 ;
        RECT 2913.495 852.195 2914.015 852.735 ;
        RECT 5.605 851.445 6.815 852.195 ;
        RECT 2910.045 851.445 2910.335 852.170 ;
        RECT 2912.805 851.445 2914.015 852.195 ;
        RECT 5.520 851.275 6.900 851.445 ;
        RECT 2909.960 851.275 2910.420 851.445 ;
        RECT 2912.720 851.275 2914.100 851.445 ;
        RECT 5.605 850.525 6.815 851.275 ;
        RECT 2912.805 850.525 2914.015 851.275 ;
        RECT 5.605 849.985 6.125 850.525 ;
        RECT 2913.495 849.985 2914.015 850.525 ;
        RECT 5.605 846.755 6.125 847.295 ;
        RECT 2913.495 846.755 2914.015 847.295 ;
        RECT 5.605 846.005 6.815 846.755 ;
        RECT 2910.045 846.005 2910.335 846.730 ;
        RECT 2912.805 846.005 2914.015 846.755 ;
        RECT 5.520 845.835 6.900 846.005 ;
        RECT 2909.960 845.835 2910.420 846.005 ;
        RECT 2912.720 845.835 2914.100 846.005 ;
        RECT 5.605 845.085 6.815 845.835 ;
        RECT 2912.805 845.085 2914.015 845.835 ;
        RECT 5.605 844.545 6.125 845.085 ;
        RECT 2913.495 844.545 2914.015 845.085 ;
        RECT 5.605 841.315 6.125 841.855 ;
        RECT 2913.495 841.315 2914.015 841.855 ;
        RECT 5.605 840.565 6.815 841.315 ;
        RECT 2910.045 840.565 2910.335 841.290 ;
        RECT 2912.805 840.565 2914.015 841.315 ;
        RECT 5.520 840.395 6.900 840.565 ;
        RECT 2909.960 840.395 2910.420 840.565 ;
        RECT 2912.720 840.395 2914.100 840.565 ;
        RECT 5.605 839.645 6.815 840.395 ;
        RECT 2912.805 839.645 2914.015 840.395 ;
        RECT 5.605 839.105 6.125 839.645 ;
        RECT 2913.495 839.105 2914.015 839.645 ;
        RECT 5.605 835.875 6.125 836.415 ;
        RECT 2913.495 835.875 2914.015 836.415 ;
        RECT 5.605 835.125 6.815 835.875 ;
        RECT 2910.045 835.125 2910.335 835.850 ;
        RECT 2912.805 835.125 2914.015 835.875 ;
        RECT 5.520 834.955 6.900 835.125 ;
        RECT 2909.960 834.955 2910.420 835.125 ;
        RECT 2912.720 834.955 2914.100 835.125 ;
        RECT 5.605 834.205 6.815 834.955 ;
        RECT 2912.805 834.205 2914.015 834.955 ;
        RECT 5.605 833.665 6.125 834.205 ;
        RECT 2913.495 833.665 2914.015 834.205 ;
        RECT 5.605 830.435 6.125 830.975 ;
        RECT 2913.495 830.435 2914.015 830.975 ;
        RECT 5.605 829.685 6.815 830.435 ;
        RECT 2910.045 829.685 2910.335 830.410 ;
        RECT 2912.805 829.685 2914.015 830.435 ;
        RECT 5.520 829.515 6.900 829.685 ;
        RECT 2909.960 829.515 2910.420 829.685 ;
        RECT 2912.720 829.515 2914.100 829.685 ;
        RECT 5.605 828.765 6.815 829.515 ;
        RECT 2912.805 828.765 2914.015 829.515 ;
        RECT 5.605 828.225 6.125 828.765 ;
        RECT 2913.495 828.225 2914.015 828.765 ;
        RECT 5.605 824.995 6.125 825.535 ;
        RECT 2913.495 824.995 2914.015 825.535 ;
        RECT 5.605 824.245 6.815 824.995 ;
        RECT 2910.045 824.245 2910.335 824.970 ;
        RECT 2912.805 824.245 2914.015 824.995 ;
        RECT 5.520 824.075 6.900 824.245 ;
        RECT 2909.960 824.075 2910.420 824.245 ;
        RECT 2912.720 824.075 2914.100 824.245 ;
        RECT 5.605 823.325 6.815 824.075 ;
        RECT 2912.805 823.325 2914.015 824.075 ;
        RECT 5.605 822.785 6.125 823.325 ;
        RECT 2913.495 822.785 2914.015 823.325 ;
        RECT 5.605 819.555 6.125 820.095 ;
        RECT 2913.495 819.555 2914.015 820.095 ;
        RECT 5.605 818.805 6.815 819.555 ;
        RECT 2910.045 818.805 2910.335 819.530 ;
        RECT 2912.805 818.805 2914.015 819.555 ;
        RECT 5.520 818.635 6.900 818.805 ;
        RECT 2909.960 818.635 2910.420 818.805 ;
        RECT 2912.720 818.635 2914.100 818.805 ;
        RECT 5.605 817.885 6.815 818.635 ;
        RECT 2912.805 817.885 2914.015 818.635 ;
        RECT 5.605 817.345 6.125 817.885 ;
        RECT 2913.495 817.345 2914.015 817.885 ;
        RECT 5.605 814.115 6.125 814.655 ;
        RECT 2913.495 814.115 2914.015 814.655 ;
        RECT 5.605 813.365 6.815 814.115 ;
        RECT 2910.045 813.365 2910.335 814.090 ;
        RECT 2912.805 813.365 2914.015 814.115 ;
        RECT 5.520 813.195 6.900 813.365 ;
        RECT 2909.040 813.195 2910.420 813.365 ;
        RECT 2912.720 813.195 2914.100 813.365 ;
        RECT 5.605 812.445 6.815 813.195 ;
        RECT 2909.815 812.535 2910.155 813.195 ;
        RECT 2912.805 812.445 2914.015 813.195 ;
        RECT 5.605 811.905 6.125 812.445 ;
        RECT 2913.495 811.905 2914.015 812.445 ;
        RECT 5.605 808.675 6.125 809.215 ;
        RECT 2913.495 808.675 2914.015 809.215 ;
        RECT 5.605 807.925 6.815 808.675 ;
        RECT 2910.045 807.925 2910.335 808.650 ;
        RECT 2912.805 807.925 2914.015 808.675 ;
        RECT 5.520 807.755 6.900 807.925 ;
        RECT 2909.960 807.755 2910.420 807.925 ;
        RECT 2912.720 807.755 2914.100 807.925 ;
        RECT 5.605 807.005 6.815 807.755 ;
        RECT 2912.805 807.005 2914.015 807.755 ;
        RECT 5.605 806.465 6.125 807.005 ;
        RECT 2913.495 806.465 2914.015 807.005 ;
        RECT 5.605 803.235 6.125 803.775 ;
        RECT 2913.495 803.235 2914.015 803.775 ;
        RECT 5.605 802.485 6.815 803.235 ;
        RECT 2910.045 802.485 2910.335 803.210 ;
        RECT 2912.805 802.485 2914.015 803.235 ;
        RECT 5.520 802.315 6.900 802.485 ;
        RECT 2909.960 802.315 2910.420 802.485 ;
        RECT 2912.720 802.315 2914.100 802.485 ;
        RECT 5.605 801.565 6.815 802.315 ;
        RECT 2912.805 801.565 2914.015 802.315 ;
        RECT 5.605 801.025 6.125 801.565 ;
        RECT 2913.495 801.025 2914.015 801.565 ;
        RECT 5.605 797.795 6.125 798.335 ;
        RECT 2913.495 797.795 2914.015 798.335 ;
        RECT 5.605 797.045 6.815 797.795 ;
        RECT 2910.045 797.045 2910.335 797.770 ;
        RECT 2912.805 797.045 2914.015 797.795 ;
        RECT 5.520 796.875 6.900 797.045 ;
        RECT 2909.960 796.875 2910.420 797.045 ;
        RECT 2912.720 796.875 2914.100 797.045 ;
        RECT 5.605 796.125 6.815 796.875 ;
        RECT 2912.805 796.125 2914.015 796.875 ;
        RECT 5.605 795.585 6.125 796.125 ;
        RECT 2913.495 795.585 2914.015 796.125 ;
        RECT 5.605 792.355 6.125 792.895 ;
        RECT 2913.495 792.355 2914.015 792.895 ;
        RECT 5.605 791.605 6.815 792.355 ;
        RECT 2910.045 791.605 2910.335 792.330 ;
        RECT 2912.805 791.605 2914.015 792.355 ;
        RECT 5.520 791.435 6.900 791.605 ;
        RECT 2909.960 791.435 2910.420 791.605 ;
        RECT 2912.720 791.435 2914.100 791.605 ;
        RECT 5.605 790.685 6.815 791.435 ;
        RECT 2912.805 790.685 2914.015 791.435 ;
        RECT 5.605 790.145 6.125 790.685 ;
        RECT 2913.495 790.145 2914.015 790.685 ;
        RECT 5.605 786.915 6.125 787.455 ;
        RECT 2913.495 786.915 2914.015 787.455 ;
        RECT 5.605 786.165 6.815 786.915 ;
        RECT 2910.045 786.165 2910.335 786.890 ;
        RECT 2912.805 786.165 2914.015 786.915 ;
        RECT 5.520 785.995 6.900 786.165 ;
        RECT 2909.960 785.995 2910.420 786.165 ;
        RECT 2912.720 785.995 2914.100 786.165 ;
        RECT 5.605 785.245 6.815 785.995 ;
        RECT 2912.805 785.245 2914.015 785.995 ;
        RECT 5.605 784.705 6.125 785.245 ;
        RECT 2913.495 784.705 2914.015 785.245 ;
        RECT 5.605 781.475 6.125 782.015 ;
        RECT 2913.495 781.475 2914.015 782.015 ;
        RECT 5.605 780.725 6.815 781.475 ;
        RECT 2910.045 780.725 2910.335 781.450 ;
        RECT 2912.805 780.725 2914.015 781.475 ;
        RECT 5.520 780.555 6.900 780.725 ;
        RECT 2909.960 780.555 2910.420 780.725 ;
        RECT 2912.720 780.555 2914.100 780.725 ;
        RECT 5.605 779.805 6.815 780.555 ;
        RECT 2912.805 779.805 2914.015 780.555 ;
        RECT 5.605 779.265 6.125 779.805 ;
        RECT 2913.495 779.265 2914.015 779.805 ;
        RECT 5.605 776.035 6.125 776.575 ;
        RECT 2913.495 776.035 2914.015 776.575 ;
        RECT 5.605 775.285 6.815 776.035 ;
        RECT 2910.045 775.285 2910.335 776.010 ;
        RECT 2912.805 775.285 2914.015 776.035 ;
        RECT 5.520 775.115 6.900 775.285 ;
        RECT 2909.960 775.115 2910.420 775.285 ;
        RECT 2912.720 775.115 2914.100 775.285 ;
        RECT 5.605 774.365 6.815 775.115 ;
        RECT 2912.805 774.365 2914.015 775.115 ;
        RECT 5.605 773.825 6.125 774.365 ;
        RECT 2913.495 773.825 2914.015 774.365 ;
        RECT 5.605 770.595 6.125 771.135 ;
        RECT 2913.495 770.595 2914.015 771.135 ;
        RECT 5.605 769.845 6.815 770.595 ;
        RECT 2910.045 769.845 2910.335 770.570 ;
        RECT 2912.805 769.845 2914.015 770.595 ;
        RECT 5.520 769.675 6.900 769.845 ;
        RECT 2909.960 769.675 2910.420 769.845 ;
        RECT 2912.720 769.675 2914.100 769.845 ;
        RECT 5.605 768.925 6.815 769.675 ;
        RECT 2912.805 768.925 2914.015 769.675 ;
        RECT 5.605 768.385 6.125 768.925 ;
        RECT 2913.495 768.385 2914.015 768.925 ;
        RECT 5.605 765.155 6.125 765.695 ;
        RECT 2913.495 765.155 2914.015 765.695 ;
        RECT 5.605 764.405 6.815 765.155 ;
        RECT 2910.045 764.405 2910.335 765.130 ;
        RECT 2912.805 764.405 2914.015 765.155 ;
        RECT 5.520 764.235 6.900 764.405 ;
        RECT 2909.960 764.235 2910.420 764.405 ;
        RECT 2912.720 764.235 2914.100 764.405 ;
        RECT 5.605 763.485 6.815 764.235 ;
        RECT 2912.805 763.485 2914.015 764.235 ;
        RECT 5.605 762.945 6.125 763.485 ;
        RECT 2913.495 762.945 2914.015 763.485 ;
        RECT 5.605 759.715 6.125 760.255 ;
        RECT 2913.495 759.715 2914.015 760.255 ;
        RECT 5.605 758.965 6.815 759.715 ;
        RECT 2910.045 758.965 2910.335 759.690 ;
        RECT 2912.805 758.965 2914.015 759.715 ;
        RECT 5.520 758.795 6.900 758.965 ;
        RECT 2909.960 758.795 2910.420 758.965 ;
        RECT 2912.720 758.795 2914.100 758.965 ;
        RECT 5.605 758.045 6.815 758.795 ;
        RECT 2912.805 758.045 2914.015 758.795 ;
        RECT 5.605 757.505 6.125 758.045 ;
        RECT 2913.495 757.505 2914.015 758.045 ;
        RECT 5.605 754.275 6.125 754.815 ;
        RECT 2913.495 754.275 2914.015 754.815 ;
        RECT 5.605 753.525 6.815 754.275 ;
        RECT 2910.045 753.525 2910.335 754.250 ;
        RECT 2912.805 753.525 2914.015 754.275 ;
        RECT 5.520 753.355 6.900 753.525 ;
        RECT 2909.960 753.355 2910.420 753.525 ;
        RECT 2912.720 753.355 2914.100 753.525 ;
        RECT 5.605 752.605 6.815 753.355 ;
        RECT 2912.805 752.605 2914.015 753.355 ;
        RECT 5.605 752.065 6.125 752.605 ;
        RECT 2913.495 752.065 2914.015 752.605 ;
        RECT 5.605 748.835 6.125 749.375 ;
        RECT 2913.495 748.835 2914.015 749.375 ;
        RECT 5.605 748.085 6.815 748.835 ;
        RECT 2910.045 748.085 2910.335 748.810 ;
        RECT 2912.805 748.085 2914.015 748.835 ;
        RECT 5.520 747.915 6.900 748.085 ;
        RECT 2909.960 747.915 2910.420 748.085 ;
        RECT 2912.720 747.915 2914.100 748.085 ;
        RECT 5.605 747.165 6.815 747.915 ;
        RECT 2912.805 747.165 2914.015 747.915 ;
        RECT 5.605 746.625 6.125 747.165 ;
        RECT 2913.495 746.625 2914.015 747.165 ;
        RECT 5.605 743.395 6.125 743.935 ;
        RECT 2913.495 743.395 2914.015 743.935 ;
        RECT 5.605 742.645 6.815 743.395 ;
        RECT 2910.045 742.645 2910.335 743.370 ;
        RECT 2912.805 742.645 2914.015 743.395 ;
        RECT 5.520 742.475 6.900 742.645 ;
        RECT 2909.960 742.475 2910.420 742.645 ;
        RECT 2912.720 742.475 2914.100 742.645 ;
        RECT 5.605 741.725 6.815 742.475 ;
        RECT 2912.805 741.725 2914.015 742.475 ;
        RECT 5.605 741.185 6.125 741.725 ;
        RECT 2913.495 741.185 2914.015 741.725 ;
        RECT 5.605 737.955 6.125 738.495 ;
        RECT 2913.495 737.955 2914.015 738.495 ;
        RECT 5.605 737.205 6.815 737.955 ;
        RECT 2910.045 737.205 2910.335 737.930 ;
        RECT 2912.805 737.205 2914.015 737.955 ;
        RECT 5.520 737.035 6.900 737.205 ;
        RECT 2909.040 737.035 2910.420 737.205 ;
        RECT 2912.720 737.035 2914.100 737.205 ;
        RECT 5.605 736.285 6.815 737.035 ;
        RECT 2909.815 736.375 2910.155 737.035 ;
        RECT 2912.805 736.285 2914.015 737.035 ;
        RECT 5.605 735.745 6.125 736.285 ;
        RECT 2913.495 735.745 2914.015 736.285 ;
        RECT 5.605 732.515 6.125 733.055 ;
        RECT 2913.495 732.515 2914.015 733.055 ;
        RECT 5.605 731.765 6.815 732.515 ;
        RECT 2910.045 731.765 2910.335 732.490 ;
        RECT 2912.805 731.765 2914.015 732.515 ;
        RECT 5.520 731.595 6.900 731.765 ;
        RECT 2909.960 731.595 2910.420 731.765 ;
        RECT 2912.720 731.595 2914.100 731.765 ;
        RECT 5.605 730.845 6.815 731.595 ;
        RECT 2912.805 730.845 2914.015 731.595 ;
        RECT 5.605 730.305 6.125 730.845 ;
        RECT 2913.495 730.305 2914.015 730.845 ;
        RECT 5.605 727.075 6.125 727.615 ;
        RECT 2913.495 727.075 2914.015 727.615 ;
        RECT 5.605 726.325 6.815 727.075 ;
        RECT 2910.045 726.325 2910.335 727.050 ;
        RECT 2912.805 726.325 2914.015 727.075 ;
        RECT 5.520 726.155 6.900 726.325 ;
        RECT 2909.960 726.155 2910.420 726.325 ;
        RECT 2912.720 726.155 2914.100 726.325 ;
        RECT 5.605 725.405 6.815 726.155 ;
        RECT 2912.805 725.405 2914.015 726.155 ;
        RECT 5.605 724.865 6.125 725.405 ;
        RECT 2913.495 724.865 2914.015 725.405 ;
        RECT 5.605 721.635 6.125 722.175 ;
        RECT 2913.495 721.635 2914.015 722.175 ;
        RECT 5.605 720.885 6.815 721.635 ;
        RECT 9.515 720.885 9.855 721.545 ;
        RECT 2910.045 720.885 2910.335 721.610 ;
        RECT 2912.805 720.885 2914.015 721.635 ;
        RECT 5.520 720.715 6.900 720.885 ;
        RECT 8.740 720.715 10.120 720.885 ;
        RECT 2909.960 720.715 2910.420 720.885 ;
        RECT 2912.720 720.715 2914.100 720.885 ;
        RECT 5.605 719.965 6.815 720.715 ;
        RECT 2912.805 719.965 2914.015 720.715 ;
        RECT 5.605 719.425 6.125 719.965 ;
        RECT 2913.495 719.425 2914.015 719.965 ;
        RECT 5.605 716.195 6.125 716.735 ;
        RECT 2913.495 716.195 2914.015 716.735 ;
        RECT 5.605 715.445 6.815 716.195 ;
        RECT 2910.045 715.445 2910.335 716.170 ;
        RECT 2912.805 715.445 2914.015 716.195 ;
        RECT 5.520 715.275 6.900 715.445 ;
        RECT 2909.960 715.275 2910.420 715.445 ;
        RECT 2912.720 715.275 2914.100 715.445 ;
        RECT 5.605 714.525 6.815 715.275 ;
        RECT 2912.805 714.525 2914.015 715.275 ;
        RECT 5.605 713.985 6.125 714.525 ;
        RECT 2913.495 713.985 2914.015 714.525 ;
        RECT 5.605 710.755 6.125 711.295 ;
        RECT 2913.495 710.755 2914.015 711.295 ;
        RECT 5.605 710.005 6.815 710.755 ;
        RECT 2910.045 710.005 2910.335 710.730 ;
        RECT 2912.805 710.005 2914.015 710.755 ;
        RECT 5.520 709.835 6.900 710.005 ;
        RECT 2909.960 709.835 2910.420 710.005 ;
        RECT 2912.720 709.835 2914.100 710.005 ;
        RECT 5.605 709.085 6.815 709.835 ;
        RECT 2912.805 709.085 2914.015 709.835 ;
        RECT 5.605 708.545 6.125 709.085 ;
        RECT 2913.495 708.545 2914.015 709.085 ;
        RECT 5.605 705.315 6.125 705.855 ;
        RECT 2913.495 705.315 2914.015 705.855 ;
        RECT 5.605 704.565 6.815 705.315 ;
        RECT 2910.045 704.565 2910.335 705.290 ;
        RECT 2912.805 704.565 2914.015 705.315 ;
        RECT 5.520 704.395 6.900 704.565 ;
        RECT 2909.960 704.395 2910.420 704.565 ;
        RECT 2912.720 704.395 2914.100 704.565 ;
        RECT 5.605 703.645 6.815 704.395 ;
        RECT 2912.805 703.645 2914.015 704.395 ;
        RECT 5.605 703.105 6.125 703.645 ;
        RECT 2913.495 703.105 2914.015 703.645 ;
        RECT 5.605 699.875 6.125 700.415 ;
        RECT 2913.495 699.875 2914.015 700.415 ;
        RECT 5.605 699.125 6.815 699.875 ;
        RECT 2910.045 699.125 2910.335 699.850 ;
        RECT 2912.805 699.125 2914.015 699.875 ;
        RECT 5.520 698.955 6.900 699.125 ;
        RECT 2909.960 698.955 2910.420 699.125 ;
        RECT 2912.720 698.955 2914.100 699.125 ;
        RECT 5.605 698.205 6.815 698.955 ;
        RECT 2912.805 698.205 2914.015 698.955 ;
        RECT 5.605 697.665 6.125 698.205 ;
        RECT 2913.495 697.665 2914.015 698.205 ;
        RECT 5.605 694.435 6.125 694.975 ;
        RECT 2913.495 694.435 2914.015 694.975 ;
        RECT 5.605 693.685 6.815 694.435 ;
        RECT 2910.045 693.685 2910.335 694.410 ;
        RECT 2912.805 693.685 2914.015 694.435 ;
        RECT 5.520 693.515 6.900 693.685 ;
        RECT 2909.960 693.515 2910.420 693.685 ;
        RECT 2912.720 693.515 2914.100 693.685 ;
        RECT 5.605 692.765 6.815 693.515 ;
        RECT 2912.805 692.765 2914.015 693.515 ;
        RECT 5.605 692.225 6.125 692.765 ;
        RECT 2913.495 692.225 2914.015 692.765 ;
        RECT 5.605 688.995 6.125 689.535 ;
        RECT 2913.495 688.995 2914.015 689.535 ;
        RECT 5.605 688.245 6.815 688.995 ;
        RECT 2910.045 688.245 2910.335 688.970 ;
        RECT 2912.805 688.245 2914.015 688.995 ;
        RECT 5.520 688.075 6.900 688.245 ;
        RECT 2909.960 688.075 2910.420 688.245 ;
        RECT 2912.720 688.075 2914.100 688.245 ;
        RECT 5.605 687.325 6.815 688.075 ;
        RECT 2912.805 687.325 2914.015 688.075 ;
        RECT 5.605 686.785 6.125 687.325 ;
        RECT 2913.495 686.785 2914.015 687.325 ;
        RECT 5.605 683.555 6.125 684.095 ;
        RECT 2913.495 683.555 2914.015 684.095 ;
        RECT 5.605 682.805 6.815 683.555 ;
        RECT 2910.045 682.805 2910.335 683.530 ;
        RECT 2912.805 682.805 2914.015 683.555 ;
        RECT 5.520 682.635 6.900 682.805 ;
        RECT 2909.960 682.635 2910.420 682.805 ;
        RECT 2912.720 682.635 2914.100 682.805 ;
        RECT 5.605 681.885 6.815 682.635 ;
        RECT 2912.805 681.885 2914.015 682.635 ;
        RECT 5.605 681.345 6.125 681.885 ;
        RECT 2913.495 681.345 2914.015 681.885 ;
        RECT 5.605 678.115 6.125 678.655 ;
        RECT 2913.495 678.115 2914.015 678.655 ;
        RECT 5.605 677.365 6.815 678.115 ;
        RECT 2910.045 677.365 2910.335 678.090 ;
        RECT 2912.805 677.365 2914.015 678.115 ;
        RECT 5.520 677.195 6.900 677.365 ;
        RECT 2909.960 677.195 2910.420 677.365 ;
        RECT 2912.720 677.195 2914.100 677.365 ;
        RECT 5.605 676.445 6.815 677.195 ;
        RECT 2912.805 676.445 2914.015 677.195 ;
        RECT 5.605 675.905 6.125 676.445 ;
        RECT 2913.495 675.905 2914.015 676.445 ;
        RECT 5.605 672.675 6.125 673.215 ;
        RECT 2913.495 672.675 2914.015 673.215 ;
        RECT 5.605 671.925 6.815 672.675 ;
        RECT 2910.045 671.925 2910.335 672.650 ;
        RECT 2912.805 671.925 2914.015 672.675 ;
        RECT 5.520 671.755 6.900 671.925 ;
        RECT 2909.960 671.755 2910.420 671.925 ;
        RECT 2912.720 671.755 2914.100 671.925 ;
        RECT 5.605 671.005 6.815 671.755 ;
        RECT 2912.805 671.005 2914.015 671.755 ;
        RECT 5.605 670.465 6.125 671.005 ;
        RECT 2913.495 670.465 2914.015 671.005 ;
        RECT 5.605 667.235 6.125 667.775 ;
        RECT 2913.495 667.235 2914.015 667.775 ;
        RECT 5.605 666.485 6.815 667.235 ;
        RECT 2910.045 666.485 2910.335 667.210 ;
        RECT 2912.805 666.485 2914.015 667.235 ;
        RECT 5.520 666.315 6.900 666.485 ;
        RECT 2909.960 666.315 2910.420 666.485 ;
        RECT 2912.720 666.315 2914.100 666.485 ;
        RECT 5.605 665.565 6.815 666.315 ;
        RECT 2912.805 665.565 2914.015 666.315 ;
        RECT 5.605 665.025 6.125 665.565 ;
        RECT 2913.495 665.025 2914.015 665.565 ;
        RECT 5.605 661.795 6.125 662.335 ;
        RECT 2913.495 661.795 2914.015 662.335 ;
        RECT 5.605 661.045 6.815 661.795 ;
        RECT 2910.045 661.045 2910.335 661.770 ;
        RECT 2912.805 661.045 2914.015 661.795 ;
        RECT 5.520 660.875 6.900 661.045 ;
        RECT 2909.960 660.875 2910.420 661.045 ;
        RECT 2912.720 660.875 2914.100 661.045 ;
        RECT 5.605 660.125 6.815 660.875 ;
        RECT 2912.805 660.125 2914.015 660.875 ;
        RECT 5.605 659.585 6.125 660.125 ;
        RECT 2913.495 659.585 2914.015 660.125 ;
        RECT 5.605 656.355 6.125 656.895 ;
        RECT 2913.495 656.355 2914.015 656.895 ;
        RECT 5.605 655.605 6.815 656.355 ;
        RECT 2910.045 655.605 2910.335 656.330 ;
        RECT 2912.805 655.605 2914.015 656.355 ;
        RECT 5.520 655.435 6.900 655.605 ;
        RECT 2909.960 655.435 2910.420 655.605 ;
        RECT 2912.720 655.435 2914.100 655.605 ;
        RECT 5.605 654.685 6.815 655.435 ;
        RECT 2912.805 654.685 2914.015 655.435 ;
        RECT 5.605 654.145 6.125 654.685 ;
        RECT 2913.495 654.145 2914.015 654.685 ;
        RECT 5.605 650.915 6.125 651.455 ;
        RECT 2913.495 650.915 2914.015 651.455 ;
        RECT 5.605 650.165 6.815 650.915 ;
        RECT 2910.045 650.165 2910.335 650.890 ;
        RECT 2912.805 650.165 2914.015 650.915 ;
        RECT 5.520 649.995 6.900 650.165 ;
        RECT 2909.960 649.995 2910.420 650.165 ;
        RECT 2912.720 649.995 2914.100 650.165 ;
        RECT 5.605 649.245 6.815 649.995 ;
        RECT 2912.805 649.245 2914.015 649.995 ;
        RECT 5.605 648.705 6.125 649.245 ;
        RECT 2913.495 648.705 2914.015 649.245 ;
        RECT 5.605 645.475 6.125 646.015 ;
        RECT 2913.495 645.475 2914.015 646.015 ;
        RECT 5.605 644.725 6.815 645.475 ;
        RECT 2910.045 644.725 2910.335 645.450 ;
        RECT 2912.805 644.725 2914.015 645.475 ;
        RECT 5.520 644.555 6.900 644.725 ;
        RECT 2909.960 644.555 2910.420 644.725 ;
        RECT 2912.720 644.555 2914.100 644.725 ;
        RECT 5.605 643.805 6.815 644.555 ;
        RECT 2912.805 643.805 2914.015 644.555 ;
        RECT 5.605 643.265 6.125 643.805 ;
        RECT 2913.495 643.265 2914.015 643.805 ;
        RECT 5.605 640.035 6.125 640.575 ;
        RECT 2913.495 640.035 2914.015 640.575 ;
        RECT 5.605 639.285 6.815 640.035 ;
        RECT 2910.045 639.285 2910.335 640.010 ;
        RECT 2912.805 639.285 2914.015 640.035 ;
        RECT 5.520 639.115 6.900 639.285 ;
        RECT 2909.960 639.115 2910.420 639.285 ;
        RECT 2912.720 639.115 2914.100 639.285 ;
        RECT 5.605 638.365 6.815 639.115 ;
        RECT 2912.805 638.365 2914.015 639.115 ;
        RECT 5.605 637.825 6.125 638.365 ;
        RECT 2913.495 637.825 2914.015 638.365 ;
        RECT 5.605 634.595 6.125 635.135 ;
        RECT 2913.495 634.595 2914.015 635.135 ;
        RECT 5.605 633.845 6.815 634.595 ;
        RECT 2910.045 633.845 2910.335 634.570 ;
        RECT 2912.805 633.845 2914.015 634.595 ;
        RECT 5.520 633.675 6.900 633.845 ;
        RECT 2909.960 633.675 2910.420 633.845 ;
        RECT 2912.720 633.675 2914.100 633.845 ;
        RECT 5.605 632.925 6.815 633.675 ;
        RECT 2912.805 632.925 2914.015 633.675 ;
        RECT 5.605 632.385 6.125 632.925 ;
        RECT 2913.495 632.385 2914.015 632.925 ;
        RECT 5.605 629.155 6.125 629.695 ;
        RECT 2913.495 629.155 2914.015 629.695 ;
        RECT 5.605 628.405 6.815 629.155 ;
        RECT 9.515 628.405 9.855 629.065 ;
        RECT 2910.045 628.405 2910.335 629.130 ;
        RECT 2912.805 628.405 2914.015 629.155 ;
        RECT 5.520 628.235 6.900 628.405 ;
        RECT 8.740 628.235 10.120 628.405 ;
        RECT 2909.960 628.235 2910.420 628.405 ;
        RECT 2912.720 628.235 2914.100 628.405 ;
        RECT 5.605 627.485 6.815 628.235 ;
        RECT 2912.805 627.485 2914.015 628.235 ;
        RECT 5.605 626.945 6.125 627.485 ;
        RECT 2913.495 626.945 2914.015 627.485 ;
        RECT 5.605 623.715 6.125 624.255 ;
        RECT 2913.495 623.715 2914.015 624.255 ;
        RECT 5.605 622.965 6.815 623.715 ;
        RECT 2910.045 622.965 2910.335 623.690 ;
        RECT 2912.805 622.965 2914.015 623.715 ;
        RECT 5.520 622.795 6.900 622.965 ;
        RECT 2909.960 622.795 2910.420 622.965 ;
        RECT 2912.720 622.795 2914.100 622.965 ;
        RECT 5.605 622.045 6.815 622.795 ;
        RECT 2912.805 622.045 2914.015 622.795 ;
        RECT 5.605 621.505 6.125 622.045 ;
        RECT 2913.495 621.505 2914.015 622.045 ;
        RECT 5.605 618.275 6.125 618.815 ;
        RECT 2913.495 618.275 2914.015 618.815 ;
        RECT 5.605 617.525 6.815 618.275 ;
        RECT 2910.045 617.525 2910.335 618.250 ;
        RECT 2912.805 617.525 2914.015 618.275 ;
        RECT 5.520 617.355 6.900 617.525 ;
        RECT 2909.960 617.355 2910.420 617.525 ;
        RECT 2912.720 617.355 2914.100 617.525 ;
        RECT 5.605 616.605 6.815 617.355 ;
        RECT 2912.805 616.605 2914.015 617.355 ;
        RECT 5.605 616.065 6.125 616.605 ;
        RECT 2913.495 616.065 2914.015 616.605 ;
        RECT 5.605 612.835 6.125 613.375 ;
        RECT 2913.495 612.835 2914.015 613.375 ;
        RECT 5.605 612.085 6.815 612.835 ;
        RECT 2910.045 612.085 2910.335 612.810 ;
        RECT 2912.805 612.085 2914.015 612.835 ;
        RECT 5.520 611.915 6.900 612.085 ;
        RECT 2909.960 611.915 2910.420 612.085 ;
        RECT 2912.720 611.915 2914.100 612.085 ;
        RECT 5.605 611.165 6.815 611.915 ;
        RECT 2912.805 611.165 2914.015 611.915 ;
        RECT 5.605 610.625 6.125 611.165 ;
        RECT 2913.495 610.625 2914.015 611.165 ;
        RECT 5.605 607.395 6.125 607.935 ;
        RECT 2913.495 607.395 2914.015 607.935 ;
        RECT 5.605 606.645 6.815 607.395 ;
        RECT 2910.045 606.645 2910.335 607.370 ;
        RECT 2912.805 606.645 2914.015 607.395 ;
        RECT 5.520 606.475 6.900 606.645 ;
        RECT 2909.960 606.475 2910.420 606.645 ;
        RECT 2912.720 606.475 2914.100 606.645 ;
        RECT 5.605 605.725 6.815 606.475 ;
        RECT 2912.805 605.725 2914.015 606.475 ;
        RECT 5.605 605.185 6.125 605.725 ;
        RECT 2913.495 605.185 2914.015 605.725 ;
        RECT 5.605 601.955 6.125 602.495 ;
        RECT 2913.495 601.955 2914.015 602.495 ;
        RECT 5.605 601.205 6.815 601.955 ;
        RECT 9.515 601.205 9.855 601.865 ;
        RECT 2910.045 601.205 2910.335 601.930 ;
        RECT 2912.805 601.205 2914.015 601.955 ;
        RECT 5.520 601.035 6.900 601.205 ;
        RECT 8.740 601.035 10.120 601.205 ;
        RECT 2909.960 601.035 2910.420 601.205 ;
        RECT 2912.720 601.035 2914.100 601.205 ;
        RECT 5.605 600.285 6.815 601.035 ;
        RECT 2912.805 600.285 2914.015 601.035 ;
        RECT 5.605 599.745 6.125 600.285 ;
        RECT 2913.495 599.745 2914.015 600.285 ;
        RECT 5.605 596.515 6.125 597.055 ;
        RECT 2913.495 596.515 2914.015 597.055 ;
        RECT 5.605 595.765 6.815 596.515 ;
        RECT 2910.045 595.765 2910.335 596.490 ;
        RECT 2912.805 595.765 2914.015 596.515 ;
        RECT 5.520 595.595 6.900 595.765 ;
        RECT 2909.960 595.595 2910.420 595.765 ;
        RECT 2912.720 595.595 2914.100 595.765 ;
        RECT 5.605 594.845 6.815 595.595 ;
        RECT 2912.805 594.845 2914.015 595.595 ;
        RECT 5.605 594.305 6.125 594.845 ;
        RECT 2913.495 594.305 2914.015 594.845 ;
        RECT 5.605 591.075 6.125 591.615 ;
        RECT 2913.495 591.075 2914.015 591.615 ;
        RECT 5.605 590.325 6.815 591.075 ;
        RECT 2910.045 590.325 2910.335 591.050 ;
        RECT 2912.805 590.325 2914.015 591.075 ;
        RECT 5.520 590.155 6.900 590.325 ;
        RECT 2909.960 590.155 2910.420 590.325 ;
        RECT 2912.720 590.155 2914.100 590.325 ;
        RECT 5.605 589.405 6.815 590.155 ;
        RECT 2912.805 589.405 2914.015 590.155 ;
        RECT 5.605 588.865 6.125 589.405 ;
        RECT 2913.495 588.865 2914.015 589.405 ;
        RECT 5.605 585.635 6.125 586.175 ;
        RECT 2913.495 585.635 2914.015 586.175 ;
        RECT 5.605 584.885 6.815 585.635 ;
        RECT 2910.045 584.885 2910.335 585.610 ;
        RECT 2912.805 584.885 2914.015 585.635 ;
        RECT 5.520 584.715 6.900 584.885 ;
        RECT 2909.960 584.715 2910.420 584.885 ;
        RECT 2912.720 584.715 2914.100 584.885 ;
        RECT 5.605 583.965 6.815 584.715 ;
        RECT 2912.805 583.965 2914.015 584.715 ;
        RECT 5.605 583.425 6.125 583.965 ;
        RECT 2913.495 583.425 2914.015 583.965 ;
        RECT 5.605 580.195 6.125 580.735 ;
        RECT 2913.495 580.195 2914.015 580.735 ;
        RECT 5.605 579.445 6.815 580.195 ;
        RECT 2910.045 579.445 2910.335 580.170 ;
        RECT 2912.805 579.445 2914.015 580.195 ;
        RECT 5.520 579.275 6.900 579.445 ;
        RECT 2909.960 579.275 2910.420 579.445 ;
        RECT 2912.720 579.275 2914.100 579.445 ;
        RECT 5.605 578.525 6.815 579.275 ;
        RECT 2912.805 578.525 2914.015 579.275 ;
        RECT 5.605 577.985 6.125 578.525 ;
        RECT 2913.495 577.985 2914.015 578.525 ;
        RECT 5.605 574.755 6.125 575.295 ;
        RECT 2913.495 574.755 2914.015 575.295 ;
        RECT 5.605 574.005 6.815 574.755 ;
        RECT 2910.045 574.005 2910.335 574.730 ;
        RECT 2912.805 574.005 2914.015 574.755 ;
        RECT 5.520 573.835 6.900 574.005 ;
        RECT 2909.960 573.835 2910.420 574.005 ;
        RECT 2912.720 573.835 2914.100 574.005 ;
        RECT 5.605 573.085 6.815 573.835 ;
        RECT 2912.805 573.085 2914.015 573.835 ;
        RECT 5.605 572.545 6.125 573.085 ;
        RECT 2913.495 572.545 2914.015 573.085 ;
        RECT 5.605 569.315 6.125 569.855 ;
        RECT 2913.495 569.315 2914.015 569.855 ;
        RECT 5.605 568.565 6.815 569.315 ;
        RECT 2910.045 568.565 2910.335 569.290 ;
        RECT 2912.805 568.565 2914.015 569.315 ;
        RECT 5.520 568.395 6.900 568.565 ;
        RECT 2909.960 568.395 2910.420 568.565 ;
        RECT 2912.720 568.395 2914.100 568.565 ;
        RECT 5.605 567.645 6.815 568.395 ;
        RECT 2912.805 567.645 2914.015 568.395 ;
        RECT 5.605 567.105 6.125 567.645 ;
        RECT 2913.495 567.105 2914.015 567.645 ;
        RECT 5.605 563.875 6.125 564.415 ;
        RECT 2913.495 563.875 2914.015 564.415 ;
        RECT 5.605 563.125 6.815 563.875 ;
        RECT 2910.045 563.125 2910.335 563.850 ;
        RECT 2912.805 563.125 2914.015 563.875 ;
        RECT 5.520 562.955 6.900 563.125 ;
        RECT 2909.960 562.955 2910.420 563.125 ;
        RECT 2912.720 562.955 2914.100 563.125 ;
        RECT 5.605 562.205 6.815 562.955 ;
        RECT 2912.805 562.205 2914.015 562.955 ;
        RECT 5.605 561.665 6.125 562.205 ;
        RECT 2913.495 561.665 2914.015 562.205 ;
        RECT 5.605 558.435 6.125 558.975 ;
        RECT 2913.495 558.435 2914.015 558.975 ;
        RECT 5.605 557.685 6.815 558.435 ;
        RECT 2910.045 557.685 2910.335 558.410 ;
        RECT 2912.805 557.685 2914.015 558.435 ;
        RECT 5.520 557.515 6.900 557.685 ;
        RECT 2909.960 557.515 2910.420 557.685 ;
        RECT 2912.720 557.515 2914.100 557.685 ;
        RECT 5.605 556.765 6.815 557.515 ;
        RECT 2912.805 556.765 2914.015 557.515 ;
        RECT 5.605 556.225 6.125 556.765 ;
        RECT 2913.495 556.225 2914.015 556.765 ;
        RECT 5.605 552.995 6.125 553.535 ;
        RECT 2913.495 552.995 2914.015 553.535 ;
        RECT 5.605 552.245 6.815 552.995 ;
        RECT 2910.045 552.245 2910.335 552.970 ;
        RECT 2912.805 552.245 2914.015 552.995 ;
        RECT 5.520 552.075 6.900 552.245 ;
        RECT 2909.960 552.075 2910.420 552.245 ;
        RECT 2912.720 552.075 2914.100 552.245 ;
        RECT 5.605 551.325 6.815 552.075 ;
        RECT 2912.805 551.325 2914.015 552.075 ;
        RECT 5.605 550.785 6.125 551.325 ;
        RECT 2913.495 550.785 2914.015 551.325 ;
        RECT 5.605 547.555 6.125 548.095 ;
        RECT 2913.495 547.555 2914.015 548.095 ;
        RECT 5.605 546.805 6.815 547.555 ;
        RECT 2910.045 546.805 2910.335 547.530 ;
        RECT 2912.805 546.805 2914.015 547.555 ;
        RECT 5.520 546.635 6.900 546.805 ;
        RECT 2909.960 546.635 2910.420 546.805 ;
        RECT 2912.720 546.635 2914.100 546.805 ;
        RECT 5.605 545.885 6.815 546.635 ;
        RECT 2912.805 545.885 2914.015 546.635 ;
        RECT 5.605 545.345 6.125 545.885 ;
        RECT 2913.495 545.345 2914.015 545.885 ;
        RECT 5.605 542.115 6.125 542.655 ;
        RECT 2913.495 542.115 2914.015 542.655 ;
        RECT 5.605 541.365 6.815 542.115 ;
        RECT 2910.045 541.365 2910.335 542.090 ;
        RECT 2912.805 541.365 2914.015 542.115 ;
        RECT 5.520 541.195 6.900 541.365 ;
        RECT 2909.960 541.195 2910.420 541.365 ;
        RECT 2912.720 541.195 2914.100 541.365 ;
        RECT 5.605 540.445 6.815 541.195 ;
        RECT 2912.805 540.445 2914.015 541.195 ;
        RECT 5.605 539.905 6.125 540.445 ;
        RECT 2913.495 539.905 2914.015 540.445 ;
        RECT 5.605 536.675 6.125 537.215 ;
        RECT 2913.495 536.675 2914.015 537.215 ;
        RECT 5.605 535.925 6.815 536.675 ;
        RECT 2910.045 535.925 2910.335 536.650 ;
        RECT 2912.805 535.925 2914.015 536.675 ;
        RECT 5.520 535.755 6.900 535.925 ;
        RECT 2909.960 535.755 2910.420 535.925 ;
        RECT 2912.720 535.755 2914.100 535.925 ;
        RECT 5.605 535.005 6.815 535.755 ;
        RECT 2912.805 535.005 2914.015 535.755 ;
        RECT 5.605 534.465 6.125 535.005 ;
        RECT 2913.495 534.465 2914.015 535.005 ;
        RECT 5.605 531.235 6.125 531.775 ;
        RECT 2913.495 531.235 2914.015 531.775 ;
        RECT 5.605 530.485 6.815 531.235 ;
        RECT 2910.045 530.485 2910.335 531.210 ;
        RECT 2912.805 530.485 2914.015 531.235 ;
        RECT 5.520 530.315 6.900 530.485 ;
        RECT 2909.960 530.315 2910.420 530.485 ;
        RECT 2912.720 530.315 2914.100 530.485 ;
        RECT 5.605 529.565 6.815 530.315 ;
        RECT 2912.805 529.565 2914.015 530.315 ;
        RECT 5.605 529.025 6.125 529.565 ;
        RECT 2913.495 529.025 2914.015 529.565 ;
        RECT 5.605 525.795 6.125 526.335 ;
        RECT 2913.495 525.795 2914.015 526.335 ;
        RECT 5.605 525.045 6.815 525.795 ;
        RECT 2910.045 525.045 2910.335 525.770 ;
        RECT 2912.805 525.045 2914.015 525.795 ;
        RECT 5.520 524.875 6.900 525.045 ;
        RECT 2909.960 524.875 2910.420 525.045 ;
        RECT 2912.720 524.875 2914.100 525.045 ;
        RECT 5.605 524.125 6.815 524.875 ;
        RECT 2912.805 524.125 2914.015 524.875 ;
        RECT 5.605 523.585 6.125 524.125 ;
        RECT 2913.495 523.585 2914.015 524.125 ;
        RECT 5.605 520.355 6.125 520.895 ;
        RECT 2913.495 520.355 2914.015 520.895 ;
        RECT 5.605 519.605 6.815 520.355 ;
        RECT 2910.045 519.605 2910.335 520.330 ;
        RECT 2912.805 519.605 2914.015 520.355 ;
        RECT 5.520 519.435 6.900 519.605 ;
        RECT 2909.960 519.435 2910.420 519.605 ;
        RECT 2912.720 519.435 2914.100 519.605 ;
        RECT 5.605 518.685 6.815 519.435 ;
        RECT 2912.805 518.685 2914.015 519.435 ;
        RECT 5.605 518.145 6.125 518.685 ;
        RECT 2913.495 518.145 2914.015 518.685 ;
        RECT 5.605 514.915 6.125 515.455 ;
        RECT 2913.495 514.915 2914.015 515.455 ;
        RECT 5.605 514.165 6.815 514.915 ;
        RECT 2910.045 514.165 2910.335 514.890 ;
        RECT 2912.805 514.165 2914.015 514.915 ;
        RECT 5.520 513.995 6.900 514.165 ;
        RECT 2909.960 513.995 2910.420 514.165 ;
        RECT 2912.720 513.995 2914.100 514.165 ;
        RECT 5.605 513.245 6.815 513.995 ;
        RECT 2912.805 513.245 2914.015 513.995 ;
        RECT 5.605 512.705 6.125 513.245 ;
        RECT 2913.495 512.705 2914.015 513.245 ;
        RECT 5.605 509.475 6.125 510.015 ;
        RECT 2913.495 509.475 2914.015 510.015 ;
        RECT 5.605 508.725 6.815 509.475 ;
        RECT 2910.045 508.725 2910.335 509.450 ;
        RECT 2912.805 508.725 2914.015 509.475 ;
        RECT 5.520 508.555 6.900 508.725 ;
        RECT 2909.960 508.555 2910.420 508.725 ;
        RECT 2912.720 508.555 2914.100 508.725 ;
        RECT 5.605 507.805 6.815 508.555 ;
        RECT 2912.805 507.805 2914.015 508.555 ;
        RECT 5.605 507.265 6.125 507.805 ;
        RECT 2913.495 507.265 2914.015 507.805 ;
        RECT 5.605 504.035 6.125 504.575 ;
        RECT 2913.495 504.035 2914.015 504.575 ;
        RECT 5.605 503.285 6.815 504.035 ;
        RECT 2910.045 503.285 2910.335 504.010 ;
        RECT 2912.805 503.285 2914.015 504.035 ;
        RECT 5.520 503.115 6.900 503.285 ;
        RECT 2909.960 503.115 2910.420 503.285 ;
        RECT 2912.720 503.115 2914.100 503.285 ;
        RECT 5.605 502.365 6.815 503.115 ;
        RECT 2912.805 502.365 2914.015 503.115 ;
        RECT 5.605 501.825 6.125 502.365 ;
        RECT 2913.495 501.825 2914.015 502.365 ;
        RECT 5.605 498.595 6.125 499.135 ;
        RECT 2913.495 498.595 2914.015 499.135 ;
        RECT 5.605 497.845 6.815 498.595 ;
        RECT 2910.045 497.845 2910.335 498.570 ;
        RECT 2912.805 497.845 2914.015 498.595 ;
        RECT 5.520 497.675 6.900 497.845 ;
        RECT 2909.960 497.675 2910.420 497.845 ;
        RECT 2912.720 497.675 2914.100 497.845 ;
        RECT 5.605 496.925 6.815 497.675 ;
        RECT 2912.805 496.925 2914.015 497.675 ;
        RECT 5.605 496.385 6.125 496.925 ;
        RECT 2913.495 496.385 2914.015 496.925 ;
        RECT 5.605 493.155 6.125 493.695 ;
        RECT 2913.495 493.155 2914.015 493.695 ;
        RECT 5.605 492.405 6.815 493.155 ;
        RECT 2910.045 492.405 2910.335 493.130 ;
        RECT 2912.805 492.405 2914.015 493.155 ;
        RECT 5.520 492.235 6.900 492.405 ;
        RECT 2909.960 492.235 2910.420 492.405 ;
        RECT 2912.720 492.235 2914.100 492.405 ;
        RECT 5.605 491.485 6.815 492.235 ;
        RECT 2912.805 491.485 2914.015 492.235 ;
        RECT 5.605 490.945 6.125 491.485 ;
        RECT 2913.495 490.945 2914.015 491.485 ;
        RECT 5.605 487.715 6.125 488.255 ;
        RECT 2913.495 487.715 2914.015 488.255 ;
        RECT 5.605 486.965 6.815 487.715 ;
        RECT 2910.045 486.965 2910.335 487.690 ;
        RECT 2912.805 486.965 2914.015 487.715 ;
        RECT 5.520 486.795 6.900 486.965 ;
        RECT 2909.960 486.795 2910.420 486.965 ;
        RECT 2912.720 486.795 2914.100 486.965 ;
        RECT 5.605 486.045 6.815 486.795 ;
        RECT 2912.805 486.045 2914.015 486.795 ;
        RECT 5.605 485.505 6.125 486.045 ;
        RECT 2913.495 485.505 2914.015 486.045 ;
        RECT 5.605 482.275 6.125 482.815 ;
        RECT 2913.495 482.275 2914.015 482.815 ;
        RECT 5.605 481.525 6.815 482.275 ;
        RECT 2910.045 481.525 2910.335 482.250 ;
        RECT 2912.805 481.525 2914.015 482.275 ;
        RECT 5.520 481.355 6.900 481.525 ;
        RECT 2909.960 481.355 2910.420 481.525 ;
        RECT 2912.720 481.355 2914.100 481.525 ;
        RECT 5.605 480.605 6.815 481.355 ;
        RECT 2912.805 480.605 2914.015 481.355 ;
        RECT 5.605 480.065 6.125 480.605 ;
        RECT 2913.495 480.065 2914.015 480.605 ;
        RECT 5.605 476.835 6.125 477.375 ;
        RECT 2913.495 476.835 2914.015 477.375 ;
        RECT 5.605 476.085 6.815 476.835 ;
        RECT 2910.045 476.085 2910.335 476.810 ;
        RECT 2912.805 476.085 2914.015 476.835 ;
        RECT 5.520 475.915 6.900 476.085 ;
        RECT 2909.960 475.915 2910.420 476.085 ;
        RECT 2912.720 475.915 2914.100 476.085 ;
        RECT 5.605 475.165 6.815 475.915 ;
        RECT 2912.805 475.165 2914.015 475.915 ;
        RECT 5.605 474.625 6.125 475.165 ;
        RECT 2913.495 474.625 2914.015 475.165 ;
        RECT 5.605 471.395 6.125 471.935 ;
        RECT 2913.495 471.395 2914.015 471.935 ;
        RECT 5.605 470.645 6.815 471.395 ;
        RECT 2910.045 470.645 2910.335 471.370 ;
        RECT 2912.805 470.645 2914.015 471.395 ;
        RECT 5.520 470.475 6.900 470.645 ;
        RECT 2909.040 470.475 2910.420 470.645 ;
        RECT 2912.720 470.475 2914.100 470.645 ;
        RECT 5.605 469.725 6.815 470.475 ;
        RECT 2909.815 469.815 2910.155 470.475 ;
        RECT 2912.805 469.725 2914.015 470.475 ;
        RECT 5.605 469.185 6.125 469.725 ;
        RECT 2913.495 469.185 2914.015 469.725 ;
        RECT 5.605 465.955 6.125 466.495 ;
        RECT 2913.495 465.955 2914.015 466.495 ;
        RECT 5.605 465.205 6.815 465.955 ;
        RECT 2910.045 465.205 2910.335 465.930 ;
        RECT 2912.805 465.205 2914.015 465.955 ;
        RECT 5.520 465.035 6.900 465.205 ;
        RECT 2909.960 465.035 2910.420 465.205 ;
        RECT 2912.720 465.035 2914.100 465.205 ;
        RECT 5.605 464.285 6.815 465.035 ;
        RECT 2912.805 464.285 2914.015 465.035 ;
        RECT 5.605 463.745 6.125 464.285 ;
        RECT 2913.495 463.745 2914.015 464.285 ;
        RECT 5.605 460.515 6.125 461.055 ;
        RECT 2913.495 460.515 2914.015 461.055 ;
        RECT 5.605 459.765 6.815 460.515 ;
        RECT 2910.045 459.765 2910.335 460.490 ;
        RECT 2912.805 459.765 2914.015 460.515 ;
        RECT 5.520 459.595 6.900 459.765 ;
        RECT 2909.960 459.595 2910.420 459.765 ;
        RECT 2912.720 459.595 2914.100 459.765 ;
        RECT 5.605 458.845 6.815 459.595 ;
        RECT 2912.805 458.845 2914.015 459.595 ;
        RECT 5.605 458.305 6.125 458.845 ;
        RECT 2913.495 458.305 2914.015 458.845 ;
        RECT 5.605 455.075 6.125 455.615 ;
        RECT 2913.495 455.075 2914.015 455.615 ;
        RECT 5.605 454.325 6.815 455.075 ;
        RECT 2910.045 454.325 2910.335 455.050 ;
        RECT 2912.805 454.325 2914.015 455.075 ;
        RECT 5.520 454.155 6.900 454.325 ;
        RECT 2909.960 454.155 2910.420 454.325 ;
        RECT 2912.720 454.155 2914.100 454.325 ;
        RECT 5.605 453.405 6.815 454.155 ;
        RECT 2912.805 453.405 2914.015 454.155 ;
        RECT 5.605 452.865 6.125 453.405 ;
        RECT 2913.495 452.865 2914.015 453.405 ;
        RECT 5.605 449.635 6.125 450.175 ;
        RECT 2913.495 449.635 2914.015 450.175 ;
        RECT 5.605 448.885 6.815 449.635 ;
        RECT 2910.045 448.885 2910.335 449.610 ;
        RECT 2911.195 448.885 2911.535 449.545 ;
        RECT 2912.805 448.885 2914.015 449.635 ;
        RECT 5.520 448.715 6.900 448.885 ;
        RECT 2909.960 448.715 2911.800 448.885 ;
        RECT 2912.720 448.715 2914.100 448.885 ;
        RECT 5.605 447.965 6.815 448.715 ;
        RECT 2912.805 447.965 2914.015 448.715 ;
        RECT 5.605 447.425 6.125 447.965 ;
        RECT 2913.495 447.425 2914.015 447.965 ;
        RECT 5.605 444.195 6.125 444.735 ;
        RECT 2913.495 444.195 2914.015 444.735 ;
        RECT 5.605 443.445 6.815 444.195 ;
        RECT 2910.045 443.445 2910.335 444.170 ;
        RECT 2912.805 443.445 2914.015 444.195 ;
        RECT 5.520 443.275 6.900 443.445 ;
        RECT 8.740 443.275 10.120 443.445 ;
        RECT 2909.960 443.275 2910.420 443.445 ;
        RECT 2912.720 443.275 2914.100 443.445 ;
        RECT 5.605 442.525 6.815 443.275 ;
        RECT 9.515 442.615 9.855 443.275 ;
        RECT 2912.805 442.525 2914.015 443.275 ;
        RECT 5.605 441.985 6.125 442.525 ;
        RECT 2913.495 441.985 2914.015 442.525 ;
        RECT 5.605 438.755 6.125 439.295 ;
        RECT 2913.495 438.755 2914.015 439.295 ;
        RECT 5.605 438.005 6.815 438.755 ;
        RECT 9.515 438.005 9.855 438.665 ;
        RECT 2910.045 438.005 2910.335 438.730 ;
        RECT 2912.805 438.005 2914.015 438.755 ;
        RECT 5.520 437.835 6.900 438.005 ;
        RECT 8.740 437.835 10.120 438.005 ;
        RECT 2909.960 437.835 2910.420 438.005 ;
        RECT 2912.720 437.835 2914.100 438.005 ;
        RECT 5.605 437.085 6.815 437.835 ;
        RECT 2912.805 437.085 2914.015 437.835 ;
        RECT 5.605 436.545 6.125 437.085 ;
        RECT 2913.495 436.545 2914.015 437.085 ;
        RECT 5.605 433.315 6.125 433.855 ;
        RECT 2913.495 433.315 2914.015 433.855 ;
        RECT 5.605 432.565 6.815 433.315 ;
        RECT 2910.045 432.565 2910.335 433.290 ;
        RECT 2912.805 432.565 2914.015 433.315 ;
        RECT 5.520 432.395 6.900 432.565 ;
        RECT 2909.960 432.395 2910.420 432.565 ;
        RECT 2912.720 432.395 2914.100 432.565 ;
        RECT 5.605 431.645 6.815 432.395 ;
        RECT 2912.805 431.645 2914.015 432.395 ;
        RECT 5.605 431.105 6.125 431.645 ;
        RECT 2913.495 431.105 2914.015 431.645 ;
        RECT 5.605 427.875 6.125 428.415 ;
        RECT 2913.495 427.875 2914.015 428.415 ;
        RECT 5.605 427.125 6.815 427.875 ;
        RECT 2910.045 427.125 2910.335 427.850 ;
        RECT 2912.805 427.125 2914.015 427.875 ;
        RECT 5.520 426.955 6.900 427.125 ;
        RECT 2909.960 426.955 2910.420 427.125 ;
        RECT 2912.720 426.955 2914.100 427.125 ;
        RECT 5.605 426.205 6.815 426.955 ;
        RECT 2912.805 426.205 2914.015 426.955 ;
        RECT 5.605 425.665 6.125 426.205 ;
        RECT 2913.495 425.665 2914.015 426.205 ;
        RECT 5.605 422.435 6.125 422.975 ;
        RECT 2913.495 422.435 2914.015 422.975 ;
        RECT 5.605 421.685 6.815 422.435 ;
        RECT 2910.045 421.685 2910.335 422.410 ;
        RECT 2912.805 421.685 2914.015 422.435 ;
        RECT 5.520 421.515 6.900 421.685 ;
        RECT 2909.960 421.515 2910.420 421.685 ;
        RECT 2912.720 421.515 2914.100 421.685 ;
        RECT 5.605 420.765 6.815 421.515 ;
        RECT 2912.805 420.765 2914.015 421.515 ;
        RECT 5.605 420.225 6.125 420.765 ;
        RECT 2913.495 420.225 2914.015 420.765 ;
        RECT 5.605 416.995 6.125 417.535 ;
        RECT 2913.495 416.995 2914.015 417.535 ;
        RECT 5.605 416.245 6.815 416.995 ;
        RECT 2910.045 416.245 2910.335 416.970 ;
        RECT 2912.805 416.245 2914.015 416.995 ;
        RECT 5.520 416.075 6.900 416.245 ;
        RECT 2909.960 416.075 2910.420 416.245 ;
        RECT 2912.720 416.075 2914.100 416.245 ;
        RECT 5.605 415.325 6.815 416.075 ;
        RECT 2912.805 415.325 2914.015 416.075 ;
        RECT 5.605 414.785 6.125 415.325 ;
        RECT 2913.495 414.785 2914.015 415.325 ;
        RECT 5.605 411.555 6.125 412.095 ;
        RECT 2913.495 411.555 2914.015 412.095 ;
        RECT 5.605 410.805 6.815 411.555 ;
        RECT 2910.045 410.805 2910.335 411.530 ;
        RECT 2912.805 410.805 2914.015 411.555 ;
        RECT 5.520 410.635 6.900 410.805 ;
        RECT 2909.960 410.635 2910.420 410.805 ;
        RECT 2912.720 410.635 2914.100 410.805 ;
        RECT 5.605 409.885 6.815 410.635 ;
        RECT 2912.805 409.885 2914.015 410.635 ;
        RECT 5.605 409.345 6.125 409.885 ;
        RECT 2913.495 409.345 2914.015 409.885 ;
        RECT 5.605 406.115 6.125 406.655 ;
        RECT 2913.495 406.115 2914.015 406.655 ;
        RECT 5.605 405.365 6.815 406.115 ;
        RECT 2910.045 405.365 2910.335 406.090 ;
        RECT 2912.805 405.365 2914.015 406.115 ;
        RECT 5.520 405.195 6.900 405.365 ;
        RECT 2909.960 405.195 2910.420 405.365 ;
        RECT 2912.720 405.195 2914.100 405.365 ;
        RECT 5.605 404.445 6.815 405.195 ;
        RECT 2912.805 404.445 2914.015 405.195 ;
        RECT 5.605 403.905 6.125 404.445 ;
        RECT 2913.495 403.905 2914.015 404.445 ;
        RECT 5.605 400.675 6.125 401.215 ;
        RECT 2913.495 400.675 2914.015 401.215 ;
        RECT 5.605 399.925 6.815 400.675 ;
        RECT 9.515 399.925 9.855 400.585 ;
        RECT 2910.045 399.925 2910.335 400.650 ;
        RECT 2912.805 399.925 2914.015 400.675 ;
        RECT 5.520 399.755 6.900 399.925 ;
        RECT 8.740 399.755 10.120 399.925 ;
        RECT 2909.960 399.755 2910.420 399.925 ;
        RECT 2912.720 399.755 2914.100 399.925 ;
        RECT 5.605 399.005 6.815 399.755 ;
        RECT 2912.805 399.005 2914.015 399.755 ;
        RECT 5.605 398.465 6.125 399.005 ;
        RECT 2913.495 398.465 2914.015 399.005 ;
        RECT 5.605 395.235 6.125 395.775 ;
        RECT 2913.495 395.235 2914.015 395.775 ;
        RECT 5.605 394.485 6.815 395.235 ;
        RECT 2910.045 394.485 2910.335 395.210 ;
        RECT 2912.805 394.485 2914.015 395.235 ;
        RECT 5.520 394.315 6.900 394.485 ;
        RECT 8.740 394.315 10.120 394.485 ;
        RECT 2909.960 394.315 2910.420 394.485 ;
        RECT 2912.720 394.315 2914.100 394.485 ;
        RECT 5.605 393.565 6.815 394.315 ;
        RECT 9.515 393.655 9.855 394.315 ;
        RECT 2912.805 393.565 2914.015 394.315 ;
        RECT 5.605 393.025 6.125 393.565 ;
        RECT 2913.495 393.025 2914.015 393.565 ;
        RECT 5.605 389.795 6.125 390.335 ;
        RECT 2913.495 389.795 2914.015 390.335 ;
        RECT 5.605 389.045 6.815 389.795 ;
        RECT 2910.045 389.045 2910.335 389.770 ;
        RECT 2912.805 389.045 2914.015 389.795 ;
        RECT 5.520 388.875 6.900 389.045 ;
        RECT 2909.960 388.875 2910.420 389.045 ;
        RECT 2912.720 388.875 2914.100 389.045 ;
        RECT 5.605 388.125 6.815 388.875 ;
        RECT 2912.805 388.125 2914.015 388.875 ;
        RECT 5.605 387.585 6.125 388.125 ;
        RECT 2913.495 387.585 2914.015 388.125 ;
        RECT 5.605 384.355 6.125 384.895 ;
        RECT 2913.495 384.355 2914.015 384.895 ;
        RECT 5.605 383.605 6.815 384.355 ;
        RECT 2910.045 383.605 2910.335 384.330 ;
        RECT 2912.805 383.605 2914.015 384.355 ;
        RECT 5.520 383.435 6.900 383.605 ;
        RECT 2909.960 383.435 2910.420 383.605 ;
        RECT 2912.720 383.435 2914.100 383.605 ;
        RECT 5.605 382.685 6.815 383.435 ;
        RECT 2912.805 382.685 2914.015 383.435 ;
        RECT 5.605 382.145 6.125 382.685 ;
        RECT 2913.495 382.145 2914.015 382.685 ;
        RECT 5.605 378.915 6.125 379.455 ;
        RECT 2913.495 378.915 2914.015 379.455 ;
        RECT 5.605 378.165 6.815 378.915 ;
        RECT 2910.045 378.165 2910.335 378.890 ;
        RECT 2912.805 378.165 2914.015 378.915 ;
        RECT 5.520 377.995 6.900 378.165 ;
        RECT 2909.960 377.995 2910.420 378.165 ;
        RECT 2912.720 377.995 2914.100 378.165 ;
        RECT 5.605 377.245 6.815 377.995 ;
        RECT 2912.805 377.245 2914.015 377.995 ;
        RECT 5.605 376.705 6.125 377.245 ;
        RECT 2913.495 376.705 2914.015 377.245 ;
        RECT 5.605 373.475 6.125 374.015 ;
        RECT 2913.495 373.475 2914.015 374.015 ;
        RECT 5.605 372.725 6.815 373.475 ;
        RECT 2910.045 372.725 2910.335 373.450 ;
        RECT 2912.805 372.725 2914.015 373.475 ;
        RECT 5.520 372.555 6.900 372.725 ;
        RECT 2909.960 372.555 2910.420 372.725 ;
        RECT 2912.720 372.555 2914.100 372.725 ;
        RECT 5.605 371.805 6.815 372.555 ;
        RECT 2912.805 371.805 2914.015 372.555 ;
        RECT 5.605 371.265 6.125 371.805 ;
        RECT 2913.495 371.265 2914.015 371.805 ;
        RECT 5.605 368.035 6.125 368.575 ;
        RECT 2913.495 368.035 2914.015 368.575 ;
        RECT 5.605 367.285 6.815 368.035 ;
        RECT 2910.045 367.285 2910.335 368.010 ;
        RECT 2912.805 367.285 2914.015 368.035 ;
        RECT 5.520 367.115 6.900 367.285 ;
        RECT 2909.960 367.115 2910.420 367.285 ;
        RECT 2912.720 367.115 2914.100 367.285 ;
        RECT 5.605 366.365 6.815 367.115 ;
        RECT 2912.805 366.365 2914.015 367.115 ;
        RECT 5.605 365.825 6.125 366.365 ;
        RECT 2913.495 365.825 2914.015 366.365 ;
        RECT 5.605 362.595 6.125 363.135 ;
        RECT 2913.495 362.595 2914.015 363.135 ;
        RECT 5.605 361.845 6.815 362.595 ;
        RECT 2910.045 361.845 2910.335 362.570 ;
        RECT 2912.805 361.845 2914.015 362.595 ;
        RECT 5.520 361.675 6.900 361.845 ;
        RECT 2909.960 361.675 2910.420 361.845 ;
        RECT 2912.720 361.675 2914.100 361.845 ;
        RECT 5.605 360.925 6.815 361.675 ;
        RECT 2912.805 360.925 2914.015 361.675 ;
        RECT 5.605 360.385 6.125 360.925 ;
        RECT 2913.495 360.385 2914.015 360.925 ;
        RECT 5.605 357.155 6.125 357.695 ;
        RECT 2913.495 357.155 2914.015 357.695 ;
        RECT 5.605 356.405 6.815 357.155 ;
        RECT 2910.045 356.405 2910.335 357.130 ;
        RECT 2912.805 356.405 2914.015 357.155 ;
        RECT 5.520 356.235 6.900 356.405 ;
        RECT 2909.960 356.235 2910.420 356.405 ;
        RECT 2912.720 356.235 2914.100 356.405 ;
        RECT 5.605 355.485 6.815 356.235 ;
        RECT 2912.805 355.485 2914.015 356.235 ;
        RECT 5.605 354.945 6.125 355.485 ;
        RECT 2913.495 354.945 2914.015 355.485 ;
        RECT 5.605 351.715 6.125 352.255 ;
        RECT 2913.495 351.715 2914.015 352.255 ;
        RECT 5.605 350.965 6.815 351.715 ;
        RECT 2910.045 350.965 2910.335 351.690 ;
        RECT 2912.805 350.965 2914.015 351.715 ;
        RECT 5.520 350.795 6.900 350.965 ;
        RECT 2909.960 350.795 2910.420 350.965 ;
        RECT 2912.720 350.795 2914.100 350.965 ;
        RECT 5.605 350.045 6.815 350.795 ;
        RECT 2912.805 350.045 2914.015 350.795 ;
        RECT 5.605 349.505 6.125 350.045 ;
        RECT 2913.495 349.505 2914.015 350.045 ;
        RECT 5.605 346.275 6.125 346.815 ;
        RECT 2913.495 346.275 2914.015 346.815 ;
        RECT 5.605 345.525 6.815 346.275 ;
        RECT 2910.045 345.525 2910.335 346.250 ;
        RECT 2912.805 345.525 2914.015 346.275 ;
        RECT 5.520 345.355 6.900 345.525 ;
        RECT 2909.960 345.355 2910.420 345.525 ;
        RECT 2912.720 345.355 2914.100 345.525 ;
        RECT 5.605 344.605 6.815 345.355 ;
        RECT 2912.805 344.605 2914.015 345.355 ;
        RECT 5.605 344.065 6.125 344.605 ;
        RECT 2913.495 344.065 2914.015 344.605 ;
        RECT 5.605 340.835 6.125 341.375 ;
        RECT 2913.495 340.835 2914.015 341.375 ;
        RECT 5.605 340.085 6.815 340.835 ;
        RECT 2910.045 340.085 2910.335 340.810 ;
        RECT 2912.805 340.085 2914.015 340.835 ;
        RECT 5.520 339.915 6.900 340.085 ;
        RECT 2909.960 339.915 2910.420 340.085 ;
        RECT 2912.720 339.915 2914.100 340.085 ;
        RECT 5.605 339.165 6.815 339.915 ;
        RECT 2912.805 339.165 2914.015 339.915 ;
        RECT 5.605 338.625 6.125 339.165 ;
        RECT 2913.495 338.625 2914.015 339.165 ;
        RECT 5.605 335.395 6.125 335.935 ;
        RECT 2913.495 335.395 2914.015 335.935 ;
        RECT 5.605 334.645 6.815 335.395 ;
        RECT 2910.045 334.645 2910.335 335.370 ;
        RECT 2912.805 334.645 2914.015 335.395 ;
        RECT 5.520 334.475 6.900 334.645 ;
        RECT 2909.960 334.475 2910.420 334.645 ;
        RECT 2912.720 334.475 2914.100 334.645 ;
        RECT 5.605 333.725 6.815 334.475 ;
        RECT 2912.805 333.725 2914.015 334.475 ;
        RECT 5.605 333.185 6.125 333.725 ;
        RECT 2913.495 333.185 2914.015 333.725 ;
        RECT 5.605 329.955 6.125 330.495 ;
        RECT 2913.495 329.955 2914.015 330.495 ;
        RECT 5.605 329.205 6.815 329.955 ;
        RECT 2910.045 329.205 2910.335 329.930 ;
        RECT 2912.805 329.205 2914.015 329.955 ;
        RECT 5.520 329.035 6.900 329.205 ;
        RECT 2909.960 329.035 2910.420 329.205 ;
        RECT 2912.720 329.035 2914.100 329.205 ;
        RECT 5.605 328.285 6.815 329.035 ;
        RECT 2912.805 328.285 2914.015 329.035 ;
        RECT 5.605 327.745 6.125 328.285 ;
        RECT 2913.495 327.745 2914.015 328.285 ;
        RECT 5.605 324.515 6.125 325.055 ;
        RECT 2913.495 324.515 2914.015 325.055 ;
        RECT 5.605 323.765 6.815 324.515 ;
        RECT 2910.045 323.765 2910.335 324.490 ;
        RECT 2912.805 323.765 2914.015 324.515 ;
        RECT 5.520 323.595 6.900 323.765 ;
        RECT 2909.960 323.595 2910.420 323.765 ;
        RECT 2912.720 323.595 2914.100 323.765 ;
        RECT 5.605 322.845 6.815 323.595 ;
        RECT 2912.805 322.845 2914.015 323.595 ;
        RECT 5.605 322.305 6.125 322.845 ;
        RECT 2913.495 322.305 2914.015 322.845 ;
        RECT 5.605 319.075 6.125 319.615 ;
        RECT 2913.495 319.075 2914.015 319.615 ;
        RECT 5.605 318.325 6.815 319.075 ;
        RECT 2910.045 318.325 2910.335 319.050 ;
        RECT 2912.805 318.325 2914.015 319.075 ;
        RECT 5.520 318.155 6.900 318.325 ;
        RECT 2909.960 318.155 2910.420 318.325 ;
        RECT 2912.720 318.155 2914.100 318.325 ;
        RECT 5.605 317.405 6.815 318.155 ;
        RECT 2912.805 317.405 2914.015 318.155 ;
        RECT 5.605 316.865 6.125 317.405 ;
        RECT 2913.495 316.865 2914.015 317.405 ;
        RECT 5.605 313.635 6.125 314.175 ;
        RECT 2913.495 313.635 2914.015 314.175 ;
        RECT 5.605 312.885 6.815 313.635 ;
        RECT 9.515 312.885 9.855 313.545 ;
        RECT 2910.045 312.885 2910.335 313.610 ;
        RECT 2912.805 312.885 2914.015 313.635 ;
        RECT 5.520 312.715 6.900 312.885 ;
        RECT 8.740 312.715 10.120 312.885 ;
        RECT 2909.960 312.715 2910.420 312.885 ;
        RECT 2912.720 312.715 2914.100 312.885 ;
        RECT 5.605 311.965 6.815 312.715 ;
        RECT 2912.805 311.965 2914.015 312.715 ;
        RECT 5.605 311.425 6.125 311.965 ;
        RECT 2913.495 311.425 2914.015 311.965 ;
        RECT 5.605 308.195 6.125 308.735 ;
        RECT 2913.495 308.195 2914.015 308.735 ;
        RECT 5.605 307.445 6.815 308.195 ;
        RECT 2910.045 307.445 2910.335 308.170 ;
        RECT 2912.805 307.445 2914.015 308.195 ;
        RECT 5.520 307.275 6.900 307.445 ;
        RECT 2909.960 307.275 2910.420 307.445 ;
        RECT 2912.720 307.275 2914.100 307.445 ;
        RECT 5.605 306.525 6.815 307.275 ;
        RECT 2912.805 306.525 2914.015 307.275 ;
        RECT 5.605 305.985 6.125 306.525 ;
        RECT 2913.495 305.985 2914.015 306.525 ;
        RECT 5.605 302.755 6.125 303.295 ;
        RECT 2913.495 302.755 2914.015 303.295 ;
        RECT 5.605 302.005 6.815 302.755 ;
        RECT 2910.045 302.005 2910.335 302.730 ;
        RECT 2912.805 302.005 2914.015 302.755 ;
        RECT 5.520 301.835 6.900 302.005 ;
        RECT 2909.960 301.835 2910.420 302.005 ;
        RECT 2912.720 301.835 2914.100 302.005 ;
        RECT 5.605 301.085 6.815 301.835 ;
        RECT 2912.805 301.085 2914.015 301.835 ;
        RECT 5.605 300.545 6.125 301.085 ;
        RECT 2913.495 300.545 2914.015 301.085 ;
        RECT 5.605 297.315 6.125 297.855 ;
        RECT 2913.495 297.315 2914.015 297.855 ;
        RECT 5.605 296.565 6.815 297.315 ;
        RECT 2910.045 296.565 2910.335 297.290 ;
        RECT 2912.805 296.565 2914.015 297.315 ;
        RECT 5.520 296.395 6.900 296.565 ;
        RECT 2909.960 296.395 2910.420 296.565 ;
        RECT 2912.720 296.395 2914.100 296.565 ;
        RECT 5.605 295.645 6.815 296.395 ;
        RECT 2912.805 295.645 2914.015 296.395 ;
        RECT 5.605 295.105 6.125 295.645 ;
        RECT 2913.495 295.105 2914.015 295.645 ;
        RECT 5.605 291.875 6.125 292.415 ;
        RECT 2913.495 291.875 2914.015 292.415 ;
        RECT 5.605 291.125 6.815 291.875 ;
        RECT 2910.045 291.125 2910.335 291.850 ;
        RECT 2912.805 291.125 2914.015 291.875 ;
        RECT 5.520 290.955 6.900 291.125 ;
        RECT 2909.040 290.955 2910.420 291.125 ;
        RECT 2912.720 290.955 2914.100 291.125 ;
        RECT 5.605 290.205 6.815 290.955 ;
        RECT 2909.815 290.295 2910.155 290.955 ;
        RECT 2912.805 290.205 2914.015 290.955 ;
        RECT 5.605 289.665 6.125 290.205 ;
        RECT 2913.495 289.665 2914.015 290.205 ;
        RECT 5.605 286.435 6.125 286.975 ;
        RECT 2913.495 286.435 2914.015 286.975 ;
        RECT 5.605 285.685 6.815 286.435 ;
        RECT 2910.045 285.685 2910.335 286.410 ;
        RECT 2912.805 285.685 2914.015 286.435 ;
        RECT 5.520 285.515 6.900 285.685 ;
        RECT 2909.960 285.515 2910.420 285.685 ;
        RECT 2912.720 285.515 2914.100 285.685 ;
        RECT 5.605 284.765 6.815 285.515 ;
        RECT 2912.805 284.765 2914.015 285.515 ;
        RECT 5.605 284.225 6.125 284.765 ;
        RECT 2913.495 284.225 2914.015 284.765 ;
        RECT 5.605 280.995 6.125 281.535 ;
        RECT 2913.495 280.995 2914.015 281.535 ;
        RECT 5.605 280.245 6.815 280.995 ;
        RECT 2910.045 280.245 2910.335 280.970 ;
        RECT 2912.805 280.245 2914.015 280.995 ;
        RECT 5.520 280.075 6.900 280.245 ;
        RECT 2909.960 280.075 2910.420 280.245 ;
        RECT 2912.720 280.075 2914.100 280.245 ;
        RECT 5.605 279.325 6.815 280.075 ;
        RECT 2912.805 279.325 2914.015 280.075 ;
        RECT 5.605 278.785 6.125 279.325 ;
        RECT 2913.495 278.785 2914.015 279.325 ;
        RECT 5.605 275.555 6.125 276.095 ;
        RECT 2913.495 275.555 2914.015 276.095 ;
        RECT 5.605 274.805 6.815 275.555 ;
        RECT 2910.045 274.805 2910.335 275.530 ;
        RECT 2912.805 274.805 2914.015 275.555 ;
        RECT 5.520 274.635 6.900 274.805 ;
        RECT 2909.960 274.635 2910.420 274.805 ;
        RECT 2912.720 274.635 2914.100 274.805 ;
        RECT 5.605 273.885 6.815 274.635 ;
        RECT 2912.805 273.885 2914.015 274.635 ;
        RECT 5.605 273.345 6.125 273.885 ;
        RECT 2913.495 273.345 2914.015 273.885 ;
        RECT 5.605 270.115 6.125 270.655 ;
        RECT 2913.495 270.115 2914.015 270.655 ;
        RECT 5.605 269.365 6.815 270.115 ;
        RECT 2910.045 269.365 2910.335 270.090 ;
        RECT 2912.805 269.365 2914.015 270.115 ;
        RECT 5.520 269.195 6.900 269.365 ;
        RECT 2909.960 269.195 2910.420 269.365 ;
        RECT 2912.720 269.195 2914.100 269.365 ;
        RECT 5.605 268.445 6.815 269.195 ;
        RECT 2912.805 268.445 2914.015 269.195 ;
        RECT 5.605 267.905 6.125 268.445 ;
        RECT 2913.495 267.905 2914.015 268.445 ;
        RECT 5.605 264.675 6.125 265.215 ;
        RECT 2913.495 264.675 2914.015 265.215 ;
        RECT 5.605 263.925 6.815 264.675 ;
        RECT 2910.045 263.925 2910.335 264.650 ;
        RECT 2912.805 263.925 2914.015 264.675 ;
        RECT 5.520 263.755 6.900 263.925 ;
        RECT 2909.960 263.755 2910.420 263.925 ;
        RECT 2912.720 263.755 2914.100 263.925 ;
        RECT 5.605 263.005 6.815 263.755 ;
        RECT 2912.805 263.005 2914.015 263.755 ;
        RECT 5.605 262.465 6.125 263.005 ;
        RECT 2913.495 262.465 2914.015 263.005 ;
        RECT 5.605 259.235 6.125 259.775 ;
        RECT 2913.495 259.235 2914.015 259.775 ;
        RECT 5.605 258.485 6.815 259.235 ;
        RECT 2910.045 258.485 2910.335 259.210 ;
        RECT 2912.805 258.485 2914.015 259.235 ;
        RECT 5.520 258.315 6.900 258.485 ;
        RECT 2909.960 258.315 2910.420 258.485 ;
        RECT 2912.720 258.315 2914.100 258.485 ;
        RECT 5.605 257.565 6.815 258.315 ;
        RECT 2912.805 257.565 2914.015 258.315 ;
        RECT 5.605 257.025 6.125 257.565 ;
        RECT 2913.495 257.025 2914.015 257.565 ;
        RECT 5.605 253.795 6.125 254.335 ;
        RECT 2913.495 253.795 2914.015 254.335 ;
        RECT 5.605 253.045 6.815 253.795 ;
        RECT 2910.045 253.045 2910.335 253.770 ;
        RECT 2912.805 253.045 2914.015 253.795 ;
        RECT 5.520 252.875 6.900 253.045 ;
        RECT 2909.960 252.875 2910.420 253.045 ;
        RECT 2912.720 252.875 2914.100 253.045 ;
        RECT 5.605 252.125 6.815 252.875 ;
        RECT 2912.805 252.125 2914.015 252.875 ;
        RECT 5.605 251.585 6.125 252.125 ;
        RECT 2913.495 251.585 2914.015 252.125 ;
        RECT 5.605 248.355 6.125 248.895 ;
        RECT 2913.495 248.355 2914.015 248.895 ;
        RECT 5.605 247.605 6.815 248.355 ;
        RECT 2910.045 247.605 2910.335 248.330 ;
        RECT 2912.805 247.605 2914.015 248.355 ;
        RECT 5.520 247.435 6.900 247.605 ;
        RECT 2909.960 247.435 2910.420 247.605 ;
        RECT 2912.720 247.435 2914.100 247.605 ;
        RECT 5.605 246.685 6.815 247.435 ;
        RECT 2912.805 246.685 2914.015 247.435 ;
        RECT 5.605 246.145 6.125 246.685 ;
        RECT 2913.495 246.145 2914.015 246.685 ;
        RECT 5.605 242.915 6.125 243.455 ;
        RECT 2913.495 242.915 2914.015 243.455 ;
        RECT 5.605 242.165 6.815 242.915 ;
        RECT 2910.045 242.165 2910.335 242.890 ;
        RECT 2912.805 242.165 2914.015 242.915 ;
        RECT 5.520 241.995 6.900 242.165 ;
        RECT 2909.960 241.995 2910.420 242.165 ;
        RECT 2912.720 241.995 2914.100 242.165 ;
        RECT 5.605 241.245 6.815 241.995 ;
        RECT 2912.805 241.245 2914.015 241.995 ;
        RECT 5.605 240.705 6.125 241.245 ;
        RECT 2913.495 240.705 2914.015 241.245 ;
        RECT 5.605 237.475 6.125 238.015 ;
        RECT 2913.495 237.475 2914.015 238.015 ;
        RECT 5.605 236.725 6.815 237.475 ;
        RECT 2910.045 236.725 2910.335 237.450 ;
        RECT 2912.805 236.725 2914.015 237.475 ;
        RECT 5.520 236.555 6.900 236.725 ;
        RECT 2909.960 236.555 2910.420 236.725 ;
        RECT 2912.720 236.555 2914.100 236.725 ;
        RECT 5.605 235.805 6.815 236.555 ;
        RECT 2912.805 235.805 2914.015 236.555 ;
        RECT 5.605 235.265 6.125 235.805 ;
        RECT 2913.495 235.265 2914.015 235.805 ;
        RECT 5.605 232.035 6.125 232.575 ;
        RECT 2913.495 232.035 2914.015 232.575 ;
        RECT 5.605 231.285 6.815 232.035 ;
        RECT 2910.045 231.285 2910.335 232.010 ;
        RECT 2911.195 231.285 2911.535 231.945 ;
        RECT 2912.805 231.285 2914.015 232.035 ;
        RECT 5.520 231.115 6.900 231.285 ;
        RECT 2909.960 231.115 2911.800 231.285 ;
        RECT 2912.720 231.115 2914.100 231.285 ;
        RECT 5.605 230.365 6.815 231.115 ;
        RECT 2912.805 230.365 2914.015 231.115 ;
        RECT 5.605 229.825 6.125 230.365 ;
        RECT 2913.495 229.825 2914.015 230.365 ;
        RECT 5.605 226.595 6.125 227.135 ;
        RECT 2913.495 226.595 2914.015 227.135 ;
        RECT 5.605 225.845 6.815 226.595 ;
        RECT 2910.045 225.845 2910.335 226.570 ;
        RECT 2912.805 225.845 2914.015 226.595 ;
        RECT 5.520 225.675 6.900 225.845 ;
        RECT 2909.960 225.675 2910.420 225.845 ;
        RECT 2912.720 225.675 2914.100 225.845 ;
        RECT 5.605 224.925 6.815 225.675 ;
        RECT 2912.805 224.925 2914.015 225.675 ;
        RECT 5.605 224.385 6.125 224.925 ;
        RECT 2913.495 224.385 2914.015 224.925 ;
        RECT 5.605 221.155 6.125 221.695 ;
        RECT 2913.495 221.155 2914.015 221.695 ;
        RECT 5.605 220.405 6.815 221.155 ;
        RECT 2910.045 220.405 2910.335 221.130 ;
        RECT 2912.805 220.405 2914.015 221.155 ;
        RECT 5.520 220.235 6.900 220.405 ;
        RECT 2909.960 220.235 2910.420 220.405 ;
        RECT 2912.720 220.235 2914.100 220.405 ;
        RECT 5.605 219.485 6.815 220.235 ;
        RECT 2912.805 219.485 2914.015 220.235 ;
        RECT 5.605 218.945 6.125 219.485 ;
        RECT 2913.495 218.945 2914.015 219.485 ;
        RECT 5.605 215.715 6.125 216.255 ;
        RECT 2913.495 215.715 2914.015 216.255 ;
        RECT 5.605 214.965 6.815 215.715 ;
        RECT 2910.045 214.965 2910.335 215.690 ;
        RECT 2912.805 214.965 2914.015 215.715 ;
        RECT 5.520 214.795 6.900 214.965 ;
        RECT 2909.960 214.795 2910.420 214.965 ;
        RECT 2912.720 214.795 2914.100 214.965 ;
        RECT 5.605 214.045 6.815 214.795 ;
        RECT 2912.805 214.045 2914.015 214.795 ;
        RECT 5.605 213.505 6.125 214.045 ;
        RECT 2913.495 213.505 2914.015 214.045 ;
        RECT 5.605 210.275 6.125 210.815 ;
        RECT 2913.495 210.275 2914.015 210.815 ;
        RECT 5.605 209.525 6.815 210.275 ;
        RECT 2910.045 209.525 2910.335 210.250 ;
        RECT 2912.805 209.525 2914.015 210.275 ;
        RECT 5.520 209.355 6.900 209.525 ;
        RECT 2909.960 209.355 2910.420 209.525 ;
        RECT 2912.720 209.355 2914.100 209.525 ;
        RECT 5.605 208.605 6.815 209.355 ;
        RECT 2912.805 208.605 2914.015 209.355 ;
        RECT 5.605 208.065 6.125 208.605 ;
        RECT 2913.495 208.065 2914.015 208.605 ;
        RECT 5.605 204.835 6.125 205.375 ;
        RECT 2913.495 204.835 2914.015 205.375 ;
        RECT 5.605 204.085 6.815 204.835 ;
        RECT 2910.045 204.085 2910.335 204.810 ;
        RECT 2912.805 204.085 2914.015 204.835 ;
        RECT 5.520 203.915 6.900 204.085 ;
        RECT 2909.960 203.915 2910.420 204.085 ;
        RECT 2912.720 203.915 2914.100 204.085 ;
        RECT 5.605 203.165 6.815 203.915 ;
        RECT 2912.805 203.165 2914.015 203.915 ;
        RECT 5.605 202.625 6.125 203.165 ;
        RECT 2913.495 202.625 2914.015 203.165 ;
        RECT 5.605 199.395 6.125 199.935 ;
        RECT 2913.495 199.395 2914.015 199.935 ;
        RECT 5.605 198.645 6.815 199.395 ;
        RECT 2910.045 198.645 2910.335 199.370 ;
        RECT 2912.805 198.645 2914.015 199.395 ;
        RECT 5.520 198.475 6.900 198.645 ;
        RECT 2909.960 198.475 2910.420 198.645 ;
        RECT 2912.720 198.475 2914.100 198.645 ;
        RECT 5.605 197.725 6.815 198.475 ;
        RECT 2912.805 197.725 2914.015 198.475 ;
        RECT 5.605 197.185 6.125 197.725 ;
        RECT 2913.495 197.185 2914.015 197.725 ;
        RECT 5.605 193.955 6.125 194.495 ;
        RECT 2913.495 193.955 2914.015 194.495 ;
        RECT 5.605 193.205 6.815 193.955 ;
        RECT 2910.045 193.205 2910.335 193.930 ;
        RECT 2912.805 193.205 2914.015 193.955 ;
        RECT 5.520 193.035 6.900 193.205 ;
        RECT 2909.960 193.035 2910.420 193.205 ;
        RECT 2912.720 193.035 2914.100 193.205 ;
        RECT 5.605 192.285 6.815 193.035 ;
        RECT 2912.805 192.285 2914.015 193.035 ;
        RECT 5.605 191.745 6.125 192.285 ;
        RECT 2913.495 191.745 2914.015 192.285 ;
        RECT 5.605 188.515 6.125 189.055 ;
        RECT 2913.495 188.515 2914.015 189.055 ;
        RECT 5.605 187.765 6.815 188.515 ;
        RECT 2910.045 187.765 2910.335 188.490 ;
        RECT 2912.805 187.765 2914.015 188.515 ;
        RECT 5.520 187.595 6.900 187.765 ;
        RECT 2909.960 187.595 2910.420 187.765 ;
        RECT 2912.720 187.595 2914.100 187.765 ;
        RECT 5.605 186.845 6.815 187.595 ;
        RECT 2912.805 186.845 2914.015 187.595 ;
        RECT 5.605 186.305 6.125 186.845 ;
        RECT 2913.495 186.305 2914.015 186.845 ;
        RECT 5.605 183.075 6.125 183.615 ;
        RECT 2913.495 183.075 2914.015 183.615 ;
        RECT 5.605 182.325 6.815 183.075 ;
        RECT 2910.045 182.325 2910.335 183.050 ;
        RECT 2912.805 182.325 2914.015 183.075 ;
        RECT 5.520 182.155 6.900 182.325 ;
        RECT 2909.960 182.155 2910.420 182.325 ;
        RECT 2912.720 182.155 2914.100 182.325 ;
        RECT 5.605 181.405 6.815 182.155 ;
        RECT 2912.805 181.405 2914.015 182.155 ;
        RECT 5.605 180.865 6.125 181.405 ;
        RECT 2913.495 180.865 2914.015 181.405 ;
        RECT 5.605 177.635 6.125 178.175 ;
        RECT 2913.495 177.635 2914.015 178.175 ;
        RECT 5.605 176.885 6.815 177.635 ;
        RECT 2910.045 176.885 2910.335 177.610 ;
        RECT 2912.805 176.885 2914.015 177.635 ;
        RECT 5.520 176.715 6.900 176.885 ;
        RECT 2909.960 176.715 2910.420 176.885 ;
        RECT 2912.720 176.715 2914.100 176.885 ;
        RECT 5.605 175.965 6.815 176.715 ;
        RECT 2912.805 175.965 2914.015 176.715 ;
        RECT 5.605 175.425 6.125 175.965 ;
        RECT 2913.495 175.425 2914.015 175.965 ;
        RECT 5.605 172.195 6.125 172.735 ;
        RECT 2913.495 172.195 2914.015 172.735 ;
        RECT 5.605 171.445 6.815 172.195 ;
        RECT 2910.045 171.445 2910.335 172.170 ;
        RECT 2912.805 171.445 2914.015 172.195 ;
        RECT 5.520 171.275 6.900 171.445 ;
        RECT 2909.960 171.275 2910.420 171.445 ;
        RECT 2912.720 171.275 2914.100 171.445 ;
        RECT 5.605 170.525 6.815 171.275 ;
        RECT 2912.805 170.525 2914.015 171.275 ;
        RECT 5.605 169.985 6.125 170.525 ;
        RECT 2913.495 169.985 2914.015 170.525 ;
        RECT 5.605 166.755 6.125 167.295 ;
        RECT 2913.495 166.755 2914.015 167.295 ;
        RECT 5.605 166.005 6.815 166.755 ;
        RECT 2910.045 166.005 2910.335 166.730 ;
        RECT 2912.805 166.005 2914.015 166.755 ;
        RECT 5.520 165.835 6.900 166.005 ;
        RECT 2909.960 165.835 2910.420 166.005 ;
        RECT 2912.720 165.835 2914.100 166.005 ;
        RECT 5.605 165.085 6.815 165.835 ;
        RECT 2912.805 165.085 2914.015 165.835 ;
        RECT 5.605 164.545 6.125 165.085 ;
        RECT 2913.495 164.545 2914.015 165.085 ;
        RECT 5.605 161.315 6.125 161.855 ;
        RECT 2913.495 161.315 2914.015 161.855 ;
        RECT 5.605 160.565 6.815 161.315 ;
        RECT 2910.045 160.565 2910.335 161.290 ;
        RECT 2912.805 160.565 2914.015 161.315 ;
        RECT 5.520 160.395 6.900 160.565 ;
        RECT 2909.960 160.395 2910.420 160.565 ;
        RECT 2912.720 160.395 2914.100 160.565 ;
        RECT 5.605 159.645 6.815 160.395 ;
        RECT 2912.805 159.645 2914.015 160.395 ;
        RECT 5.605 159.105 6.125 159.645 ;
        RECT 2913.495 159.105 2914.015 159.645 ;
        RECT 5.605 155.875 6.125 156.415 ;
        RECT 2913.495 155.875 2914.015 156.415 ;
        RECT 5.605 155.125 6.815 155.875 ;
        RECT 2910.045 155.125 2910.335 155.850 ;
        RECT 2912.805 155.125 2914.015 155.875 ;
        RECT 5.520 154.955 6.900 155.125 ;
        RECT 2909.960 154.955 2910.420 155.125 ;
        RECT 2912.720 154.955 2914.100 155.125 ;
        RECT 5.605 154.205 6.815 154.955 ;
        RECT 2912.805 154.205 2914.015 154.955 ;
        RECT 5.605 153.665 6.125 154.205 ;
        RECT 2913.495 153.665 2914.015 154.205 ;
        RECT 5.605 150.435 6.125 150.975 ;
        RECT 2913.495 150.435 2914.015 150.975 ;
        RECT 5.605 149.685 6.815 150.435 ;
        RECT 2910.045 149.685 2910.335 150.410 ;
        RECT 2912.805 149.685 2914.015 150.435 ;
        RECT 5.520 149.515 6.900 149.685 ;
        RECT 2909.960 149.515 2910.420 149.685 ;
        RECT 2912.720 149.515 2914.100 149.685 ;
        RECT 5.605 148.765 6.815 149.515 ;
        RECT 2912.805 148.765 2914.015 149.515 ;
        RECT 5.605 148.225 6.125 148.765 ;
        RECT 2913.495 148.225 2914.015 148.765 ;
        RECT 5.605 144.995 6.125 145.535 ;
        RECT 2913.495 144.995 2914.015 145.535 ;
        RECT 5.605 144.245 6.815 144.995 ;
        RECT 2910.045 144.245 2910.335 144.970 ;
        RECT 2912.805 144.245 2914.015 144.995 ;
        RECT 5.520 144.075 6.900 144.245 ;
        RECT 2909.960 144.075 2910.420 144.245 ;
        RECT 2912.720 144.075 2914.100 144.245 ;
        RECT 5.605 143.325 6.815 144.075 ;
        RECT 2912.805 143.325 2914.015 144.075 ;
        RECT 5.605 142.785 6.125 143.325 ;
        RECT 2913.495 142.785 2914.015 143.325 ;
        RECT 5.605 139.555 6.125 140.095 ;
        RECT 2913.495 139.555 2914.015 140.095 ;
        RECT 5.605 138.805 6.815 139.555 ;
        RECT 2910.045 138.805 2910.335 139.530 ;
        RECT 2912.805 138.805 2914.015 139.555 ;
        RECT 5.520 138.635 6.900 138.805 ;
        RECT 2909.960 138.635 2910.420 138.805 ;
        RECT 2912.720 138.635 2914.100 138.805 ;
        RECT 5.605 137.885 6.815 138.635 ;
        RECT 2912.805 137.885 2914.015 138.635 ;
        RECT 5.605 137.345 6.125 137.885 ;
        RECT 2913.495 137.345 2914.015 137.885 ;
        RECT 5.605 134.115 6.125 134.655 ;
        RECT 2913.495 134.115 2914.015 134.655 ;
        RECT 5.605 133.365 6.815 134.115 ;
        RECT 2910.045 133.365 2910.335 134.090 ;
        RECT 2912.805 133.365 2914.015 134.115 ;
        RECT 5.520 133.195 6.900 133.365 ;
        RECT 2909.960 133.195 2910.420 133.365 ;
        RECT 2912.720 133.195 2914.100 133.365 ;
        RECT 5.605 132.445 6.815 133.195 ;
        RECT 2912.805 132.445 2914.015 133.195 ;
        RECT 5.605 131.905 6.125 132.445 ;
        RECT 2913.495 131.905 2914.015 132.445 ;
        RECT 5.605 128.675 6.125 129.215 ;
        RECT 2913.495 128.675 2914.015 129.215 ;
        RECT 5.605 127.925 6.815 128.675 ;
        RECT 2910.045 127.925 2910.335 128.650 ;
        RECT 2912.805 127.925 2914.015 128.675 ;
        RECT 5.520 127.755 13.700 127.925 ;
        RECT 2909.960 127.755 2910.420 127.925 ;
        RECT 2912.720 127.755 2914.100 127.925 ;
        RECT 5.605 127.005 6.815 127.755 ;
        RECT 7.415 127.375 7.745 127.755 ;
        RECT 8.355 127.295 8.605 127.755 ;
        RECT 10.300 127.255 10.670 127.755 ;
        RECT 12.525 127.225 12.695 127.755 ;
        RECT 13.525 127.275 13.695 127.755 ;
        RECT 2912.805 127.005 2914.015 127.755 ;
        RECT 5.605 126.465 6.125 127.005 ;
        RECT 2913.495 126.465 2914.015 127.005 ;
        RECT 5.605 123.235 6.125 123.775 ;
        RECT 2913.495 123.235 2914.015 123.775 ;
        RECT 5.605 122.485 6.815 123.235 ;
        RECT 2910.045 122.485 2910.335 123.210 ;
        RECT 2912.805 122.485 2914.015 123.235 ;
        RECT 5.520 122.315 6.900 122.485 ;
        RECT 2909.960 122.315 2910.420 122.485 ;
        RECT 2912.720 122.315 2914.100 122.485 ;
        RECT 5.605 121.565 6.815 122.315 ;
        RECT 2912.805 121.565 2914.015 122.315 ;
        RECT 5.605 121.025 6.125 121.565 ;
        RECT 2913.495 121.025 2914.015 121.565 ;
        RECT 5.605 117.795 6.125 118.335 ;
        RECT 2913.495 117.795 2914.015 118.335 ;
        RECT 5.605 117.045 6.815 117.795 ;
        RECT 2910.045 117.045 2910.335 117.770 ;
        RECT 2912.805 117.045 2914.015 117.795 ;
        RECT 5.520 116.875 6.900 117.045 ;
        RECT 2909.960 116.875 2910.420 117.045 ;
        RECT 2912.720 116.875 2914.100 117.045 ;
        RECT 5.605 116.125 6.815 116.875 ;
        RECT 2912.805 116.125 2914.015 116.875 ;
        RECT 5.605 115.585 6.125 116.125 ;
        RECT 2913.495 115.585 2914.015 116.125 ;
        RECT 5.605 112.355 6.125 112.895 ;
        RECT 2913.495 112.355 2914.015 112.895 ;
        RECT 5.605 111.605 6.815 112.355 ;
        RECT 2910.045 111.605 2910.335 112.330 ;
        RECT 2912.805 111.605 2914.015 112.355 ;
        RECT 5.520 111.435 6.900 111.605 ;
        RECT 2909.960 111.435 2910.420 111.605 ;
        RECT 2912.720 111.435 2914.100 111.605 ;
        RECT 5.605 110.685 6.815 111.435 ;
        RECT 2912.805 110.685 2914.015 111.435 ;
        RECT 5.605 110.145 6.125 110.685 ;
        RECT 2913.495 110.145 2914.015 110.685 ;
        RECT 5.605 106.915 6.125 107.455 ;
        RECT 2913.495 106.915 2914.015 107.455 ;
        RECT 5.605 106.165 6.815 106.915 ;
        RECT 2910.045 106.165 2910.335 106.890 ;
        RECT 2912.805 106.165 2914.015 106.915 ;
        RECT 5.520 105.995 6.900 106.165 ;
        RECT 8.740 105.995 10.120 106.165 ;
        RECT 2909.960 105.995 2910.420 106.165 ;
        RECT 2912.720 105.995 2914.100 106.165 ;
        RECT 5.605 105.245 6.815 105.995 ;
        RECT 5.605 104.705 6.125 105.245 ;
        RECT 8.865 105.175 9.095 105.995 ;
        RECT 9.765 105.175 9.975 105.995 ;
        RECT 2912.805 105.245 2914.015 105.995 ;
        RECT 2913.495 104.705 2914.015 105.245 ;
        RECT 5.605 101.475 6.125 102.015 ;
        RECT 2913.495 101.475 2914.015 102.015 ;
        RECT 5.605 100.725 6.815 101.475 ;
        RECT 2910.045 100.725 2910.335 101.450 ;
        RECT 2912.805 100.725 2914.015 101.475 ;
        RECT 5.520 100.555 6.900 100.725 ;
        RECT 2909.960 100.555 2910.420 100.725 ;
        RECT 2912.720 100.555 2914.100 100.725 ;
        RECT 5.605 99.805 6.815 100.555 ;
        RECT 2912.805 99.805 2914.015 100.555 ;
        RECT 5.605 99.265 6.125 99.805 ;
        RECT 2913.495 99.265 2914.015 99.805 ;
        RECT 5.605 96.035 6.125 96.575 ;
        RECT 2913.495 96.035 2914.015 96.575 ;
        RECT 5.605 95.285 6.815 96.035 ;
        RECT 2910.045 95.285 2910.335 96.010 ;
        RECT 2912.805 95.285 2914.015 96.035 ;
        RECT 5.520 95.115 6.900 95.285 ;
        RECT 2909.960 95.115 2910.420 95.285 ;
        RECT 2912.720 95.115 2914.100 95.285 ;
        RECT 5.605 94.365 6.815 95.115 ;
        RECT 2912.805 94.365 2914.015 95.115 ;
        RECT 5.605 93.825 6.125 94.365 ;
        RECT 2913.495 93.825 2914.015 94.365 ;
        RECT 5.605 90.595 6.125 91.135 ;
        RECT 2913.495 90.595 2914.015 91.135 ;
        RECT 5.605 89.845 6.815 90.595 ;
        RECT 2910.045 89.845 2910.335 90.570 ;
        RECT 2912.805 89.845 2914.015 90.595 ;
        RECT 5.520 89.675 6.900 89.845 ;
        RECT 2909.960 89.675 2910.420 89.845 ;
        RECT 2912.720 89.675 2914.100 89.845 ;
        RECT 5.605 88.925 6.815 89.675 ;
        RECT 2912.805 88.925 2914.015 89.675 ;
        RECT 5.605 88.385 6.125 88.925 ;
        RECT 2913.495 88.385 2914.015 88.925 ;
        RECT 5.605 85.155 6.125 85.695 ;
        RECT 2913.495 85.155 2914.015 85.695 ;
        RECT 5.605 84.405 6.815 85.155 ;
        RECT 2910.045 84.405 2910.335 85.130 ;
        RECT 2912.805 84.405 2914.015 85.155 ;
        RECT 5.520 84.235 6.900 84.405 ;
        RECT 2909.960 84.235 2910.420 84.405 ;
        RECT 2912.720 84.235 2914.100 84.405 ;
        RECT 5.605 83.485 6.815 84.235 ;
        RECT 2912.805 83.485 2914.015 84.235 ;
        RECT 5.605 82.945 6.125 83.485 ;
        RECT 2913.495 82.945 2914.015 83.485 ;
        RECT 5.605 79.715 6.125 80.255 ;
        RECT 2913.495 79.715 2914.015 80.255 ;
        RECT 5.605 78.965 6.815 79.715 ;
        RECT 2910.045 78.965 2910.335 79.690 ;
        RECT 2912.805 78.965 2914.015 79.715 ;
        RECT 5.520 78.795 6.900 78.965 ;
        RECT 2909.960 78.795 2910.420 78.965 ;
        RECT 2912.720 78.795 2914.100 78.965 ;
        RECT 5.605 78.045 6.815 78.795 ;
        RECT 2912.805 78.045 2914.015 78.795 ;
        RECT 5.605 77.505 6.125 78.045 ;
        RECT 2913.495 77.505 2914.015 78.045 ;
        RECT 5.605 74.275 6.125 74.815 ;
        RECT 2913.495 74.275 2914.015 74.815 ;
        RECT 5.605 73.525 6.815 74.275 ;
        RECT 2910.045 73.525 2910.335 74.250 ;
        RECT 2912.805 73.525 2914.015 74.275 ;
        RECT 5.520 73.355 6.900 73.525 ;
        RECT 2909.960 73.355 2910.420 73.525 ;
        RECT 2912.720 73.355 2914.100 73.525 ;
        RECT 5.605 72.605 6.815 73.355 ;
        RECT 2912.805 72.605 2914.015 73.355 ;
        RECT 5.605 72.065 6.125 72.605 ;
        RECT 2913.495 72.065 2914.015 72.605 ;
        RECT 5.605 68.835 6.125 69.375 ;
        RECT 2913.495 68.835 2914.015 69.375 ;
        RECT 5.605 68.085 6.815 68.835 ;
        RECT 2910.045 68.085 2910.335 68.810 ;
        RECT 2912.805 68.085 2914.015 68.835 ;
        RECT 5.520 67.915 6.900 68.085 ;
        RECT 2909.960 67.915 2910.420 68.085 ;
        RECT 2912.720 67.915 2914.100 68.085 ;
        RECT 5.605 67.165 6.815 67.915 ;
        RECT 2912.805 67.165 2914.015 67.915 ;
        RECT 5.605 66.625 6.125 67.165 ;
        RECT 2913.495 66.625 2914.015 67.165 ;
        RECT 5.605 63.395 6.125 63.935 ;
        RECT 2913.495 63.395 2914.015 63.935 ;
        RECT 5.605 62.645 6.815 63.395 ;
        RECT 2910.045 62.645 2910.335 63.370 ;
        RECT 2912.805 62.645 2914.015 63.395 ;
        RECT 5.520 62.475 6.900 62.645 ;
        RECT 2909.040 62.475 2910.420 62.645 ;
        RECT 2912.720 62.475 2914.100 62.645 ;
        RECT 5.605 61.725 6.815 62.475 ;
        RECT 2909.815 61.815 2910.155 62.475 ;
        RECT 2912.805 61.725 2914.015 62.475 ;
        RECT 5.605 61.185 6.125 61.725 ;
        RECT 2913.495 61.185 2914.015 61.725 ;
        RECT 5.605 57.955 6.125 58.495 ;
        RECT 2913.495 57.955 2914.015 58.495 ;
        RECT 5.605 57.205 6.815 57.955 ;
        RECT 2910.045 57.205 2910.335 57.930 ;
        RECT 2912.805 57.205 2914.015 57.955 ;
        RECT 5.520 57.035 6.900 57.205 ;
        RECT 2909.960 57.035 2910.420 57.205 ;
        RECT 2912.720 57.035 2914.100 57.205 ;
        RECT 5.605 56.285 6.815 57.035 ;
        RECT 2912.805 56.285 2914.015 57.035 ;
        RECT 5.605 55.745 6.125 56.285 ;
        RECT 2913.495 55.745 2914.015 56.285 ;
        RECT 5.605 52.515 6.125 53.055 ;
        RECT 2913.495 52.515 2914.015 53.055 ;
        RECT 5.605 51.765 6.815 52.515 ;
        RECT 2910.045 51.765 2910.335 52.490 ;
        RECT 2912.805 51.765 2914.015 52.515 ;
        RECT 5.520 51.595 6.900 51.765 ;
        RECT 2909.960 51.595 2910.420 51.765 ;
        RECT 2912.720 51.595 2914.100 51.765 ;
        RECT 5.605 50.845 6.815 51.595 ;
        RECT 2912.805 50.845 2914.015 51.595 ;
        RECT 5.605 50.305 6.125 50.845 ;
        RECT 2913.495 50.305 2914.015 50.845 ;
        RECT 5.605 47.075 6.125 47.615 ;
        RECT 2913.495 47.075 2914.015 47.615 ;
        RECT 5.605 46.325 6.815 47.075 ;
        RECT 2910.045 46.325 2910.335 47.050 ;
        RECT 2912.805 46.325 2914.015 47.075 ;
        RECT 5.520 46.155 6.900 46.325 ;
        RECT 2909.960 46.155 2910.420 46.325 ;
        RECT 2912.720 46.155 2914.100 46.325 ;
        RECT 5.605 45.405 6.815 46.155 ;
        RECT 2912.805 45.405 2914.015 46.155 ;
        RECT 5.605 44.865 6.125 45.405 ;
        RECT 2913.495 44.865 2914.015 45.405 ;
        RECT 5.605 41.635 6.125 42.175 ;
        RECT 2913.495 41.635 2914.015 42.175 ;
        RECT 5.605 40.885 6.815 41.635 ;
        RECT 7.415 40.885 7.745 41.265 ;
        RECT 8.355 40.885 8.605 41.345 ;
        RECT 10.300 40.885 10.670 41.385 ;
        RECT 12.525 40.885 12.695 41.415 ;
        RECT 13.525 40.885 13.695 41.365 ;
        RECT 2910.045 40.885 2910.335 41.610 ;
        RECT 2912.805 40.885 2914.015 41.635 ;
        RECT 5.520 40.715 13.700 40.885 ;
        RECT 2909.960 40.715 2910.420 40.885 ;
        RECT 2912.720 40.715 2914.100 40.885 ;
        RECT 5.605 39.965 6.815 40.715 ;
        RECT 2912.805 39.965 2914.015 40.715 ;
        RECT 5.605 39.425 6.125 39.965 ;
        RECT 2913.495 39.425 2914.015 39.965 ;
        RECT 5.605 36.195 6.125 36.735 ;
        RECT 2913.495 36.195 2914.015 36.735 ;
        RECT 5.605 35.445 6.815 36.195 ;
        RECT 2910.045 35.445 2910.335 36.170 ;
        RECT 2912.805 35.445 2914.015 36.195 ;
        RECT 5.520 35.275 6.900 35.445 ;
        RECT 2909.960 35.275 2910.420 35.445 ;
        RECT 2912.720 35.275 2914.100 35.445 ;
        RECT 5.605 34.525 6.815 35.275 ;
        RECT 2912.805 34.525 2914.015 35.275 ;
        RECT 5.605 33.985 6.125 34.525 ;
        RECT 2913.495 33.985 2914.015 34.525 ;
        RECT 5.605 30.755 6.125 31.295 ;
        RECT 2913.495 30.755 2914.015 31.295 ;
        RECT 5.605 30.005 6.815 30.755 ;
        RECT 2910.045 30.005 2910.335 30.730 ;
        RECT 2912.805 30.005 2914.015 30.755 ;
        RECT 5.520 29.835 6.900 30.005 ;
        RECT 2909.960 29.835 2910.420 30.005 ;
        RECT 2912.720 29.835 2914.100 30.005 ;
        RECT 5.605 29.085 6.815 29.835 ;
        RECT 2912.805 29.085 2914.015 29.835 ;
        RECT 5.605 28.545 6.125 29.085 ;
        RECT 2913.495 28.545 2914.015 29.085 ;
        RECT 5.605 25.315 6.125 25.855 ;
        RECT 2913.495 25.315 2914.015 25.855 ;
        RECT 5.605 24.565 6.815 25.315 ;
        RECT 2910.045 24.565 2910.335 25.290 ;
        RECT 2912.805 24.565 2914.015 25.315 ;
        RECT 5.520 24.395 6.900 24.565 ;
        RECT 2909.960 24.395 2910.420 24.565 ;
        RECT 2912.720 24.395 2914.100 24.565 ;
        RECT 5.605 23.645 6.815 24.395 ;
        RECT 2912.805 23.645 2914.015 24.395 ;
        RECT 5.605 23.105 6.125 23.645 ;
        RECT 2913.495 23.105 2914.015 23.645 ;
        RECT 5.605 19.875 6.125 20.415 ;
        RECT 5.605 19.125 6.815 19.875 ;
        RECT 7.075 19.125 7.245 19.935 ;
        RECT 8.755 19.125 8.925 19.595 ;
        RECT 9.595 19.125 10.285 19.595 ;
        RECT 10.955 19.125 11.125 19.595 ;
        RECT 11.795 19.125 11.965 19.935 ;
        RECT 2913.495 19.875 2914.015 20.415 ;
        RECT 12.635 19.125 12.805 19.595 ;
        RECT 13.475 19.125 13.645 19.595 ;
        RECT 2910.045 19.125 2910.335 19.850 ;
        RECT 2912.805 19.125 2914.015 19.875 ;
        RECT 5.520 18.955 13.700 19.125 ;
        RECT 2909.040 18.955 2911.800 19.125 ;
        RECT 2912.720 18.955 2914.100 19.125 ;
        RECT 5.605 18.205 6.815 18.955 ;
        RECT 7.415 18.575 7.745 18.955 ;
        RECT 8.355 18.495 8.605 18.955 ;
        RECT 10.300 18.455 10.670 18.955 ;
        RECT 12.525 18.425 12.695 18.955 ;
        RECT 13.525 18.475 13.695 18.955 ;
        RECT 2909.815 18.295 2910.155 18.955 ;
        RECT 2911.195 18.295 2911.535 18.955 ;
        RECT 2912.805 18.205 2914.015 18.955 ;
        RECT 5.605 17.665 6.125 18.205 ;
        RECT 2913.495 17.665 2914.015 18.205 ;
        RECT 5.605 14.435 6.125 14.975 ;
        RECT 2913.495 14.435 2914.015 14.975 ;
        RECT 5.605 13.685 6.815 14.435 ;
        RECT 7.415 13.685 7.745 14.065 ;
        RECT 8.355 13.685 8.605 14.145 ;
        RECT 10.300 13.685 10.670 14.185 ;
        RECT 12.525 13.685 12.695 14.215 ;
        RECT 13.525 13.685 13.695 14.165 ;
        RECT 14.395 13.685 14.565 13.700 ;
        RECT 15.245 13.685 15.415 13.700 ;
        RECT 17.120 13.685 17.450 13.700 ;
        RECT 18.050 13.685 18.310 13.700 ;
        RECT 19.865 13.685 20.155 13.700 ;
        RECT 47.925 13.685 48.215 13.700 ;
        RECT 58.085 13.685 58.315 13.700 ;
        RECT 58.985 13.685 59.195 13.700 ;
        RECT 59.600 13.685 59.770 13.700 ;
        RECT 60.440 13.685 60.610 13.700 ;
        RECT 61.280 13.685 61.450 13.700 ;
        RECT 63.980 13.685 64.150 13.700 ;
        RECT 64.820 13.685 64.990 13.700 ;
        RECT 75.985 13.685 76.275 13.700 ;
        RECT 79.185 13.685 79.515 13.700 ;
        RECT 80.090 13.685 80.420 13.700 ;
        RECT 80.950 13.685 81.280 13.700 ;
        RECT 83.315 13.685 83.645 13.700 ;
        RECT 84.255 13.685 84.505 13.700 ;
        RECT 86.200 13.685 86.570 13.700 ;
        RECT 88.425 13.685 88.595 13.700 ;
        RECT 89.425 13.685 89.595 13.700 ;
        RECT 90.295 13.685 90.465 13.700 ;
        RECT 91.145 13.685 91.315 13.700 ;
        RECT 101.760 13.685 102.090 13.700 ;
        RECT 102.690 13.685 102.950 13.700 ;
        RECT 104.045 13.685 104.335 13.700 ;
        RECT 104.595 13.685 104.765 13.700 ;
        RECT 106.275 13.685 106.445 13.700 ;
        RECT 107.115 13.685 107.805 13.700 ;
        RECT 108.475 13.685 108.645 13.700 ;
        RECT 109.315 13.685 109.485 13.700 ;
        RECT 110.155 13.685 110.325 13.700 ;
        RECT 110.995 13.685 111.165 13.700 ;
        RECT 120.185 13.685 120.415 13.700 ;
        RECT 121.085 13.685 121.295 13.700 ;
        RECT 132.105 13.685 132.395 13.700 ;
        RECT 134.580 13.685 134.750 13.700 ;
        RECT 135.420 13.685 135.590 13.700 ;
        RECT 136.260 13.685 136.430 13.700 ;
        RECT 138.960 13.685 139.130 13.700 ;
        RECT 139.800 13.685 139.970 13.700 ;
        RECT 144.165 13.685 144.475 13.700 ;
        RECT 145.015 13.685 145.345 13.700 ;
        RECT 145.855 13.685 146.185 13.700 ;
        RECT 146.840 13.685 147.170 13.700 ;
        RECT 147.770 13.685 148.030 13.700 ;
        RECT 152.895 13.685 153.065 13.700 ;
        RECT 154.575 13.685 154.745 13.700 ;
        RECT 155.415 13.685 156.105 13.700 ;
        RECT 156.775 13.685 156.945 13.700 ;
        RECT 157.615 13.685 157.785 13.700 ;
        RECT 158.455 13.685 158.625 13.700 ;
        RECT 159.295 13.685 159.465 13.700 ;
        RECT 160.165 13.685 160.455 13.700 ;
        RECT 160.665 13.685 160.895 13.700 ;
        RECT 161.565 13.685 161.775 13.700 ;
        RECT 162.895 13.685 163.225 13.700 ;
        RECT 163.835 13.685 164.085 13.700 ;
        RECT 165.780 13.685 166.150 13.700 ;
        RECT 168.005 13.685 168.175 13.700 ;
        RECT 169.005 13.685 169.175 13.700 ;
        RECT 169.875 13.685 170.045 13.700 ;
        RECT 170.725 13.685 170.895 13.700 ;
        RECT 181.500 13.685 181.670 13.700 ;
        RECT 182.340 13.685 182.510 13.700 ;
        RECT 183.180 13.685 183.350 13.700 ;
        RECT 185.880 13.685 186.050 13.700 ;
        RECT 186.720 13.685 186.890 13.700 ;
        RECT 188.225 13.685 188.515 13.700 ;
        RECT 196.025 13.685 196.355 13.700 ;
        RECT 196.930 13.685 197.260 13.700 ;
        RECT 197.790 13.685 198.120 13.700 ;
        RECT 200.165 13.685 200.495 13.700 ;
        RECT 201.070 13.685 201.400 13.700 ;
        RECT 201.930 13.685 202.260 13.700 ;
        RECT 208.555 13.685 208.725 13.700 ;
        RECT 210.235 13.685 210.405 13.700 ;
        RECT 211.075 13.685 211.765 13.700 ;
        RECT 212.435 13.685 212.605 13.700 ;
        RECT 213.275 13.685 213.445 13.700 ;
        RECT 214.115 13.685 214.285 13.700 ;
        RECT 214.955 13.685 215.125 13.700 ;
        RECT 216.285 13.685 216.575 13.700 ;
        RECT 218.300 13.685 218.470 13.700 ;
        RECT 219.140 13.685 219.310 13.700 ;
        RECT 219.980 13.685 220.150 13.700 ;
        RECT 222.680 13.685 222.850 13.700 ;
        RECT 223.520 13.685 223.690 13.700 ;
        RECT 228.215 13.685 228.545 13.700 ;
        RECT 229.155 13.685 229.405 13.700 ;
        RECT 231.100 13.685 231.470 13.700 ;
        RECT 233.325 13.685 233.495 13.700 ;
        RECT 234.325 13.685 234.495 13.700 ;
        RECT 235.195 13.685 235.365 13.700 ;
        RECT 236.045 13.685 236.215 13.700 ;
        RECT 237.075 13.685 237.245 13.700 ;
        RECT 238.755 13.685 238.925 13.700 ;
        RECT 239.595 13.685 240.285 13.700 ;
        RECT 240.955 13.685 241.125 13.700 ;
        RECT 241.795 13.685 241.965 13.700 ;
        RECT 242.635 13.685 242.805 13.700 ;
        RECT 243.475 13.685 243.645 13.700 ;
        RECT 244.345 13.685 244.635 13.700 ;
        RECT 259.495 13.685 259.825 13.700 ;
        RECT 260.435 13.685 260.685 13.700 ;
        RECT 262.380 13.685 262.750 13.700 ;
        RECT 264.605 13.685 264.775 13.700 ;
        RECT 265.605 13.685 265.775 13.700 ;
        RECT 266.475 13.685 266.645 13.700 ;
        RECT 267.325 13.685 267.495 13.700 ;
        RECT 268.280 13.685 268.610 13.700 ;
        RECT 269.210 13.685 269.470 13.700 ;
        RECT 272.405 13.685 272.695 13.700 ;
        RECT 277.505 13.685 277.735 13.700 ;
        RECT 278.405 13.685 278.615 13.700 ;
        RECT 283.460 13.685 283.790 13.700 ;
        RECT 284.390 13.685 284.650 13.700 ;
        RECT 289.005 13.685 289.235 13.700 ;
        RECT 289.905 13.685 290.115 13.700 ;
        RECT 292.820 13.685 292.990 13.700 ;
        RECT 293.660 13.685 293.830 13.700 ;
        RECT 294.500 13.685 294.670 13.700 ;
        RECT 297.200 13.685 297.370 13.700 ;
        RECT 298.040 13.685 298.210 13.700 ;
        RECT 300.465 13.685 300.755 13.700 ;
        RECT 304.645 13.685 304.875 13.700 ;
        RECT 305.545 13.685 305.755 13.700 ;
        RECT 306.025 13.685 306.255 13.700 ;
        RECT 306.925 13.685 307.135 13.700 ;
        RECT 308.300 13.685 308.630 13.700 ;
        RECT 309.230 13.685 309.490 13.700 ;
        RECT 310.140 13.685 310.470 13.700 ;
        RECT 311.070 13.685 311.330 13.700 ;
        RECT 314.305 13.685 314.535 13.700 ;
        RECT 315.205 13.685 315.415 13.700 ;
        RECT 317.915 13.685 318.245 13.700 ;
        RECT 318.855 13.685 319.105 13.700 ;
        RECT 320.800 13.685 321.170 13.700 ;
        RECT 323.025 13.685 323.195 13.700 ;
        RECT 324.025 13.685 324.195 13.700 ;
        RECT 324.895 13.685 325.065 13.700 ;
        RECT 325.745 13.685 325.915 13.700 ;
        RECT 328.525 13.685 328.815 13.700 ;
        RECT 329.415 13.685 329.745 13.700 ;
        RECT 330.355 13.685 330.605 13.700 ;
        RECT 332.300 13.685 332.670 13.700 ;
        RECT 334.525 13.685 334.695 13.700 ;
        RECT 335.525 13.685 335.695 13.700 ;
        RECT 336.395 13.685 336.565 13.700 ;
        RECT 337.245 13.685 337.415 13.700 ;
        RECT 339.580 13.685 339.910 13.700 ;
        RECT 340.510 13.685 340.770 13.700 ;
        RECT 348.275 13.685 348.605 13.700 ;
        RECT 349.215 13.685 349.465 13.700 ;
        RECT 351.160 13.685 351.530 13.700 ;
        RECT 353.385 13.685 353.555 13.700 ;
        RECT 354.385 13.685 354.555 13.700 ;
        RECT 355.255 13.685 355.425 13.700 ;
        RECT 356.105 13.685 356.275 13.700 ;
        RECT 356.585 13.685 356.875 13.700 ;
        RECT 357.520 13.685 357.850 13.700 ;
        RECT 358.450 13.685 358.710 13.700 ;
        RECT 359.895 13.685 360.065 13.700 ;
        RECT 361.575 13.685 361.745 13.700 ;
        RECT 362.415 13.685 363.105 13.700 ;
        RECT 363.775 13.685 363.945 13.700 ;
        RECT 364.615 13.685 364.785 13.700 ;
        RECT 365.455 13.685 365.625 13.700 ;
        RECT 366.295 13.685 366.465 13.700 ;
        RECT 368.175 13.685 368.345 13.700 ;
        RECT 369.855 13.685 370.025 13.700 ;
        RECT 370.695 13.685 371.385 13.700 ;
        RECT 372.055 13.685 372.225 13.700 ;
        RECT 372.895 13.685 373.065 13.700 ;
        RECT 373.735 13.685 373.905 13.700 ;
        RECT 374.575 13.685 374.745 13.700 ;
        RECT 384.645 13.685 384.935 13.700 ;
        RECT 385.195 13.685 385.365 13.700 ;
        RECT 386.875 13.685 387.045 13.700 ;
        RECT 387.715 13.685 388.405 13.700 ;
        RECT 389.075 13.685 389.245 13.700 ;
        RECT 389.915 13.685 390.085 13.700 ;
        RECT 390.755 13.685 390.925 13.700 ;
        RECT 391.595 13.685 391.765 13.700 ;
        RECT 394.320 13.685 394.650 13.700 ;
        RECT 395.250 13.685 395.510 13.700 ;
        RECT 396.115 13.685 396.445 13.700 ;
        RECT 397.055 13.685 397.305 13.700 ;
        RECT 399.000 13.685 399.370 13.700 ;
        RECT 401.225 13.685 401.395 13.700 ;
        RECT 402.225 13.685 402.395 13.700 ;
        RECT 403.095 13.685 403.265 13.700 ;
        RECT 403.945 13.685 404.115 13.700 ;
        RECT 412.705 13.685 412.995 13.700 ;
        RECT 413.715 13.685 413.885 13.700 ;
        RECT 415.395 13.685 415.565 13.700 ;
        RECT 416.235 13.685 416.925 13.700 ;
        RECT 417.595 13.685 417.765 13.700 ;
        RECT 418.435 13.685 418.605 13.700 ;
        RECT 419.275 13.685 419.445 13.700 ;
        RECT 420.115 13.685 420.285 13.700 ;
        RECT 426.015 13.685 426.345 13.700 ;
        RECT 426.955 13.685 427.205 13.700 ;
        RECT 428.900 13.685 429.270 13.700 ;
        RECT 431.125 13.685 431.295 13.700 ;
        RECT 432.125 13.685 432.295 13.700 ;
        RECT 432.995 13.685 433.165 13.700 ;
        RECT 433.845 13.685 434.015 13.700 ;
        RECT 440.765 13.685 441.055 13.700 ;
        RECT 445.795 13.685 446.125 13.700 ;
        RECT 446.735 13.685 446.985 13.700 ;
        RECT 448.680 13.685 449.050 13.700 ;
        RECT 450.905 13.685 451.075 13.700 ;
        RECT 451.905 13.685 452.075 13.700 ;
        RECT 452.775 13.685 452.945 13.700 ;
        RECT 453.625 13.685 453.795 13.700 ;
        RECT 458.215 13.685 458.545 13.700 ;
        RECT 459.155 13.685 459.405 13.700 ;
        RECT 461.100 13.685 461.470 13.700 ;
        RECT 463.325 13.685 463.495 13.700 ;
        RECT 464.325 13.685 464.495 13.700 ;
        RECT 465.195 13.685 465.365 13.700 ;
        RECT 466.045 13.685 466.215 13.700 ;
        RECT 467.460 13.685 467.790 13.700 ;
        RECT 468.390 13.685 468.650 13.700 ;
        RECT 468.825 13.685 469.115 13.700 ;
        RECT 481.260 13.685 481.590 13.700 ;
        RECT 482.190 13.685 482.450 13.700 ;
        RECT 494.625 13.685 494.855 13.700 ;
        RECT 495.525 13.685 495.735 13.700 ;
        RECT 496.885 13.685 497.175 13.700 ;
        RECT 524.945 13.685 525.235 13.700 ;
        RECT 527.880 13.685 528.050 13.700 ;
        RECT 528.720 13.685 528.890 13.700 ;
        RECT 529.560 13.685 529.730 13.700 ;
        RECT 532.260 13.685 532.430 13.700 ;
        RECT 533.100 13.685 533.270 13.700 ;
        RECT 536.025 13.685 536.255 13.700 ;
        RECT 536.925 13.685 537.135 13.700 ;
        RECT 539.220 13.685 539.550 13.700 ;
        RECT 540.150 13.685 540.410 13.700 ;
        RECT 553.005 13.685 553.295 13.700 ;
        RECT 564.520 13.685 564.850 13.700 ;
        RECT 565.450 13.685 565.710 13.700 ;
        RECT 572.295 13.685 572.625 13.700 ;
        RECT 573.235 13.685 573.485 13.700 ;
        RECT 575.180 13.685 575.550 13.700 ;
        RECT 577.405 13.685 577.575 13.700 ;
        RECT 578.405 13.685 578.575 13.700 ;
        RECT 579.275 13.685 579.445 13.700 ;
        RECT 580.125 13.685 580.295 13.700 ;
        RECT 581.065 13.685 581.355 13.700 ;
        RECT 609.125 13.685 609.415 13.700 ;
        RECT 637.185 13.685 637.475 13.700 ;
        RECT 665.245 13.685 665.535 13.700 ;
        RECT 693.305 13.685 693.595 13.700 ;
        RECT 721.365 13.685 721.655 13.700 ;
        RECT 749.425 13.685 749.715 13.700 ;
        RECT 777.485 13.685 777.775 13.700 ;
        RECT 805.545 13.685 805.835 13.700 ;
        RECT 833.605 13.685 833.895 13.700 ;
        RECT 861.665 13.685 861.955 13.700 ;
        RECT 889.725 13.685 890.015 13.700 ;
        RECT 917.785 13.685 918.075 13.700 ;
        RECT 945.845 13.685 946.135 13.700 ;
        RECT 973.905 13.685 974.195 13.700 ;
        RECT 1001.965 13.685 1002.255 13.700 ;
        RECT 1030.025 13.685 1030.315 13.700 ;
        RECT 1058.085 13.685 1058.375 13.700 ;
        RECT 1086.145 13.685 1086.435 13.700 ;
        RECT 1114.205 13.685 1114.495 13.700 ;
        RECT 1142.265 13.685 1142.555 13.700 ;
        RECT 1170.325 13.685 1170.615 13.700 ;
        RECT 1198.385 13.685 1198.675 13.700 ;
        RECT 1226.445 13.685 1226.735 13.700 ;
        RECT 1254.505 13.685 1254.795 13.700 ;
        RECT 1282.565 13.685 1282.855 13.700 ;
        RECT 1310.625 13.685 1310.915 13.700 ;
        RECT 1338.685 13.685 1338.975 13.700 ;
        RECT 1366.745 13.685 1367.035 13.700 ;
        RECT 1383.075 13.685 1383.415 13.700 ;
        RECT 1394.805 13.685 1395.095 13.700 ;
        RECT 1401.475 13.685 1401.815 13.700 ;
        RECT 1422.865 13.685 1423.155 13.700 ;
        RECT 1450.925 13.685 1451.215 13.700 ;
        RECT 1478.985 13.685 1479.275 13.700 ;
        RECT 1504.515 13.685 1504.855 13.700 ;
        RECT 1507.045 13.685 1507.335 13.700 ;
        RECT 1526.595 13.685 1526.935 13.700 ;
        RECT 1535.105 13.685 1535.395 13.700 ;
        RECT 1536.255 13.685 1536.595 13.700 ;
        RECT 1539.935 13.685 1540.275 13.700 ;
        RECT 1543.155 13.685 1543.495 13.700 ;
        RECT 1559.715 13.685 1560.055 13.700 ;
        RECT 1563.165 13.685 1563.455 13.700 ;
        RECT 1576.275 13.685 1576.615 13.700 ;
        RECT 1589.155 13.685 1589.495 13.700 ;
        RECT 1591.225 13.685 1591.515 13.700 ;
        RECT 1619.285 13.685 1619.575 13.700 ;
        RECT 1626.415 13.685 1626.755 13.700 ;
        RECT 1647.345 13.685 1647.635 13.700 ;
        RECT 1649.415 13.685 1649.755 13.700 ;
        RECT 1675.405 13.685 1675.695 13.700 ;
        RECT 1703.465 13.685 1703.755 13.700 ;
        RECT 1731.525 13.685 1731.815 13.700 ;
        RECT 1759.585 13.685 1759.875 13.700 ;
        RECT 1760.735 13.685 1761.075 13.700 ;
        RECT 1774.535 13.685 1774.875 13.700 ;
        RECT 1787.645 13.685 1787.935 13.700 ;
        RECT 1815.705 13.685 1815.995 13.700 ;
        RECT 1830.655 13.685 1830.995 13.700 ;
        RECT 1843.765 13.685 1844.055 13.700 ;
        RECT 1871.825 13.685 1872.115 13.700 ;
        RECT 1899.885 13.685 1900.175 13.700 ;
        RECT 1913.915 13.685 1914.255 13.700 ;
        RECT 1926.335 13.685 1926.675 13.700 ;
        RECT 1927.945 13.685 1928.235 13.700 ;
        RECT 1932.315 13.685 1932.655 13.700 ;
        RECT 1948.415 13.685 1948.755 13.700 ;
        RECT 1956.005 13.685 1956.295 13.700 ;
        RECT 1973.715 13.685 1974.055 13.700 ;
        RECT 1983.375 13.685 1983.715 13.700 ;
        RECT 1984.065 13.685 1984.355 13.700 ;
        RECT 1992.575 13.685 1992.915 13.700 ;
        RECT 1995.795 13.685 1996.135 13.700 ;
        RECT 2000.395 13.685 2000.735 13.700 ;
        RECT 2012.125 13.685 2012.415 13.700 ;
        RECT 2018.795 13.685 2019.135 13.700 ;
        RECT 2025.235 13.685 2025.575 13.700 ;
        RECT 2038.115 13.685 2038.455 13.700 ;
        RECT 2040.185 13.685 2040.475 13.700 ;
        RECT 2059.735 13.685 2060.075 13.700 ;
        RECT 2061.115 13.685 2061.455 13.700 ;
        RECT 2068.245 13.685 2068.535 13.700 ;
        RECT 2074.455 13.685 2074.795 13.700 ;
        RECT 2090.555 13.685 2090.895 13.700 ;
        RECT 2096.305 13.685 2096.595 13.700 ;
        RECT 2105.735 13.685 2106.075 13.700 ;
        RECT 2124.365 13.685 2124.655 13.700 ;
        RECT 2125.515 13.685 2125.855 13.700 ;
        RECT 2136.095 13.685 2136.435 13.700 ;
        RECT 2137.475 13.685 2137.815 13.700 ;
        RECT 2141.615 13.685 2141.955 13.700 ;
        RECT 2152.425 13.685 2152.715 13.700 ;
        RECT 2174.735 13.685 2175.075 13.700 ;
        RECT 2179.795 13.685 2180.135 13.700 ;
        RECT 2180.485 13.685 2180.775 13.700 ;
        RECT 2190.375 13.685 2190.715 13.700 ;
        RECT 2192.675 13.685 2193.015 13.700 ;
        RECT 2208.545 13.685 2208.835 13.700 ;
        RECT 2234.535 13.685 2234.875 13.700 ;
        RECT 2236.605 13.685 2236.895 13.700 ;
        RECT 2239.135 13.685 2239.475 13.700 ;
        RECT 2241.435 13.685 2241.775 13.700 ;
        RECT 2264.665 13.685 2264.955 13.700 ;
        RECT 2272.255 13.685 2272.595 13.700 ;
        RECT 2277.315 13.685 2277.655 13.700 ;
        RECT 2292.725 13.685 2293.015 13.700 ;
        RECT 2297.095 13.685 2297.435 13.700 ;
        RECT 2320.785 13.685 2321.075 13.700 ;
        RECT 2321.935 13.685 2322.275 13.700 ;
        RECT 2348.845 13.685 2349.135 13.700 ;
        RECT 2376.905 13.685 2377.195 13.700 ;
        RECT 2404.965 13.685 2405.255 13.700 ;
        RECT 2428.195 13.685 2428.535 13.700 ;
        RECT 2433.025 13.685 2433.315 13.700 ;
        RECT 2440.155 13.685 2440.495 13.700 ;
        RECT 2461.085 13.685 2461.375 13.700 ;
        RECT 2489.145 13.685 2489.435 13.700 ;
        RECT 2490.755 13.685 2491.095 13.700 ;
        RECT 2496.735 13.685 2497.075 13.700 ;
        RECT 2498.115 13.685 2498.455 13.700 ;
        RECT 2500.875 13.685 2501.215 13.700 ;
        RECT 2502.255 13.685 2502.595 13.700 ;
        RECT 2510.075 13.685 2510.415 13.700 ;
        RECT 2517.205 13.685 2517.495 13.700 ;
        RECT 2525.715 13.685 2526.055 13.700 ;
        RECT 2530.775 13.685 2531.115 13.700 ;
        RECT 2534.455 13.685 2534.795 13.700 ;
        RECT 2545.265 13.685 2545.555 13.700 ;
        RECT 2548.255 13.685 2548.595 13.700 ;
        RECT 2551.935 13.685 2552.275 13.700 ;
        RECT 2554.695 13.685 2555.035 13.700 ;
        RECT 2569.875 13.685 2570.215 13.700 ;
        RECT 2573.325 13.685 2573.615 13.700 ;
        RECT 2581.375 13.685 2581.715 13.700 ;
        RECT 2586.435 13.685 2586.775 13.700 ;
        RECT 2593.335 13.685 2593.675 13.700 ;
        RECT 2598.395 13.685 2598.735 13.700 ;
        RECT 2601.385 13.685 2601.675 13.700 ;
        RECT 2609.895 13.685 2610.235 13.700 ;
        RECT 2629.445 13.685 2629.735 13.700 ;
        RECT 2655.895 13.685 2656.235 13.700 ;
        RECT 2657.505 13.685 2657.795 13.700 ;
        RECT 2685.565 13.685 2685.855 13.700 ;
        RECT 2686.715 13.685 2687.055 13.700 ;
        RECT 2689.015 13.685 2689.355 13.700 ;
        RECT 2713.625 13.685 2713.915 13.700 ;
        RECT 2726.275 13.685 2726.615 13.700 ;
        RECT 2727.655 13.685 2727.995 13.700 ;
        RECT 2730.875 13.685 2731.215 13.700 ;
        RECT 2741.685 13.685 2741.975 13.700 ;
        RECT 2769.745 13.685 2770.035 13.700 ;
        RECT 2797.805 13.685 2798.095 13.700 ;
        RECT 2825.865 13.685 2826.155 13.700 ;
        RECT 2853.925 13.685 2854.215 13.700 ;
        RECT 2855.995 13.685 2856.335 13.700 ;
        RECT 2881.985 13.685 2882.275 13.700 ;
        RECT 2907.975 13.685 2908.315 14.345 ;
        RECT 2909.355 13.685 2909.695 14.345 ;
        RECT 2910.045 13.685 2910.335 14.410 ;
        RECT 2911.195 13.685 2911.535 14.345 ;
        RECT 2912.805 13.685 2914.015 14.435 ;
        RECT 5.520 13.515 15.640 13.685 ;
        RECT 16.560 13.515 18.400 13.685 ;
        RECT 19.780 13.515 20.240 13.685 ;
        RECT 34.040 13.515 34.500 13.685 ;
        RECT 47.840 13.515 48.760 13.685 ;
        RECT 57.960 13.515 65.780 13.685 ;
        RECT 75.900 13.515 76.360 13.685 ;
        RECT 76.820 13.515 81.420 13.685 ;
        RECT 81.880 13.515 91.540 13.685 ;
        RECT 101.200 13.515 103.040 13.685 ;
        RECT 103.960 13.515 111.780 13.685 ;
        RECT 119.600 13.515 121.440 13.685 ;
        RECT 132.020 13.515 132.480 13.685 ;
        RECT 133.860 13.515 140.760 13.685 ;
        RECT 142.140 13.515 148.580 13.685 ;
        RECT 152.720 13.515 161.920 13.685 ;
        RECT 162.380 13.515 171.120 13.685 ;
        RECT 176.640 13.515 177.100 13.685 ;
        RECT 181.240 13.515 187.680 13.685 ;
        RECT 188.140 13.515 188.600 13.685 ;
        RECT 190.900 13.515 191.360 13.685 ;
        RECT 194.120 13.515 202.400 13.685 ;
        RECT 205.160 13.515 215.740 13.685 ;
        RECT 216.200 13.515 216.660 13.685 ;
        RECT 218.040 13.515 224.480 13.685 ;
        RECT 225.400 13.515 236.440 13.685 ;
        RECT 236.900 13.515 244.720 13.685 ;
        RECT 247.940 13.515 248.400 13.685 ;
        RECT 258.980 13.515 269.560 13.685 ;
        RECT 272.320 13.515 272.780 13.685 ;
        RECT 276.460 13.515 276.920 13.685 ;
        RECT 277.380 13.515 278.760 13.685 ;
        RECT 282.900 13.515 284.740 13.685 ;
        RECT 288.880 13.515 290.260 13.685 ;
        RECT 290.720 13.515 291.180 13.685 ;
        RECT 292.560 13.515 299.000 13.685 ;
        RECT 300.380 13.515 300.840 13.685 ;
        RECT 304.520 13.515 307.280 13.685 ;
        RECT 307.740 13.515 311.420 13.685 ;
        RECT 314.180 13.515 315.560 13.685 ;
        RECT 317.400 13.515 326.140 13.685 ;
        RECT 328.440 13.515 337.640 13.685 ;
        RECT 339.020 13.515 340.860 13.685 ;
        RECT 347.760 13.515 358.800 13.685 ;
        RECT 359.720 13.515 367.080 13.685 ;
        RECT 368.000 13.515 375.360 13.685 ;
        RECT 376.280 13.515 376.740 13.685 ;
        RECT 384.560 13.515 404.340 13.685 ;
        RECT 404.800 13.515 405.260 13.685 ;
        RECT 412.620 13.515 413.080 13.685 ;
        RECT 413.540 13.515 420.900 13.685 ;
        RECT 425.500 13.515 434.240 13.685 ;
        RECT 440.680 13.515 441.140 13.685 ;
        RECT 445.280 13.515 457.240 13.685 ;
        RECT 457.700 13.515 466.440 13.685 ;
        RECT 466.900 13.515 469.200 13.685 ;
        RECT 476.100 13.515 476.560 13.685 ;
        RECT 480.700 13.515 482.540 13.685 ;
        RECT 490.360 13.515 490.820 13.685 ;
        RECT 494.500 13.515 495.880 13.685 ;
        RECT 496.800 13.515 497.260 13.685 ;
        RECT 504.620 13.515 505.080 13.685 ;
        RECT 518.880 13.515 519.340 13.685 ;
        RECT 524.860 13.515 525.320 13.685 ;
        RECT 527.620 13.515 534.060 13.685 ;
        RECT 535.900 13.515 537.280 13.685 ;
        RECT 538.660 13.515 540.500 13.685 ;
        RECT 547.400 13.515 547.860 13.685 ;
        RECT 552.920 13.515 553.380 13.685 ;
        RECT 561.660 13.515 562.120 13.685 ;
        RECT 563.960 13.515 565.800 13.685 ;
        RECT 570.860 13.515 580.520 13.685 ;
        RECT 580.980 13.515 581.440 13.685 ;
        RECT 590.180 13.515 590.640 13.685 ;
        RECT 604.440 13.515 604.900 13.685 ;
        RECT 609.040 13.515 609.500 13.685 ;
        RECT 618.700 13.515 619.160 13.685 ;
        RECT 632.960 13.515 633.420 13.685 ;
        RECT 637.100 13.515 637.560 13.685 ;
        RECT 647.220 13.515 647.680 13.685 ;
        RECT 661.480 13.515 661.940 13.685 ;
        RECT 665.160 13.515 665.620 13.685 ;
        RECT 675.740 13.515 676.200 13.685 ;
        RECT 690.000 13.515 690.460 13.685 ;
        RECT 693.220 13.515 693.680 13.685 ;
        RECT 704.260 13.515 704.720 13.685 ;
        RECT 718.520 13.515 718.980 13.685 ;
        RECT 721.280 13.515 721.740 13.685 ;
        RECT 732.780 13.515 733.240 13.685 ;
        RECT 747.040 13.515 747.500 13.685 ;
        RECT 749.340 13.515 749.800 13.685 ;
        RECT 761.300 13.515 761.760 13.685 ;
        RECT 775.560 13.515 776.020 13.685 ;
        RECT 777.400 13.515 777.860 13.685 ;
        RECT 789.820 13.515 790.280 13.685 ;
        RECT 804.080 13.515 804.540 13.685 ;
        RECT 805.460 13.515 805.920 13.685 ;
        RECT 818.340 13.515 818.800 13.685 ;
        RECT 832.600 13.515 833.060 13.685 ;
        RECT 833.520 13.515 833.980 13.685 ;
        RECT 846.860 13.515 847.320 13.685 ;
        RECT 861.120 13.515 862.040 13.685 ;
        RECT 875.380 13.515 875.840 13.685 ;
        RECT 889.640 13.515 890.100 13.685 ;
        RECT 903.900 13.515 904.360 13.685 ;
        RECT 917.700 13.515 918.620 13.685 ;
        RECT 932.420 13.515 932.880 13.685 ;
        RECT 945.760 13.515 946.220 13.685 ;
        RECT 946.680 13.515 947.140 13.685 ;
        RECT 960.940 13.515 961.400 13.685 ;
        RECT 973.820 13.515 974.280 13.685 ;
        RECT 975.200 13.515 975.660 13.685 ;
        RECT 989.460 13.515 989.920 13.685 ;
        RECT 1001.880 13.515 1002.340 13.685 ;
        RECT 1003.720 13.515 1004.180 13.685 ;
        RECT 1017.980 13.515 1018.440 13.685 ;
        RECT 1029.940 13.515 1030.400 13.685 ;
        RECT 1032.240 13.515 1032.700 13.685 ;
        RECT 1046.500 13.515 1046.960 13.685 ;
        RECT 1058.000 13.515 1058.460 13.685 ;
        RECT 1060.760 13.515 1061.220 13.685 ;
        RECT 1075.020 13.515 1075.480 13.685 ;
        RECT 1086.060 13.515 1086.520 13.685 ;
        RECT 1089.280 13.515 1089.740 13.685 ;
        RECT 1103.540 13.515 1104.000 13.685 ;
        RECT 1114.120 13.515 1114.580 13.685 ;
        RECT 1117.800 13.515 1118.260 13.685 ;
        RECT 1132.060 13.515 1132.520 13.685 ;
        RECT 1142.180 13.515 1142.640 13.685 ;
        RECT 1146.320 13.515 1146.780 13.685 ;
        RECT 1160.580 13.515 1161.040 13.685 ;
        RECT 1170.240 13.515 1170.700 13.685 ;
        RECT 1174.840 13.515 1175.300 13.685 ;
        RECT 1189.100 13.515 1189.560 13.685 ;
        RECT 1198.300 13.515 1198.760 13.685 ;
        RECT 1203.360 13.515 1203.820 13.685 ;
        RECT 1217.620 13.515 1218.080 13.685 ;
        RECT 1226.360 13.515 1226.820 13.685 ;
        RECT 1231.880 13.515 1232.340 13.685 ;
        RECT 1246.140 13.515 1246.600 13.685 ;
        RECT 1254.420 13.515 1254.880 13.685 ;
        RECT 1260.400 13.515 1260.860 13.685 ;
        RECT 1274.660 13.515 1275.120 13.685 ;
        RECT 1282.480 13.515 1282.940 13.685 ;
        RECT 1288.920 13.515 1289.380 13.685 ;
        RECT 1303.180 13.515 1303.640 13.685 ;
        RECT 1310.540 13.515 1311.000 13.685 ;
        RECT 1317.440 13.515 1317.900 13.685 ;
        RECT 1331.700 13.515 1332.160 13.685 ;
        RECT 1338.600 13.515 1339.060 13.685 ;
        RECT 1345.960 13.515 1346.420 13.685 ;
        RECT 1360.220 13.515 1360.680 13.685 ;
        RECT 1366.660 13.515 1367.120 13.685 ;
        RECT 1374.480 13.515 1374.940 13.685 ;
        RECT 1382.300 13.515 1383.680 13.685 ;
        RECT 1388.740 13.515 1389.200 13.685 ;
        RECT 1394.720 13.515 1395.180 13.685 ;
        RECT 1400.700 13.515 1402.080 13.685 ;
        RECT 1403.000 13.515 1403.460 13.685 ;
        RECT 1417.260 13.515 1417.720 13.685 ;
        RECT 1422.780 13.515 1423.240 13.685 ;
        RECT 1431.520 13.515 1431.980 13.685 ;
        RECT 1445.780 13.515 1446.240 13.685 ;
        RECT 1450.840 13.515 1451.300 13.685 ;
        RECT 1460.040 13.515 1460.500 13.685 ;
        RECT 1474.300 13.515 1474.760 13.685 ;
        RECT 1478.900 13.515 1479.360 13.685 ;
        RECT 1488.560 13.515 1489.020 13.685 ;
        RECT 1502.820 13.515 1503.280 13.685 ;
        RECT 1503.740 13.515 1505.120 13.685 ;
        RECT 1506.960 13.515 1507.420 13.685 ;
        RECT 1517.080 13.515 1517.540 13.685 ;
        RECT 1525.820 13.515 1527.200 13.685 ;
        RECT 1531.340 13.515 1531.800 13.685 ;
        RECT 1535.020 13.515 1536.860 13.685 ;
        RECT 1539.160 13.515 1540.540 13.685 ;
        RECT 1542.380 13.515 1543.760 13.685 ;
        RECT 1545.600 13.515 1546.060 13.685 ;
        RECT 1558.940 13.515 1560.320 13.685 ;
        RECT 1563.080 13.515 1563.540 13.685 ;
        RECT 1574.120 13.515 1574.580 13.685 ;
        RECT 1575.500 13.515 1576.880 13.685 ;
        RECT 1588.380 13.515 1589.760 13.685 ;
        RECT 1591.140 13.515 1591.600 13.685 ;
        RECT 1602.640 13.515 1603.100 13.685 ;
        RECT 1616.900 13.515 1617.360 13.685 ;
        RECT 1619.200 13.515 1619.660 13.685 ;
        RECT 1625.640 13.515 1627.020 13.685 ;
        RECT 1631.160 13.515 1631.620 13.685 ;
        RECT 1645.420 13.515 1645.880 13.685 ;
        RECT 1647.260 13.515 1647.720 13.685 ;
        RECT 1648.640 13.515 1650.020 13.685 ;
        RECT 1659.680 13.515 1660.140 13.685 ;
        RECT 1673.940 13.515 1674.400 13.685 ;
        RECT 1675.320 13.515 1675.780 13.685 ;
        RECT 1688.200 13.515 1688.660 13.685 ;
        RECT 1702.460 13.515 1702.920 13.685 ;
        RECT 1703.380 13.515 1703.840 13.685 ;
        RECT 1716.720 13.515 1717.180 13.685 ;
        RECT 1730.980 13.515 1731.900 13.685 ;
        RECT 1745.240 13.515 1745.700 13.685 ;
        RECT 1759.500 13.515 1761.340 13.685 ;
        RECT 1773.760 13.515 1775.140 13.685 ;
        RECT 1787.560 13.515 1788.480 13.685 ;
        RECT 1802.280 13.515 1802.740 13.685 ;
        RECT 1815.620 13.515 1816.080 13.685 ;
        RECT 1816.540 13.515 1817.000 13.685 ;
        RECT 1829.880 13.515 1831.260 13.685 ;
        RECT 1843.680 13.515 1844.140 13.685 ;
        RECT 1845.060 13.515 1845.520 13.685 ;
        RECT 1859.320 13.515 1859.780 13.685 ;
        RECT 1871.740 13.515 1872.200 13.685 ;
        RECT 1873.580 13.515 1874.040 13.685 ;
        RECT 1887.840 13.515 1888.300 13.685 ;
        RECT 1899.800 13.515 1900.260 13.685 ;
        RECT 1902.100 13.515 1902.560 13.685 ;
        RECT 1913.140 13.515 1914.520 13.685 ;
        RECT 1916.360 13.515 1916.820 13.685 ;
        RECT 1925.560 13.515 1926.940 13.685 ;
        RECT 1927.860 13.515 1928.320 13.685 ;
        RECT 1930.620 13.515 1931.080 13.685 ;
        RECT 1931.540 13.515 1932.920 13.685 ;
        RECT 1944.880 13.515 1945.340 13.685 ;
        RECT 1947.640 13.515 1949.020 13.685 ;
        RECT 1955.920 13.515 1956.380 13.685 ;
        RECT 1959.140 13.515 1959.600 13.685 ;
        RECT 1972.940 13.515 1974.320 13.685 ;
        RECT 1982.600 13.515 1984.440 13.685 ;
        RECT 1987.660 13.515 1988.120 13.685 ;
        RECT 1991.800 13.515 1993.180 13.685 ;
        RECT 1995.020 13.515 1996.400 13.685 ;
        RECT 1999.620 13.515 2001.000 13.685 ;
        RECT 2001.920 13.515 2002.380 13.685 ;
        RECT 2012.040 13.515 2012.500 13.685 ;
        RECT 2016.180 13.515 2016.640 13.685 ;
        RECT 2018.020 13.515 2019.400 13.685 ;
        RECT 2024.460 13.515 2025.840 13.685 ;
        RECT 2030.440 13.515 2030.900 13.685 ;
        RECT 2037.340 13.515 2038.720 13.685 ;
        RECT 2040.100 13.515 2040.560 13.685 ;
        RECT 2044.700 13.515 2045.160 13.685 ;
        RECT 2058.960 13.515 2061.720 13.685 ;
        RECT 2068.160 13.515 2068.620 13.685 ;
        RECT 2073.220 13.515 2075.060 13.685 ;
        RECT 2087.480 13.515 2087.940 13.685 ;
        RECT 2089.780 13.515 2091.160 13.685 ;
        RECT 2096.220 13.515 2096.680 13.685 ;
        RECT 2101.740 13.515 2102.200 13.685 ;
        RECT 2104.960 13.515 2106.340 13.685 ;
        RECT 2116.000 13.515 2116.460 13.685 ;
        RECT 2124.280 13.515 2126.120 13.685 ;
        RECT 2130.260 13.515 2130.720 13.685 ;
        RECT 2135.320 13.515 2138.080 13.685 ;
        RECT 2140.840 13.515 2142.220 13.685 ;
        RECT 2144.520 13.515 2144.980 13.685 ;
        RECT 2152.340 13.515 2152.800 13.685 ;
        RECT 2158.780 13.515 2159.240 13.685 ;
        RECT 2173.040 13.515 2173.500 13.685 ;
        RECT 2173.960 13.515 2175.340 13.685 ;
        RECT 2179.020 13.515 2180.860 13.685 ;
        RECT 2187.300 13.515 2187.760 13.685 ;
        RECT 2189.600 13.515 2190.980 13.685 ;
        RECT 2191.900 13.515 2193.280 13.685 ;
        RECT 2201.560 13.515 2202.020 13.685 ;
        RECT 2208.460 13.515 2208.920 13.685 ;
        RECT 2215.820 13.515 2216.280 13.685 ;
        RECT 2230.080 13.515 2230.540 13.685 ;
        RECT 2233.760 13.515 2235.140 13.685 ;
        RECT 2236.520 13.515 2236.980 13.685 ;
        RECT 2238.360 13.515 2239.740 13.685 ;
        RECT 2240.660 13.515 2242.040 13.685 ;
        RECT 2244.340 13.515 2244.800 13.685 ;
        RECT 2258.600 13.515 2259.060 13.685 ;
        RECT 2264.580 13.515 2265.040 13.685 ;
        RECT 2271.480 13.515 2273.320 13.685 ;
        RECT 2276.540 13.515 2277.920 13.685 ;
        RECT 2287.120 13.515 2287.580 13.685 ;
        RECT 2292.640 13.515 2293.100 13.685 ;
        RECT 2296.320 13.515 2297.700 13.685 ;
        RECT 2301.380 13.515 2301.840 13.685 ;
        RECT 2315.640 13.515 2316.100 13.685 ;
        RECT 2320.700 13.515 2322.540 13.685 ;
        RECT 2329.900 13.515 2330.360 13.685 ;
        RECT 2344.160 13.515 2344.620 13.685 ;
        RECT 2348.760 13.515 2349.220 13.685 ;
        RECT 2358.420 13.515 2358.880 13.685 ;
        RECT 2372.680 13.515 2373.140 13.685 ;
        RECT 2376.820 13.515 2377.280 13.685 ;
        RECT 2386.940 13.515 2387.400 13.685 ;
        RECT 2401.200 13.515 2401.660 13.685 ;
        RECT 2404.880 13.515 2405.340 13.685 ;
        RECT 2415.460 13.515 2415.920 13.685 ;
        RECT 2427.420 13.515 2428.800 13.685 ;
        RECT 2429.720 13.515 2430.180 13.685 ;
        RECT 2432.940 13.515 2433.400 13.685 ;
        RECT 2439.380 13.515 2440.760 13.685 ;
        RECT 2443.980 13.515 2444.440 13.685 ;
        RECT 2458.240 13.515 2458.700 13.685 ;
        RECT 2461.000 13.515 2461.460 13.685 ;
        RECT 2472.500 13.515 2472.960 13.685 ;
        RECT 2486.760 13.515 2487.220 13.685 ;
        RECT 2489.060 13.515 2489.520 13.685 ;
        RECT 2489.980 13.515 2491.360 13.685 ;
        RECT 2495.960 13.515 2498.720 13.685 ;
        RECT 2500.100 13.515 2502.860 13.685 ;
        RECT 2509.300 13.515 2510.680 13.685 ;
        RECT 2515.280 13.515 2515.740 13.685 ;
        RECT 2517.120 13.515 2517.580 13.685 ;
        RECT 2524.940 13.515 2526.320 13.685 ;
        RECT 2529.540 13.515 2531.380 13.685 ;
        RECT 2533.680 13.515 2535.060 13.685 ;
        RECT 2543.800 13.515 2544.260 13.685 ;
        RECT 2545.180 13.515 2545.640 13.685 ;
        RECT 2547.480 13.515 2548.860 13.685 ;
        RECT 2551.160 13.515 2552.540 13.685 ;
        RECT 2553.920 13.515 2555.300 13.685 ;
        RECT 2558.060 13.515 2558.520 13.685 ;
        RECT 2569.100 13.515 2570.480 13.685 ;
        RECT 2572.320 13.515 2572.780 13.685 ;
        RECT 2573.240 13.515 2573.700 13.685 ;
        RECT 2580.600 13.515 2581.980 13.685 ;
        RECT 2585.660 13.515 2587.040 13.685 ;
        RECT 2592.560 13.515 2593.940 13.685 ;
        RECT 2597.620 13.515 2599.000 13.685 ;
        RECT 2600.840 13.515 2601.760 13.685 ;
        RECT 2609.120 13.515 2610.500 13.685 ;
        RECT 2615.100 13.515 2615.560 13.685 ;
        RECT 2629.360 13.515 2629.820 13.685 ;
        RECT 2643.620 13.515 2644.080 13.685 ;
        RECT 2655.120 13.515 2656.500 13.685 ;
        RECT 2657.420 13.515 2658.340 13.685 ;
        RECT 2672.140 13.515 2672.600 13.685 ;
        RECT 2685.480 13.515 2687.320 13.685 ;
        RECT 2688.240 13.515 2689.620 13.685 ;
        RECT 2700.660 13.515 2701.120 13.685 ;
        RECT 2713.540 13.515 2714.000 13.685 ;
        RECT 2714.920 13.515 2715.380 13.685 ;
        RECT 2725.500 13.515 2728.260 13.685 ;
        RECT 2729.180 13.515 2729.640 13.685 ;
        RECT 2730.100 13.515 2731.480 13.685 ;
        RECT 2741.600 13.515 2742.060 13.685 ;
        RECT 2743.440 13.515 2743.900 13.685 ;
        RECT 2757.700 13.515 2758.160 13.685 ;
        RECT 2769.660 13.515 2770.120 13.685 ;
        RECT 2771.960 13.515 2772.420 13.685 ;
        RECT 2786.220 13.515 2786.680 13.685 ;
        RECT 2797.720 13.515 2798.180 13.685 ;
        RECT 2800.480 13.515 2800.940 13.685 ;
        RECT 2814.740 13.515 2815.200 13.685 ;
        RECT 2825.780 13.515 2826.240 13.685 ;
        RECT 2829.000 13.515 2829.460 13.685 ;
        RECT 2843.260 13.515 2843.720 13.685 ;
        RECT 2853.840 13.515 2854.300 13.685 ;
        RECT 2855.220 13.515 2856.600 13.685 ;
        RECT 2857.520 13.515 2857.980 13.685 ;
        RECT 2871.780 13.515 2872.240 13.685 ;
        RECT 2881.900 13.515 2882.360 13.685 ;
        RECT 2886.040 13.515 2886.500 13.685 ;
        RECT 2900.300 13.515 2900.760 13.685 ;
        RECT 2907.200 13.515 2911.800 13.685 ;
        RECT 2912.720 13.515 2914.100 13.685 ;
        RECT 5.605 12.765 6.815 13.515 ;
        RECT 5.605 12.225 6.125 12.765 ;
        RECT 8.865 12.695 9.095 13.515 ;
        RECT 9.765 12.695 9.975 13.515 ;
        RECT 10.895 12.855 11.235 13.515 ;
        RECT 19.865 12.790 20.155 13.515 ;
        RECT 34.125 12.790 34.415 13.515 ;
        RECT 48.385 12.790 48.675 13.515 ;
        RECT 62.645 12.790 62.935 13.515 ;
        RECT 76.905 12.790 77.195 13.515 ;
        RECT 82.395 13.135 82.725 13.515 ;
        RECT 83.335 13.055 83.585 13.515 ;
        RECT 85.280 13.015 85.650 13.515 ;
        RECT 87.505 12.985 87.675 13.515 ;
        RECT 88.505 13.035 88.675 13.515 ;
        RECT 89.375 13.040 89.545 13.515 ;
        RECT 90.225 13.040 90.395 13.515 ;
        RECT 91.165 12.790 91.455 13.515 ;
        RECT 105.425 12.790 105.715 13.515 ;
        RECT 119.685 12.790 119.975 13.515 ;
        RECT 133.945 12.790 134.235 13.515 ;
        RECT 148.205 12.790 148.495 13.515 ;
        RECT 162.465 12.790 162.755 13.515 ;
        RECT 176.725 12.790 177.015 13.515 ;
        RECT 190.985 12.790 191.275 13.515 ;
        RECT 205.245 12.790 205.535 13.515 ;
        RECT 205.795 12.705 205.965 13.515 ;
        RECT 207.475 13.045 207.645 13.515 ;
        RECT 208.315 13.045 209.005 13.515 ;
        RECT 209.675 13.045 209.845 13.515 ;
        RECT 210.515 12.705 210.685 13.515 ;
        RECT 211.355 13.045 211.525 13.515 ;
        RECT 212.195 13.045 212.365 13.515 ;
        RECT 219.505 12.790 219.795 13.515 ;
        RECT 225.660 13.045 225.830 13.515 ;
        RECT 226.500 13.045 226.670 13.515 ;
        RECT 227.340 13.045 227.510 13.515 ;
        RECT 230.040 13.045 230.210 13.515 ;
        RECT 230.880 13.045 231.050 13.515 ;
        RECT 233.765 12.790 234.055 13.515 ;
        RECT 242.025 13.155 242.355 13.515 ;
        RECT 242.930 13.155 243.260 13.515 ;
        RECT 243.790 13.155 244.120 13.515 ;
        RECT 248.025 12.790 248.315 13.515 ;
        RECT 262.285 12.790 262.575 13.515 ;
        RECT 262.920 13.045 263.090 13.515 ;
        RECT 263.760 13.045 263.930 13.515 ;
        RECT 264.600 13.045 264.770 13.515 ;
        RECT 267.300 13.045 267.470 13.515 ;
        RECT 268.140 13.045 268.310 13.515 ;
        RECT 276.545 12.790 276.835 13.515 ;
        RECT 290.805 12.790 291.095 13.515 ;
        RECT 305.065 12.790 305.355 13.515 ;
        RECT 319.325 12.790 319.615 13.515 ;
        RECT 333.585 12.790 333.875 13.515 ;
        RECT 347.845 12.790 348.135 13.515 ;
        RECT 352.485 12.695 352.715 13.515 ;
        RECT 353.385 12.695 353.595 13.515 ;
        RECT 362.105 12.790 362.395 13.515 ;
        RECT 376.365 12.790 376.655 13.515 ;
        RECT 390.625 12.790 390.915 13.515 ;
        RECT 391.515 13.135 391.845 13.515 ;
        RECT 392.455 13.055 392.705 13.515 ;
        RECT 394.400 13.015 394.770 13.515 ;
        RECT 396.625 12.985 396.795 13.515 ;
        RECT 397.625 13.035 397.795 13.515 ;
        RECT 398.495 13.040 398.665 13.515 ;
        RECT 399.345 13.040 399.515 13.515 ;
        RECT 399.865 12.695 400.095 13.515 ;
        RECT 400.765 12.695 400.975 13.515 ;
        RECT 404.885 12.790 405.175 13.515 ;
        RECT 419.145 12.790 419.435 13.515 ;
        RECT 433.405 12.790 433.695 13.515 ;
        RECT 447.665 12.790 447.955 13.515 ;
        RECT 451.060 13.045 451.230 13.515 ;
        RECT 451.900 13.045 452.070 13.515 ;
        RECT 452.740 13.045 452.910 13.515 ;
        RECT 455.440 13.045 455.610 13.515 ;
        RECT 456.280 13.045 456.450 13.515 ;
        RECT 461.925 12.790 462.215 13.515 ;
        RECT 476.185 12.790 476.475 13.515 ;
        RECT 490.445 12.790 490.735 13.515 ;
        RECT 504.705 12.790 504.995 13.515 ;
        RECT 518.965 12.790 519.255 13.515 ;
        RECT 533.225 12.790 533.515 13.515 ;
        RECT 547.485 12.790 547.775 13.515 ;
        RECT 561.745 12.790 562.035 13.515 ;
        RECT 576.005 12.790 576.295 13.515 ;
        RECT 590.265 12.790 590.555 13.515 ;
        RECT 604.525 12.790 604.815 13.515 ;
        RECT 618.785 12.790 619.075 13.515 ;
        RECT 633.045 12.790 633.335 13.515 ;
        RECT 647.305 12.790 647.595 13.515 ;
        RECT 661.565 12.790 661.855 13.515 ;
        RECT 675.825 12.790 676.115 13.515 ;
        RECT 690.085 12.790 690.375 13.515 ;
        RECT 704.345 12.790 704.635 13.515 ;
        RECT 718.605 12.790 718.895 13.515 ;
        RECT 732.865 12.790 733.155 13.515 ;
        RECT 747.125 12.790 747.415 13.515 ;
        RECT 761.385 12.790 761.675 13.515 ;
        RECT 775.645 12.790 775.935 13.515 ;
        RECT 789.905 12.790 790.195 13.515 ;
        RECT 804.165 12.790 804.455 13.515 ;
        RECT 818.425 12.790 818.715 13.515 ;
        RECT 832.685 12.790 832.975 13.515 ;
        RECT 846.945 12.790 847.235 13.515 ;
        RECT 861.205 12.790 861.495 13.515 ;
        RECT 875.465 12.790 875.755 13.515 ;
        RECT 889.725 12.790 890.015 13.515 ;
        RECT 903.985 12.790 904.275 13.515 ;
        RECT 918.245 12.790 918.535 13.515 ;
        RECT 932.505 12.790 932.795 13.515 ;
        RECT 946.765 12.790 947.055 13.515 ;
        RECT 961.025 12.790 961.315 13.515 ;
        RECT 975.285 12.790 975.575 13.515 ;
        RECT 989.545 12.790 989.835 13.515 ;
        RECT 1003.805 12.790 1004.095 13.515 ;
        RECT 1018.065 12.790 1018.355 13.515 ;
        RECT 1032.325 12.790 1032.615 13.515 ;
        RECT 1046.585 12.790 1046.875 13.515 ;
        RECT 1060.845 12.790 1061.135 13.515 ;
        RECT 1075.105 12.790 1075.395 13.515 ;
        RECT 1089.365 12.790 1089.655 13.515 ;
        RECT 1103.625 12.790 1103.915 13.515 ;
        RECT 1117.885 12.790 1118.175 13.515 ;
        RECT 1132.145 12.790 1132.435 13.515 ;
        RECT 1146.405 12.790 1146.695 13.515 ;
        RECT 1160.665 12.790 1160.955 13.515 ;
        RECT 1174.925 12.790 1175.215 13.515 ;
        RECT 1189.185 12.790 1189.475 13.515 ;
        RECT 1203.445 12.790 1203.735 13.515 ;
        RECT 1217.705 12.790 1217.995 13.515 ;
        RECT 1231.965 12.790 1232.255 13.515 ;
        RECT 1246.225 12.790 1246.515 13.515 ;
        RECT 1260.485 12.790 1260.775 13.515 ;
        RECT 1274.745 12.790 1275.035 13.515 ;
        RECT 1289.005 12.790 1289.295 13.515 ;
        RECT 1303.265 12.790 1303.555 13.515 ;
        RECT 1317.525 12.790 1317.815 13.515 ;
        RECT 1331.785 12.790 1332.075 13.515 ;
        RECT 1346.045 12.790 1346.335 13.515 ;
        RECT 1360.305 12.790 1360.595 13.515 ;
        RECT 1374.565 12.790 1374.855 13.515 ;
        RECT 1388.825 12.790 1389.115 13.515 ;
        RECT 1403.085 12.790 1403.375 13.515 ;
        RECT 1417.345 12.790 1417.635 13.515 ;
        RECT 1431.605 12.790 1431.895 13.515 ;
        RECT 1445.865 12.790 1446.155 13.515 ;
        RECT 1460.125 12.790 1460.415 13.515 ;
        RECT 1474.385 12.790 1474.675 13.515 ;
        RECT 1488.645 12.790 1488.935 13.515 ;
        RECT 1502.905 12.790 1503.195 13.515 ;
        RECT 1517.165 12.790 1517.455 13.515 ;
        RECT 1531.425 12.790 1531.715 13.515 ;
        RECT 1545.685 12.790 1545.975 13.515 ;
        RECT 1559.945 12.790 1560.235 13.515 ;
        RECT 1574.205 12.790 1574.495 13.515 ;
        RECT 1588.465 12.790 1588.755 13.515 ;
        RECT 1602.725 12.790 1603.015 13.515 ;
        RECT 1616.985 12.790 1617.275 13.515 ;
        RECT 1631.245 12.790 1631.535 13.515 ;
        RECT 1645.505 12.790 1645.795 13.515 ;
        RECT 1659.765 12.790 1660.055 13.515 ;
        RECT 1674.025 12.790 1674.315 13.515 ;
        RECT 1688.285 12.790 1688.575 13.515 ;
        RECT 1702.545 12.790 1702.835 13.515 ;
        RECT 1716.805 12.790 1717.095 13.515 ;
        RECT 1731.065 12.790 1731.355 13.515 ;
        RECT 1745.325 12.790 1745.615 13.515 ;
        RECT 1759.585 12.790 1759.875 13.515 ;
        RECT 1773.845 12.790 1774.135 13.515 ;
        RECT 1788.105 12.790 1788.395 13.515 ;
        RECT 1802.365 12.790 1802.655 13.515 ;
        RECT 1816.625 12.790 1816.915 13.515 ;
        RECT 1830.885 12.790 1831.175 13.515 ;
        RECT 1845.145 12.790 1845.435 13.515 ;
        RECT 1859.405 12.790 1859.695 13.515 ;
        RECT 1873.665 12.790 1873.955 13.515 ;
        RECT 1887.925 12.790 1888.215 13.515 ;
        RECT 1902.185 12.790 1902.475 13.515 ;
        RECT 1916.445 12.790 1916.735 13.515 ;
        RECT 1930.705 12.790 1930.995 13.515 ;
        RECT 1944.965 12.790 1945.255 13.515 ;
        RECT 1959.225 12.790 1959.515 13.515 ;
        RECT 1973.485 12.790 1973.775 13.515 ;
        RECT 1987.745 12.790 1988.035 13.515 ;
        RECT 2002.005 12.790 2002.295 13.515 ;
        RECT 2016.265 12.790 2016.555 13.515 ;
        RECT 2030.525 12.790 2030.815 13.515 ;
        RECT 2044.785 12.790 2045.075 13.515 ;
        RECT 2059.045 12.790 2059.335 13.515 ;
        RECT 2073.305 12.790 2073.595 13.515 ;
        RECT 2087.565 12.790 2087.855 13.515 ;
        RECT 2101.825 12.790 2102.115 13.515 ;
        RECT 2116.085 12.790 2116.375 13.515 ;
        RECT 2130.345 12.790 2130.635 13.515 ;
        RECT 2144.605 12.790 2144.895 13.515 ;
        RECT 2158.865 12.790 2159.155 13.515 ;
        RECT 2173.125 12.790 2173.415 13.515 ;
        RECT 2187.385 12.790 2187.675 13.515 ;
        RECT 2201.645 12.790 2201.935 13.515 ;
        RECT 2215.905 12.790 2216.195 13.515 ;
        RECT 2230.165 12.790 2230.455 13.515 ;
        RECT 2244.425 12.790 2244.715 13.515 ;
        RECT 2258.685 12.790 2258.975 13.515 ;
        RECT 2272.945 12.790 2273.235 13.515 ;
        RECT 2287.205 12.790 2287.495 13.515 ;
        RECT 2301.465 12.790 2301.755 13.515 ;
        RECT 2315.725 12.790 2316.015 13.515 ;
        RECT 2329.985 12.790 2330.275 13.515 ;
        RECT 2344.245 12.790 2344.535 13.515 ;
        RECT 2358.505 12.790 2358.795 13.515 ;
        RECT 2372.765 12.790 2373.055 13.515 ;
        RECT 2387.025 12.790 2387.315 13.515 ;
        RECT 2401.285 12.790 2401.575 13.515 ;
        RECT 2415.545 12.790 2415.835 13.515 ;
        RECT 2429.805 12.790 2430.095 13.515 ;
        RECT 2444.065 12.790 2444.355 13.515 ;
        RECT 2458.325 12.790 2458.615 13.515 ;
        RECT 2472.585 12.790 2472.875 13.515 ;
        RECT 2486.845 12.790 2487.135 13.515 ;
        RECT 2501.105 12.790 2501.395 13.515 ;
        RECT 2515.365 12.790 2515.655 13.515 ;
        RECT 2529.625 12.790 2529.915 13.515 ;
        RECT 2543.885 12.790 2544.175 13.515 ;
        RECT 2558.145 12.790 2558.435 13.515 ;
        RECT 2572.405 12.790 2572.695 13.515 ;
        RECT 2586.665 12.790 2586.955 13.515 ;
        RECT 2600.925 12.790 2601.215 13.515 ;
        RECT 2615.185 12.790 2615.475 13.515 ;
        RECT 2629.445 12.790 2629.735 13.515 ;
        RECT 2643.705 12.790 2643.995 13.515 ;
        RECT 2657.965 12.790 2658.255 13.515 ;
        RECT 2672.225 12.790 2672.515 13.515 ;
        RECT 2686.485 12.790 2686.775 13.515 ;
        RECT 2700.745 12.790 2701.035 13.515 ;
        RECT 2715.005 12.790 2715.295 13.515 ;
        RECT 2729.265 12.790 2729.555 13.515 ;
        RECT 2743.525 12.790 2743.815 13.515 ;
        RECT 2757.785 12.790 2758.075 13.515 ;
        RECT 2772.045 12.790 2772.335 13.515 ;
        RECT 2786.305 12.790 2786.595 13.515 ;
        RECT 2800.565 12.790 2800.855 13.515 ;
        RECT 2814.825 12.790 2815.115 13.515 ;
        RECT 2829.085 12.790 2829.375 13.515 ;
        RECT 2843.345 12.790 2843.635 13.515 ;
        RECT 2857.605 12.790 2857.895 13.515 ;
        RECT 2871.865 12.790 2872.155 13.515 ;
        RECT 2886.125 12.790 2886.415 13.515 ;
        RECT 2900.385 12.790 2900.675 13.515 ;
        RECT 2909.815 12.855 2910.155 13.515 ;
        RECT 2912.805 12.765 2914.015 13.515 ;
        RECT 2913.495 12.225 2914.015 12.765 ;
      LAYER mcon ;
        RECT 5.665 3505.995 5.835 3506.165 ;
        RECT 6.125 3505.995 6.295 3506.165 ;
        RECT 6.585 3505.995 6.755 3506.165 ;
        RECT 9.805 3505.995 9.975 3506.165 ;
        RECT 10.265 3505.995 10.435 3506.165 ;
        RECT 10.725 3505.995 10.895 3506.165 ;
        RECT 11.185 3505.995 11.355 3506.165 ;
        RECT 11.645 3505.995 11.815 3506.165 ;
        RECT 12.105 3505.995 12.275 3506.165 ;
        RECT 2909.185 3505.995 2909.355 3506.165 ;
        RECT 2909.645 3505.995 2909.815 3506.165 ;
        RECT 2910.105 3505.995 2910.275 3506.165 ;
        RECT 2910.565 3505.995 2910.735 3506.165 ;
        RECT 2911.025 3505.995 2911.195 3506.165 ;
        RECT 2911.485 3505.995 2911.655 3506.165 ;
        RECT 2912.865 3505.995 2913.035 3506.165 ;
        RECT 2913.325 3505.995 2913.495 3506.165 ;
        RECT 2913.785 3505.995 2913.955 3506.165 ;
        RECT 5.665 3500.555 5.835 3500.725 ;
        RECT 6.125 3500.555 6.295 3500.725 ;
        RECT 6.585 3500.555 6.755 3500.725 ;
        RECT 2910.105 3500.555 2910.275 3500.725 ;
        RECT 2912.865 3500.555 2913.035 3500.725 ;
        RECT 2913.325 3500.555 2913.495 3500.725 ;
        RECT 2913.785 3500.555 2913.955 3500.725 ;
        RECT 5.665 3495.115 5.835 3495.285 ;
        RECT 6.125 3495.115 6.295 3495.285 ;
        RECT 6.585 3495.115 6.755 3495.285 ;
        RECT 2910.105 3495.115 2910.275 3495.285 ;
        RECT 2912.865 3495.115 2913.035 3495.285 ;
        RECT 2913.325 3495.115 2913.495 3495.285 ;
        RECT 2913.785 3495.115 2913.955 3495.285 ;
        RECT 5.665 3489.675 5.835 3489.845 ;
        RECT 6.125 3489.675 6.295 3489.845 ;
        RECT 6.585 3489.675 6.755 3489.845 ;
        RECT 2910.105 3489.675 2910.275 3489.845 ;
        RECT 2912.865 3489.675 2913.035 3489.845 ;
        RECT 2913.325 3489.675 2913.495 3489.845 ;
        RECT 2913.785 3489.675 2913.955 3489.845 ;
        RECT 5.665 3484.235 5.835 3484.405 ;
        RECT 6.125 3484.235 6.295 3484.405 ;
        RECT 6.585 3484.235 6.755 3484.405 ;
        RECT 2910.105 3484.235 2910.275 3484.405 ;
        RECT 2912.865 3484.235 2913.035 3484.405 ;
        RECT 2913.325 3484.235 2913.495 3484.405 ;
        RECT 2913.785 3484.235 2913.955 3484.405 ;
        RECT 5.665 3478.795 5.835 3478.965 ;
        RECT 6.125 3478.795 6.295 3478.965 ;
        RECT 6.585 3478.795 6.755 3478.965 ;
        RECT 2910.105 3478.795 2910.275 3478.965 ;
        RECT 2912.865 3478.795 2913.035 3478.965 ;
        RECT 2913.325 3478.795 2913.495 3478.965 ;
        RECT 2913.785 3478.795 2913.955 3478.965 ;
        RECT 5.665 3473.355 5.835 3473.525 ;
        RECT 6.125 3473.355 6.295 3473.525 ;
        RECT 6.585 3473.355 6.755 3473.525 ;
        RECT 2910.105 3473.355 2910.275 3473.525 ;
        RECT 2912.865 3473.355 2913.035 3473.525 ;
        RECT 2913.325 3473.355 2913.495 3473.525 ;
        RECT 2913.785 3473.355 2913.955 3473.525 ;
        RECT 5.665 3467.915 5.835 3468.085 ;
        RECT 6.125 3467.915 6.295 3468.085 ;
        RECT 6.585 3467.915 6.755 3468.085 ;
        RECT 2910.105 3467.915 2910.275 3468.085 ;
        RECT 2912.865 3467.915 2913.035 3468.085 ;
        RECT 2913.325 3467.915 2913.495 3468.085 ;
        RECT 2913.785 3467.915 2913.955 3468.085 ;
        RECT 5.665 3462.475 5.835 3462.645 ;
        RECT 6.125 3462.475 6.295 3462.645 ;
        RECT 6.585 3462.475 6.755 3462.645 ;
        RECT 2910.105 3462.475 2910.275 3462.645 ;
        RECT 2912.865 3462.475 2913.035 3462.645 ;
        RECT 2913.325 3462.475 2913.495 3462.645 ;
        RECT 2913.785 3462.475 2913.955 3462.645 ;
        RECT 5.665 3457.035 5.835 3457.205 ;
        RECT 6.125 3457.035 6.295 3457.205 ;
        RECT 6.585 3457.035 6.755 3457.205 ;
        RECT 2910.105 3457.035 2910.275 3457.205 ;
        RECT 2912.865 3457.035 2913.035 3457.205 ;
        RECT 2913.325 3457.035 2913.495 3457.205 ;
        RECT 2913.785 3457.035 2913.955 3457.205 ;
        RECT 5.665 3451.595 5.835 3451.765 ;
        RECT 6.125 3451.595 6.295 3451.765 ;
        RECT 6.585 3451.595 6.755 3451.765 ;
        RECT 2910.105 3451.595 2910.275 3451.765 ;
        RECT 2912.865 3451.595 2913.035 3451.765 ;
        RECT 2913.325 3451.595 2913.495 3451.765 ;
        RECT 2913.785 3451.595 2913.955 3451.765 ;
        RECT 5.665 3446.155 5.835 3446.325 ;
        RECT 6.125 3446.155 6.295 3446.325 ;
        RECT 6.585 3446.155 6.755 3446.325 ;
        RECT 2910.105 3446.155 2910.275 3446.325 ;
        RECT 2912.865 3446.155 2913.035 3446.325 ;
        RECT 2913.325 3446.155 2913.495 3446.325 ;
        RECT 2913.785 3446.155 2913.955 3446.325 ;
        RECT 5.665 3440.715 5.835 3440.885 ;
        RECT 6.125 3440.715 6.295 3440.885 ;
        RECT 6.585 3440.715 6.755 3440.885 ;
        RECT 2910.105 3440.715 2910.275 3440.885 ;
        RECT 2912.865 3440.715 2913.035 3440.885 ;
        RECT 2913.325 3440.715 2913.495 3440.885 ;
        RECT 2913.785 3440.715 2913.955 3440.885 ;
        RECT 5.665 3435.275 5.835 3435.445 ;
        RECT 6.125 3435.275 6.295 3435.445 ;
        RECT 6.585 3435.275 6.755 3435.445 ;
        RECT 2910.105 3435.275 2910.275 3435.445 ;
        RECT 2912.865 3435.275 2913.035 3435.445 ;
        RECT 2913.325 3435.275 2913.495 3435.445 ;
        RECT 2913.785 3435.275 2913.955 3435.445 ;
        RECT 5.665 3429.835 5.835 3430.005 ;
        RECT 6.125 3429.835 6.295 3430.005 ;
        RECT 6.585 3429.835 6.755 3430.005 ;
        RECT 2910.105 3429.835 2910.275 3430.005 ;
        RECT 2912.865 3429.835 2913.035 3430.005 ;
        RECT 2913.325 3429.835 2913.495 3430.005 ;
        RECT 2913.785 3429.835 2913.955 3430.005 ;
        RECT 5.665 3424.395 5.835 3424.565 ;
        RECT 6.125 3424.395 6.295 3424.565 ;
        RECT 6.585 3424.395 6.755 3424.565 ;
        RECT 2910.105 3424.395 2910.275 3424.565 ;
        RECT 2912.865 3424.395 2913.035 3424.565 ;
        RECT 2913.325 3424.395 2913.495 3424.565 ;
        RECT 2913.785 3424.395 2913.955 3424.565 ;
        RECT 5.665 3418.955 5.835 3419.125 ;
        RECT 6.125 3418.955 6.295 3419.125 ;
        RECT 6.585 3418.955 6.755 3419.125 ;
        RECT 2910.105 3418.955 2910.275 3419.125 ;
        RECT 2912.865 3418.955 2913.035 3419.125 ;
        RECT 2913.325 3418.955 2913.495 3419.125 ;
        RECT 2913.785 3418.955 2913.955 3419.125 ;
        RECT 5.665 3413.515 5.835 3413.685 ;
        RECT 6.125 3413.515 6.295 3413.685 ;
        RECT 6.585 3413.515 6.755 3413.685 ;
        RECT 2910.105 3413.515 2910.275 3413.685 ;
        RECT 2912.865 3413.515 2913.035 3413.685 ;
        RECT 2913.325 3413.515 2913.495 3413.685 ;
        RECT 2913.785 3413.515 2913.955 3413.685 ;
        RECT 5.665 3408.075 5.835 3408.245 ;
        RECT 6.125 3408.075 6.295 3408.245 ;
        RECT 6.585 3408.075 6.755 3408.245 ;
        RECT 2910.105 3408.075 2910.275 3408.245 ;
        RECT 2912.865 3408.075 2913.035 3408.245 ;
        RECT 2913.325 3408.075 2913.495 3408.245 ;
        RECT 2913.785 3408.075 2913.955 3408.245 ;
        RECT 5.665 3402.635 5.835 3402.805 ;
        RECT 6.125 3402.635 6.295 3402.805 ;
        RECT 6.585 3402.635 6.755 3402.805 ;
        RECT 2909.185 3402.635 2909.355 3402.805 ;
        RECT 2909.645 3402.635 2909.815 3402.805 ;
        RECT 2910.105 3402.635 2910.275 3402.805 ;
        RECT 2912.865 3402.635 2913.035 3402.805 ;
        RECT 2913.325 3402.635 2913.495 3402.805 ;
        RECT 2913.785 3402.635 2913.955 3402.805 ;
        RECT 5.665 3397.195 5.835 3397.365 ;
        RECT 6.125 3397.195 6.295 3397.365 ;
        RECT 6.585 3397.195 6.755 3397.365 ;
        RECT 2910.105 3397.195 2910.275 3397.365 ;
        RECT 2912.865 3397.195 2913.035 3397.365 ;
        RECT 2913.325 3397.195 2913.495 3397.365 ;
        RECT 2913.785 3397.195 2913.955 3397.365 ;
        RECT 5.665 3391.755 5.835 3391.925 ;
        RECT 6.125 3391.755 6.295 3391.925 ;
        RECT 6.585 3391.755 6.755 3391.925 ;
        RECT 2910.105 3391.755 2910.275 3391.925 ;
        RECT 2912.865 3391.755 2913.035 3391.925 ;
        RECT 2913.325 3391.755 2913.495 3391.925 ;
        RECT 2913.785 3391.755 2913.955 3391.925 ;
        RECT 5.665 3386.315 5.835 3386.485 ;
        RECT 6.125 3386.315 6.295 3386.485 ;
        RECT 6.585 3386.315 6.755 3386.485 ;
        RECT 2910.105 3386.315 2910.275 3386.485 ;
        RECT 2912.865 3386.315 2913.035 3386.485 ;
        RECT 2913.325 3386.315 2913.495 3386.485 ;
        RECT 2913.785 3386.315 2913.955 3386.485 ;
        RECT 5.665 3380.875 5.835 3381.045 ;
        RECT 6.125 3380.875 6.295 3381.045 ;
        RECT 6.585 3380.875 6.755 3381.045 ;
        RECT 2910.105 3380.875 2910.275 3381.045 ;
        RECT 2912.865 3380.875 2913.035 3381.045 ;
        RECT 2913.325 3380.875 2913.495 3381.045 ;
        RECT 2913.785 3380.875 2913.955 3381.045 ;
        RECT 5.665 3375.435 5.835 3375.605 ;
        RECT 6.125 3375.435 6.295 3375.605 ;
        RECT 6.585 3375.435 6.755 3375.605 ;
        RECT 2910.105 3375.435 2910.275 3375.605 ;
        RECT 2912.865 3375.435 2913.035 3375.605 ;
        RECT 2913.325 3375.435 2913.495 3375.605 ;
        RECT 2913.785 3375.435 2913.955 3375.605 ;
        RECT 5.665 3369.995 5.835 3370.165 ;
        RECT 6.125 3369.995 6.295 3370.165 ;
        RECT 6.585 3369.995 6.755 3370.165 ;
        RECT 2910.105 3369.995 2910.275 3370.165 ;
        RECT 2912.865 3369.995 2913.035 3370.165 ;
        RECT 2913.325 3369.995 2913.495 3370.165 ;
        RECT 2913.785 3369.995 2913.955 3370.165 ;
        RECT 5.665 3364.555 5.835 3364.725 ;
        RECT 6.125 3364.555 6.295 3364.725 ;
        RECT 6.585 3364.555 6.755 3364.725 ;
        RECT 2910.105 3364.555 2910.275 3364.725 ;
        RECT 2910.565 3364.555 2910.735 3364.725 ;
        RECT 2911.025 3364.555 2911.195 3364.725 ;
        RECT 2911.485 3364.555 2911.655 3364.725 ;
        RECT 2912.865 3364.555 2913.035 3364.725 ;
        RECT 2913.325 3364.555 2913.495 3364.725 ;
        RECT 2913.785 3364.555 2913.955 3364.725 ;
        RECT 5.665 3359.115 5.835 3359.285 ;
        RECT 6.125 3359.115 6.295 3359.285 ;
        RECT 6.585 3359.115 6.755 3359.285 ;
        RECT 2910.105 3359.115 2910.275 3359.285 ;
        RECT 2912.865 3359.115 2913.035 3359.285 ;
        RECT 2913.325 3359.115 2913.495 3359.285 ;
        RECT 2913.785 3359.115 2913.955 3359.285 ;
        RECT 5.665 3353.675 5.835 3353.845 ;
        RECT 6.125 3353.675 6.295 3353.845 ;
        RECT 6.585 3353.675 6.755 3353.845 ;
        RECT 2910.105 3353.675 2910.275 3353.845 ;
        RECT 2912.865 3353.675 2913.035 3353.845 ;
        RECT 2913.325 3353.675 2913.495 3353.845 ;
        RECT 2913.785 3353.675 2913.955 3353.845 ;
        RECT 5.665 3348.235 5.835 3348.405 ;
        RECT 6.125 3348.235 6.295 3348.405 ;
        RECT 6.585 3348.235 6.755 3348.405 ;
        RECT 2910.105 3348.235 2910.275 3348.405 ;
        RECT 2912.865 3348.235 2913.035 3348.405 ;
        RECT 2913.325 3348.235 2913.495 3348.405 ;
        RECT 2913.785 3348.235 2913.955 3348.405 ;
        RECT 5.665 3342.795 5.835 3342.965 ;
        RECT 6.125 3342.795 6.295 3342.965 ;
        RECT 6.585 3342.795 6.755 3342.965 ;
        RECT 2910.105 3342.795 2910.275 3342.965 ;
        RECT 2912.865 3342.795 2913.035 3342.965 ;
        RECT 2913.325 3342.795 2913.495 3342.965 ;
        RECT 2913.785 3342.795 2913.955 3342.965 ;
        RECT 5.665 3337.355 5.835 3337.525 ;
        RECT 6.125 3337.355 6.295 3337.525 ;
        RECT 6.585 3337.355 6.755 3337.525 ;
        RECT 2910.105 3337.355 2910.275 3337.525 ;
        RECT 2912.865 3337.355 2913.035 3337.525 ;
        RECT 2913.325 3337.355 2913.495 3337.525 ;
        RECT 2913.785 3337.355 2913.955 3337.525 ;
        RECT 5.665 3331.915 5.835 3332.085 ;
        RECT 6.125 3331.915 6.295 3332.085 ;
        RECT 6.585 3331.915 6.755 3332.085 ;
        RECT 2910.105 3331.915 2910.275 3332.085 ;
        RECT 2912.865 3331.915 2913.035 3332.085 ;
        RECT 2913.325 3331.915 2913.495 3332.085 ;
        RECT 2913.785 3331.915 2913.955 3332.085 ;
        RECT 5.665 3326.475 5.835 3326.645 ;
        RECT 6.125 3326.475 6.295 3326.645 ;
        RECT 6.585 3326.475 6.755 3326.645 ;
        RECT 2910.105 3326.475 2910.275 3326.645 ;
        RECT 2912.865 3326.475 2913.035 3326.645 ;
        RECT 2913.325 3326.475 2913.495 3326.645 ;
        RECT 2913.785 3326.475 2913.955 3326.645 ;
        RECT 5.665 3321.035 5.835 3321.205 ;
        RECT 6.125 3321.035 6.295 3321.205 ;
        RECT 6.585 3321.035 6.755 3321.205 ;
        RECT 2910.105 3321.035 2910.275 3321.205 ;
        RECT 2912.865 3321.035 2913.035 3321.205 ;
        RECT 2913.325 3321.035 2913.495 3321.205 ;
        RECT 2913.785 3321.035 2913.955 3321.205 ;
        RECT 5.665 3315.595 5.835 3315.765 ;
        RECT 6.125 3315.595 6.295 3315.765 ;
        RECT 6.585 3315.595 6.755 3315.765 ;
        RECT 2910.105 3315.595 2910.275 3315.765 ;
        RECT 2912.865 3315.595 2913.035 3315.765 ;
        RECT 2913.325 3315.595 2913.495 3315.765 ;
        RECT 2913.785 3315.595 2913.955 3315.765 ;
        RECT 5.665 3310.155 5.835 3310.325 ;
        RECT 6.125 3310.155 6.295 3310.325 ;
        RECT 6.585 3310.155 6.755 3310.325 ;
        RECT 2910.105 3310.155 2910.275 3310.325 ;
        RECT 2912.865 3310.155 2913.035 3310.325 ;
        RECT 2913.325 3310.155 2913.495 3310.325 ;
        RECT 2913.785 3310.155 2913.955 3310.325 ;
        RECT 5.665 3304.715 5.835 3304.885 ;
        RECT 6.125 3304.715 6.295 3304.885 ;
        RECT 6.585 3304.715 6.755 3304.885 ;
        RECT 2910.105 3304.715 2910.275 3304.885 ;
        RECT 2912.865 3304.715 2913.035 3304.885 ;
        RECT 2913.325 3304.715 2913.495 3304.885 ;
        RECT 2913.785 3304.715 2913.955 3304.885 ;
        RECT 5.665 3299.275 5.835 3299.445 ;
        RECT 6.125 3299.275 6.295 3299.445 ;
        RECT 6.585 3299.275 6.755 3299.445 ;
        RECT 2910.105 3299.275 2910.275 3299.445 ;
        RECT 2912.865 3299.275 2913.035 3299.445 ;
        RECT 2913.325 3299.275 2913.495 3299.445 ;
        RECT 2913.785 3299.275 2913.955 3299.445 ;
        RECT 5.665 3293.835 5.835 3294.005 ;
        RECT 6.125 3293.835 6.295 3294.005 ;
        RECT 6.585 3293.835 6.755 3294.005 ;
        RECT 2910.105 3293.835 2910.275 3294.005 ;
        RECT 2912.865 3293.835 2913.035 3294.005 ;
        RECT 2913.325 3293.835 2913.495 3294.005 ;
        RECT 2913.785 3293.835 2913.955 3294.005 ;
        RECT 5.665 3288.395 5.835 3288.565 ;
        RECT 6.125 3288.395 6.295 3288.565 ;
        RECT 6.585 3288.395 6.755 3288.565 ;
        RECT 2910.105 3288.395 2910.275 3288.565 ;
        RECT 2912.865 3288.395 2913.035 3288.565 ;
        RECT 2913.325 3288.395 2913.495 3288.565 ;
        RECT 2913.785 3288.395 2913.955 3288.565 ;
        RECT 5.665 3282.955 5.835 3283.125 ;
        RECT 6.125 3282.955 6.295 3283.125 ;
        RECT 6.585 3282.955 6.755 3283.125 ;
        RECT 2910.105 3282.955 2910.275 3283.125 ;
        RECT 2912.865 3282.955 2913.035 3283.125 ;
        RECT 2913.325 3282.955 2913.495 3283.125 ;
        RECT 2913.785 3282.955 2913.955 3283.125 ;
        RECT 5.665 3277.515 5.835 3277.685 ;
        RECT 6.125 3277.515 6.295 3277.685 ;
        RECT 6.585 3277.515 6.755 3277.685 ;
        RECT 2910.105 3277.515 2910.275 3277.685 ;
        RECT 2912.865 3277.515 2913.035 3277.685 ;
        RECT 2913.325 3277.515 2913.495 3277.685 ;
        RECT 2913.785 3277.515 2913.955 3277.685 ;
        RECT 5.665 3272.075 5.835 3272.245 ;
        RECT 6.125 3272.075 6.295 3272.245 ;
        RECT 6.585 3272.075 6.755 3272.245 ;
        RECT 2910.105 3272.075 2910.275 3272.245 ;
        RECT 2912.865 3272.075 2913.035 3272.245 ;
        RECT 2913.325 3272.075 2913.495 3272.245 ;
        RECT 2913.785 3272.075 2913.955 3272.245 ;
        RECT 5.665 3266.635 5.835 3266.805 ;
        RECT 6.125 3266.635 6.295 3266.805 ;
        RECT 6.585 3266.635 6.755 3266.805 ;
        RECT 2910.105 3266.635 2910.275 3266.805 ;
        RECT 2912.865 3266.635 2913.035 3266.805 ;
        RECT 2913.325 3266.635 2913.495 3266.805 ;
        RECT 2913.785 3266.635 2913.955 3266.805 ;
        RECT 5.665 3261.195 5.835 3261.365 ;
        RECT 6.125 3261.195 6.295 3261.365 ;
        RECT 6.585 3261.195 6.755 3261.365 ;
        RECT 2910.105 3261.195 2910.275 3261.365 ;
        RECT 2912.865 3261.195 2913.035 3261.365 ;
        RECT 2913.325 3261.195 2913.495 3261.365 ;
        RECT 2913.785 3261.195 2913.955 3261.365 ;
        RECT 5.665 3255.755 5.835 3255.925 ;
        RECT 6.125 3255.755 6.295 3255.925 ;
        RECT 6.585 3255.755 6.755 3255.925 ;
        RECT 2910.105 3255.755 2910.275 3255.925 ;
        RECT 2912.865 3255.755 2913.035 3255.925 ;
        RECT 2913.325 3255.755 2913.495 3255.925 ;
        RECT 2913.785 3255.755 2913.955 3255.925 ;
        RECT 5.665 3250.315 5.835 3250.485 ;
        RECT 6.125 3250.315 6.295 3250.485 ;
        RECT 6.585 3250.315 6.755 3250.485 ;
        RECT 2910.105 3250.315 2910.275 3250.485 ;
        RECT 2912.865 3250.315 2913.035 3250.485 ;
        RECT 2913.325 3250.315 2913.495 3250.485 ;
        RECT 2913.785 3250.315 2913.955 3250.485 ;
        RECT 5.665 3244.875 5.835 3245.045 ;
        RECT 6.125 3244.875 6.295 3245.045 ;
        RECT 6.585 3244.875 6.755 3245.045 ;
        RECT 2910.105 3244.875 2910.275 3245.045 ;
        RECT 2912.865 3244.875 2913.035 3245.045 ;
        RECT 2913.325 3244.875 2913.495 3245.045 ;
        RECT 2913.785 3244.875 2913.955 3245.045 ;
        RECT 5.665 3239.435 5.835 3239.605 ;
        RECT 6.125 3239.435 6.295 3239.605 ;
        RECT 6.585 3239.435 6.755 3239.605 ;
        RECT 2910.105 3239.435 2910.275 3239.605 ;
        RECT 2912.865 3239.435 2913.035 3239.605 ;
        RECT 2913.325 3239.435 2913.495 3239.605 ;
        RECT 2913.785 3239.435 2913.955 3239.605 ;
        RECT 5.665 3233.995 5.835 3234.165 ;
        RECT 6.125 3233.995 6.295 3234.165 ;
        RECT 6.585 3233.995 6.755 3234.165 ;
        RECT 2910.105 3233.995 2910.275 3234.165 ;
        RECT 2912.865 3233.995 2913.035 3234.165 ;
        RECT 2913.325 3233.995 2913.495 3234.165 ;
        RECT 2913.785 3233.995 2913.955 3234.165 ;
        RECT 5.665 3228.555 5.835 3228.725 ;
        RECT 6.125 3228.555 6.295 3228.725 ;
        RECT 6.585 3228.555 6.755 3228.725 ;
        RECT 2910.105 3228.555 2910.275 3228.725 ;
        RECT 2912.865 3228.555 2913.035 3228.725 ;
        RECT 2913.325 3228.555 2913.495 3228.725 ;
        RECT 2913.785 3228.555 2913.955 3228.725 ;
        RECT 5.665 3223.115 5.835 3223.285 ;
        RECT 6.125 3223.115 6.295 3223.285 ;
        RECT 6.585 3223.115 6.755 3223.285 ;
        RECT 8.885 3223.115 9.055 3223.285 ;
        RECT 9.345 3223.115 9.515 3223.285 ;
        RECT 9.805 3223.115 9.975 3223.285 ;
        RECT 2910.105 3223.115 2910.275 3223.285 ;
        RECT 2912.865 3223.115 2913.035 3223.285 ;
        RECT 2913.325 3223.115 2913.495 3223.285 ;
        RECT 2913.785 3223.115 2913.955 3223.285 ;
        RECT 5.665 3217.675 5.835 3217.845 ;
        RECT 6.125 3217.675 6.295 3217.845 ;
        RECT 6.585 3217.675 6.755 3217.845 ;
        RECT 2910.105 3217.675 2910.275 3217.845 ;
        RECT 2912.865 3217.675 2913.035 3217.845 ;
        RECT 2913.325 3217.675 2913.495 3217.845 ;
        RECT 2913.785 3217.675 2913.955 3217.845 ;
        RECT 5.665 3212.235 5.835 3212.405 ;
        RECT 6.125 3212.235 6.295 3212.405 ;
        RECT 6.585 3212.235 6.755 3212.405 ;
        RECT 2910.105 3212.235 2910.275 3212.405 ;
        RECT 2912.865 3212.235 2913.035 3212.405 ;
        RECT 2913.325 3212.235 2913.495 3212.405 ;
        RECT 2913.785 3212.235 2913.955 3212.405 ;
        RECT 5.665 3206.795 5.835 3206.965 ;
        RECT 6.125 3206.795 6.295 3206.965 ;
        RECT 6.585 3206.795 6.755 3206.965 ;
        RECT 2910.105 3206.795 2910.275 3206.965 ;
        RECT 2912.865 3206.795 2913.035 3206.965 ;
        RECT 2913.325 3206.795 2913.495 3206.965 ;
        RECT 2913.785 3206.795 2913.955 3206.965 ;
        RECT 5.665 3201.355 5.835 3201.525 ;
        RECT 6.125 3201.355 6.295 3201.525 ;
        RECT 6.585 3201.355 6.755 3201.525 ;
        RECT 2910.105 3201.355 2910.275 3201.525 ;
        RECT 2910.565 3201.355 2910.735 3201.525 ;
        RECT 2911.025 3201.355 2911.195 3201.525 ;
        RECT 2911.485 3201.355 2911.655 3201.525 ;
        RECT 2912.865 3201.355 2913.035 3201.525 ;
        RECT 2913.325 3201.355 2913.495 3201.525 ;
        RECT 2913.785 3201.355 2913.955 3201.525 ;
        RECT 5.665 3195.915 5.835 3196.085 ;
        RECT 6.125 3195.915 6.295 3196.085 ;
        RECT 6.585 3195.915 6.755 3196.085 ;
        RECT 2910.105 3195.915 2910.275 3196.085 ;
        RECT 2912.865 3195.915 2913.035 3196.085 ;
        RECT 2913.325 3195.915 2913.495 3196.085 ;
        RECT 2913.785 3195.915 2913.955 3196.085 ;
        RECT 5.665 3190.475 5.835 3190.645 ;
        RECT 6.125 3190.475 6.295 3190.645 ;
        RECT 6.585 3190.475 6.755 3190.645 ;
        RECT 2910.105 3190.475 2910.275 3190.645 ;
        RECT 2912.865 3190.475 2913.035 3190.645 ;
        RECT 2913.325 3190.475 2913.495 3190.645 ;
        RECT 2913.785 3190.475 2913.955 3190.645 ;
        RECT 5.665 3185.035 5.835 3185.205 ;
        RECT 6.125 3185.035 6.295 3185.205 ;
        RECT 6.585 3185.035 6.755 3185.205 ;
        RECT 2910.105 3185.035 2910.275 3185.205 ;
        RECT 2912.865 3185.035 2913.035 3185.205 ;
        RECT 2913.325 3185.035 2913.495 3185.205 ;
        RECT 2913.785 3185.035 2913.955 3185.205 ;
        RECT 5.665 3179.595 5.835 3179.765 ;
        RECT 6.125 3179.595 6.295 3179.765 ;
        RECT 6.585 3179.595 6.755 3179.765 ;
        RECT 2910.105 3179.595 2910.275 3179.765 ;
        RECT 2912.865 3179.595 2913.035 3179.765 ;
        RECT 2913.325 3179.595 2913.495 3179.765 ;
        RECT 2913.785 3179.595 2913.955 3179.765 ;
        RECT 5.665 3174.155 5.835 3174.325 ;
        RECT 6.125 3174.155 6.295 3174.325 ;
        RECT 6.585 3174.155 6.755 3174.325 ;
        RECT 2910.105 3174.155 2910.275 3174.325 ;
        RECT 2912.865 3174.155 2913.035 3174.325 ;
        RECT 2913.325 3174.155 2913.495 3174.325 ;
        RECT 2913.785 3174.155 2913.955 3174.325 ;
        RECT 5.665 3168.715 5.835 3168.885 ;
        RECT 6.125 3168.715 6.295 3168.885 ;
        RECT 6.585 3168.715 6.755 3168.885 ;
        RECT 2910.105 3168.715 2910.275 3168.885 ;
        RECT 2912.865 3168.715 2913.035 3168.885 ;
        RECT 2913.325 3168.715 2913.495 3168.885 ;
        RECT 2913.785 3168.715 2913.955 3168.885 ;
        RECT 5.665 3163.275 5.835 3163.445 ;
        RECT 6.125 3163.275 6.295 3163.445 ;
        RECT 6.585 3163.275 6.755 3163.445 ;
        RECT 2910.105 3163.275 2910.275 3163.445 ;
        RECT 2912.865 3163.275 2913.035 3163.445 ;
        RECT 2913.325 3163.275 2913.495 3163.445 ;
        RECT 2913.785 3163.275 2913.955 3163.445 ;
        RECT 5.665 3157.835 5.835 3158.005 ;
        RECT 6.125 3157.835 6.295 3158.005 ;
        RECT 6.585 3157.835 6.755 3158.005 ;
        RECT 2910.105 3157.835 2910.275 3158.005 ;
        RECT 2912.865 3157.835 2913.035 3158.005 ;
        RECT 2913.325 3157.835 2913.495 3158.005 ;
        RECT 2913.785 3157.835 2913.955 3158.005 ;
        RECT 5.665 3152.395 5.835 3152.565 ;
        RECT 6.125 3152.395 6.295 3152.565 ;
        RECT 6.585 3152.395 6.755 3152.565 ;
        RECT 2910.105 3152.395 2910.275 3152.565 ;
        RECT 2912.865 3152.395 2913.035 3152.565 ;
        RECT 2913.325 3152.395 2913.495 3152.565 ;
        RECT 2913.785 3152.395 2913.955 3152.565 ;
        RECT 5.665 3146.955 5.835 3147.125 ;
        RECT 6.125 3146.955 6.295 3147.125 ;
        RECT 6.585 3146.955 6.755 3147.125 ;
        RECT 2910.105 3146.955 2910.275 3147.125 ;
        RECT 2912.865 3146.955 2913.035 3147.125 ;
        RECT 2913.325 3146.955 2913.495 3147.125 ;
        RECT 2913.785 3146.955 2913.955 3147.125 ;
        RECT 5.665 3141.515 5.835 3141.685 ;
        RECT 6.125 3141.515 6.295 3141.685 ;
        RECT 6.585 3141.515 6.755 3141.685 ;
        RECT 2910.105 3141.515 2910.275 3141.685 ;
        RECT 2912.865 3141.515 2913.035 3141.685 ;
        RECT 2913.325 3141.515 2913.495 3141.685 ;
        RECT 2913.785 3141.515 2913.955 3141.685 ;
        RECT 5.665 3136.075 5.835 3136.245 ;
        RECT 6.125 3136.075 6.295 3136.245 ;
        RECT 6.585 3136.075 6.755 3136.245 ;
        RECT 2910.105 3136.075 2910.275 3136.245 ;
        RECT 2912.865 3136.075 2913.035 3136.245 ;
        RECT 2913.325 3136.075 2913.495 3136.245 ;
        RECT 2913.785 3136.075 2913.955 3136.245 ;
        RECT 5.665 3130.635 5.835 3130.805 ;
        RECT 6.125 3130.635 6.295 3130.805 ;
        RECT 6.585 3130.635 6.755 3130.805 ;
        RECT 2910.105 3130.635 2910.275 3130.805 ;
        RECT 2912.865 3130.635 2913.035 3130.805 ;
        RECT 2913.325 3130.635 2913.495 3130.805 ;
        RECT 2913.785 3130.635 2913.955 3130.805 ;
        RECT 5.665 3125.195 5.835 3125.365 ;
        RECT 6.125 3125.195 6.295 3125.365 ;
        RECT 6.585 3125.195 6.755 3125.365 ;
        RECT 2910.105 3125.195 2910.275 3125.365 ;
        RECT 2912.865 3125.195 2913.035 3125.365 ;
        RECT 2913.325 3125.195 2913.495 3125.365 ;
        RECT 2913.785 3125.195 2913.955 3125.365 ;
        RECT 5.665 3119.755 5.835 3119.925 ;
        RECT 6.125 3119.755 6.295 3119.925 ;
        RECT 6.585 3119.755 6.755 3119.925 ;
        RECT 2910.105 3119.755 2910.275 3119.925 ;
        RECT 2912.865 3119.755 2913.035 3119.925 ;
        RECT 2913.325 3119.755 2913.495 3119.925 ;
        RECT 2913.785 3119.755 2913.955 3119.925 ;
        RECT 5.665 3114.315 5.835 3114.485 ;
        RECT 6.125 3114.315 6.295 3114.485 ;
        RECT 6.585 3114.315 6.755 3114.485 ;
        RECT 2910.105 3114.315 2910.275 3114.485 ;
        RECT 2912.865 3114.315 2913.035 3114.485 ;
        RECT 2913.325 3114.315 2913.495 3114.485 ;
        RECT 2913.785 3114.315 2913.955 3114.485 ;
        RECT 5.665 3108.875 5.835 3109.045 ;
        RECT 6.125 3108.875 6.295 3109.045 ;
        RECT 6.585 3108.875 6.755 3109.045 ;
        RECT 2910.105 3108.875 2910.275 3109.045 ;
        RECT 2912.865 3108.875 2913.035 3109.045 ;
        RECT 2913.325 3108.875 2913.495 3109.045 ;
        RECT 2913.785 3108.875 2913.955 3109.045 ;
        RECT 5.665 3103.435 5.835 3103.605 ;
        RECT 6.125 3103.435 6.295 3103.605 ;
        RECT 6.585 3103.435 6.755 3103.605 ;
        RECT 2910.105 3103.435 2910.275 3103.605 ;
        RECT 2912.865 3103.435 2913.035 3103.605 ;
        RECT 2913.325 3103.435 2913.495 3103.605 ;
        RECT 2913.785 3103.435 2913.955 3103.605 ;
        RECT 5.665 3097.995 5.835 3098.165 ;
        RECT 6.125 3097.995 6.295 3098.165 ;
        RECT 6.585 3097.995 6.755 3098.165 ;
        RECT 2909.185 3097.995 2909.355 3098.165 ;
        RECT 2909.645 3097.995 2909.815 3098.165 ;
        RECT 2910.105 3097.995 2910.275 3098.165 ;
        RECT 2912.865 3097.995 2913.035 3098.165 ;
        RECT 2913.325 3097.995 2913.495 3098.165 ;
        RECT 2913.785 3097.995 2913.955 3098.165 ;
        RECT 5.665 3092.555 5.835 3092.725 ;
        RECT 6.125 3092.555 6.295 3092.725 ;
        RECT 6.585 3092.555 6.755 3092.725 ;
        RECT 2910.105 3092.555 2910.275 3092.725 ;
        RECT 2912.865 3092.555 2913.035 3092.725 ;
        RECT 2913.325 3092.555 2913.495 3092.725 ;
        RECT 2913.785 3092.555 2913.955 3092.725 ;
        RECT 5.665 3087.115 5.835 3087.285 ;
        RECT 6.125 3087.115 6.295 3087.285 ;
        RECT 6.585 3087.115 6.755 3087.285 ;
        RECT 2910.105 3087.115 2910.275 3087.285 ;
        RECT 2912.865 3087.115 2913.035 3087.285 ;
        RECT 2913.325 3087.115 2913.495 3087.285 ;
        RECT 2913.785 3087.115 2913.955 3087.285 ;
        RECT 5.665 3081.675 5.835 3081.845 ;
        RECT 6.125 3081.675 6.295 3081.845 ;
        RECT 6.585 3081.675 6.755 3081.845 ;
        RECT 2910.105 3081.675 2910.275 3081.845 ;
        RECT 2912.865 3081.675 2913.035 3081.845 ;
        RECT 2913.325 3081.675 2913.495 3081.845 ;
        RECT 2913.785 3081.675 2913.955 3081.845 ;
        RECT 5.665 3076.235 5.835 3076.405 ;
        RECT 6.125 3076.235 6.295 3076.405 ;
        RECT 6.585 3076.235 6.755 3076.405 ;
        RECT 2910.105 3076.235 2910.275 3076.405 ;
        RECT 2912.865 3076.235 2913.035 3076.405 ;
        RECT 2913.325 3076.235 2913.495 3076.405 ;
        RECT 2913.785 3076.235 2913.955 3076.405 ;
        RECT 5.665 3070.795 5.835 3070.965 ;
        RECT 6.125 3070.795 6.295 3070.965 ;
        RECT 6.585 3070.795 6.755 3070.965 ;
        RECT 2910.105 3070.795 2910.275 3070.965 ;
        RECT 2912.865 3070.795 2913.035 3070.965 ;
        RECT 2913.325 3070.795 2913.495 3070.965 ;
        RECT 2913.785 3070.795 2913.955 3070.965 ;
        RECT 5.665 3065.355 5.835 3065.525 ;
        RECT 6.125 3065.355 6.295 3065.525 ;
        RECT 6.585 3065.355 6.755 3065.525 ;
        RECT 2910.105 3065.355 2910.275 3065.525 ;
        RECT 2912.865 3065.355 2913.035 3065.525 ;
        RECT 2913.325 3065.355 2913.495 3065.525 ;
        RECT 2913.785 3065.355 2913.955 3065.525 ;
        RECT 5.665 3059.915 5.835 3060.085 ;
        RECT 6.125 3059.915 6.295 3060.085 ;
        RECT 6.585 3059.915 6.755 3060.085 ;
        RECT 2910.105 3059.915 2910.275 3060.085 ;
        RECT 2912.865 3059.915 2913.035 3060.085 ;
        RECT 2913.325 3059.915 2913.495 3060.085 ;
        RECT 2913.785 3059.915 2913.955 3060.085 ;
        RECT 5.665 3054.475 5.835 3054.645 ;
        RECT 6.125 3054.475 6.295 3054.645 ;
        RECT 6.585 3054.475 6.755 3054.645 ;
        RECT 2910.105 3054.475 2910.275 3054.645 ;
        RECT 2912.865 3054.475 2913.035 3054.645 ;
        RECT 2913.325 3054.475 2913.495 3054.645 ;
        RECT 2913.785 3054.475 2913.955 3054.645 ;
        RECT 5.665 3049.035 5.835 3049.205 ;
        RECT 6.125 3049.035 6.295 3049.205 ;
        RECT 6.585 3049.035 6.755 3049.205 ;
        RECT 2910.105 3049.035 2910.275 3049.205 ;
        RECT 2912.865 3049.035 2913.035 3049.205 ;
        RECT 2913.325 3049.035 2913.495 3049.205 ;
        RECT 2913.785 3049.035 2913.955 3049.205 ;
        RECT 5.665 3043.595 5.835 3043.765 ;
        RECT 6.125 3043.595 6.295 3043.765 ;
        RECT 6.585 3043.595 6.755 3043.765 ;
        RECT 2910.105 3043.595 2910.275 3043.765 ;
        RECT 2912.865 3043.595 2913.035 3043.765 ;
        RECT 2913.325 3043.595 2913.495 3043.765 ;
        RECT 2913.785 3043.595 2913.955 3043.765 ;
        RECT 5.665 3038.155 5.835 3038.325 ;
        RECT 6.125 3038.155 6.295 3038.325 ;
        RECT 6.585 3038.155 6.755 3038.325 ;
        RECT 2910.105 3038.155 2910.275 3038.325 ;
        RECT 2912.865 3038.155 2913.035 3038.325 ;
        RECT 2913.325 3038.155 2913.495 3038.325 ;
        RECT 2913.785 3038.155 2913.955 3038.325 ;
        RECT 5.665 3032.715 5.835 3032.885 ;
        RECT 6.125 3032.715 6.295 3032.885 ;
        RECT 6.585 3032.715 6.755 3032.885 ;
        RECT 2910.105 3032.715 2910.275 3032.885 ;
        RECT 2912.865 3032.715 2913.035 3032.885 ;
        RECT 2913.325 3032.715 2913.495 3032.885 ;
        RECT 2913.785 3032.715 2913.955 3032.885 ;
        RECT 5.665 3027.275 5.835 3027.445 ;
        RECT 6.125 3027.275 6.295 3027.445 ;
        RECT 6.585 3027.275 6.755 3027.445 ;
        RECT 2910.105 3027.275 2910.275 3027.445 ;
        RECT 2912.865 3027.275 2913.035 3027.445 ;
        RECT 2913.325 3027.275 2913.495 3027.445 ;
        RECT 2913.785 3027.275 2913.955 3027.445 ;
        RECT 5.665 3021.835 5.835 3022.005 ;
        RECT 6.125 3021.835 6.295 3022.005 ;
        RECT 6.585 3021.835 6.755 3022.005 ;
        RECT 2910.105 3021.835 2910.275 3022.005 ;
        RECT 2912.865 3021.835 2913.035 3022.005 ;
        RECT 2913.325 3021.835 2913.495 3022.005 ;
        RECT 2913.785 3021.835 2913.955 3022.005 ;
        RECT 5.665 3016.395 5.835 3016.565 ;
        RECT 6.125 3016.395 6.295 3016.565 ;
        RECT 6.585 3016.395 6.755 3016.565 ;
        RECT 2910.105 3016.395 2910.275 3016.565 ;
        RECT 2912.865 3016.395 2913.035 3016.565 ;
        RECT 2913.325 3016.395 2913.495 3016.565 ;
        RECT 2913.785 3016.395 2913.955 3016.565 ;
        RECT 5.665 3010.955 5.835 3011.125 ;
        RECT 6.125 3010.955 6.295 3011.125 ;
        RECT 6.585 3010.955 6.755 3011.125 ;
        RECT 8.885 3010.955 9.055 3011.125 ;
        RECT 9.345 3010.955 9.515 3011.125 ;
        RECT 9.805 3010.955 9.975 3011.125 ;
        RECT 2910.105 3010.955 2910.275 3011.125 ;
        RECT 2912.865 3010.955 2913.035 3011.125 ;
        RECT 2913.325 3010.955 2913.495 3011.125 ;
        RECT 2913.785 3010.955 2913.955 3011.125 ;
        RECT 5.665 3005.515 5.835 3005.685 ;
        RECT 6.125 3005.515 6.295 3005.685 ;
        RECT 6.585 3005.515 6.755 3005.685 ;
        RECT 2910.105 3005.515 2910.275 3005.685 ;
        RECT 2912.865 3005.515 2913.035 3005.685 ;
        RECT 2913.325 3005.515 2913.495 3005.685 ;
        RECT 2913.785 3005.515 2913.955 3005.685 ;
        RECT 5.665 3000.075 5.835 3000.245 ;
        RECT 6.125 3000.075 6.295 3000.245 ;
        RECT 6.585 3000.075 6.755 3000.245 ;
        RECT 2910.105 3000.075 2910.275 3000.245 ;
        RECT 2912.865 3000.075 2913.035 3000.245 ;
        RECT 2913.325 3000.075 2913.495 3000.245 ;
        RECT 2913.785 3000.075 2913.955 3000.245 ;
        RECT 5.665 2994.635 5.835 2994.805 ;
        RECT 6.125 2994.635 6.295 2994.805 ;
        RECT 6.585 2994.635 6.755 2994.805 ;
        RECT 2910.105 2994.635 2910.275 2994.805 ;
        RECT 2912.865 2994.635 2913.035 2994.805 ;
        RECT 2913.325 2994.635 2913.495 2994.805 ;
        RECT 2913.785 2994.635 2913.955 2994.805 ;
        RECT 5.665 2989.195 5.835 2989.365 ;
        RECT 6.125 2989.195 6.295 2989.365 ;
        RECT 6.585 2989.195 6.755 2989.365 ;
        RECT 2910.105 2989.195 2910.275 2989.365 ;
        RECT 2912.865 2989.195 2913.035 2989.365 ;
        RECT 2913.325 2989.195 2913.495 2989.365 ;
        RECT 2913.785 2989.195 2913.955 2989.365 ;
        RECT 5.665 2983.755 5.835 2983.925 ;
        RECT 6.125 2983.755 6.295 2983.925 ;
        RECT 6.585 2983.755 6.755 2983.925 ;
        RECT 2910.105 2983.755 2910.275 2983.925 ;
        RECT 2912.865 2983.755 2913.035 2983.925 ;
        RECT 2913.325 2983.755 2913.495 2983.925 ;
        RECT 2913.785 2983.755 2913.955 2983.925 ;
        RECT 5.665 2978.315 5.835 2978.485 ;
        RECT 6.125 2978.315 6.295 2978.485 ;
        RECT 6.585 2978.315 6.755 2978.485 ;
        RECT 2910.105 2978.315 2910.275 2978.485 ;
        RECT 2912.865 2978.315 2913.035 2978.485 ;
        RECT 2913.325 2978.315 2913.495 2978.485 ;
        RECT 2913.785 2978.315 2913.955 2978.485 ;
        RECT 5.665 2972.875 5.835 2973.045 ;
        RECT 6.125 2972.875 6.295 2973.045 ;
        RECT 6.585 2972.875 6.755 2973.045 ;
        RECT 8.885 2972.875 9.055 2973.045 ;
        RECT 9.345 2972.875 9.515 2973.045 ;
        RECT 9.805 2972.875 9.975 2973.045 ;
        RECT 2910.105 2972.875 2910.275 2973.045 ;
        RECT 2912.865 2972.875 2913.035 2973.045 ;
        RECT 2913.325 2972.875 2913.495 2973.045 ;
        RECT 2913.785 2972.875 2913.955 2973.045 ;
        RECT 5.665 2967.435 5.835 2967.605 ;
        RECT 6.125 2967.435 6.295 2967.605 ;
        RECT 6.585 2967.435 6.755 2967.605 ;
        RECT 2910.105 2967.435 2910.275 2967.605 ;
        RECT 2912.865 2967.435 2913.035 2967.605 ;
        RECT 2913.325 2967.435 2913.495 2967.605 ;
        RECT 2913.785 2967.435 2913.955 2967.605 ;
        RECT 5.665 2961.995 5.835 2962.165 ;
        RECT 6.125 2961.995 6.295 2962.165 ;
        RECT 6.585 2961.995 6.755 2962.165 ;
        RECT 2910.105 2961.995 2910.275 2962.165 ;
        RECT 2912.865 2961.995 2913.035 2962.165 ;
        RECT 2913.325 2961.995 2913.495 2962.165 ;
        RECT 2913.785 2961.995 2913.955 2962.165 ;
        RECT 5.665 2956.555 5.835 2956.725 ;
        RECT 6.125 2956.555 6.295 2956.725 ;
        RECT 6.585 2956.555 6.755 2956.725 ;
        RECT 8.885 2956.555 9.055 2956.725 ;
        RECT 9.345 2956.555 9.515 2956.725 ;
        RECT 9.805 2956.555 9.975 2956.725 ;
        RECT 2910.105 2956.555 2910.275 2956.725 ;
        RECT 2912.865 2956.555 2913.035 2956.725 ;
        RECT 2913.325 2956.555 2913.495 2956.725 ;
        RECT 2913.785 2956.555 2913.955 2956.725 ;
        RECT 5.665 2951.115 5.835 2951.285 ;
        RECT 6.125 2951.115 6.295 2951.285 ;
        RECT 6.585 2951.115 6.755 2951.285 ;
        RECT 2910.105 2951.115 2910.275 2951.285 ;
        RECT 2912.865 2951.115 2913.035 2951.285 ;
        RECT 2913.325 2951.115 2913.495 2951.285 ;
        RECT 2913.785 2951.115 2913.955 2951.285 ;
        RECT 5.665 2945.675 5.835 2945.845 ;
        RECT 6.125 2945.675 6.295 2945.845 ;
        RECT 6.585 2945.675 6.755 2945.845 ;
        RECT 2910.105 2945.675 2910.275 2945.845 ;
        RECT 2912.865 2945.675 2913.035 2945.845 ;
        RECT 2913.325 2945.675 2913.495 2945.845 ;
        RECT 2913.785 2945.675 2913.955 2945.845 ;
        RECT 5.665 2940.235 5.835 2940.405 ;
        RECT 6.125 2940.235 6.295 2940.405 ;
        RECT 6.585 2940.235 6.755 2940.405 ;
        RECT 2910.105 2940.235 2910.275 2940.405 ;
        RECT 2912.865 2940.235 2913.035 2940.405 ;
        RECT 2913.325 2940.235 2913.495 2940.405 ;
        RECT 2913.785 2940.235 2913.955 2940.405 ;
        RECT 5.665 2934.795 5.835 2934.965 ;
        RECT 6.125 2934.795 6.295 2934.965 ;
        RECT 6.585 2934.795 6.755 2934.965 ;
        RECT 2910.105 2934.795 2910.275 2934.965 ;
        RECT 2912.865 2934.795 2913.035 2934.965 ;
        RECT 2913.325 2934.795 2913.495 2934.965 ;
        RECT 2913.785 2934.795 2913.955 2934.965 ;
        RECT 5.665 2929.355 5.835 2929.525 ;
        RECT 6.125 2929.355 6.295 2929.525 ;
        RECT 6.585 2929.355 6.755 2929.525 ;
        RECT 2910.105 2929.355 2910.275 2929.525 ;
        RECT 2912.865 2929.355 2913.035 2929.525 ;
        RECT 2913.325 2929.355 2913.495 2929.525 ;
        RECT 2913.785 2929.355 2913.955 2929.525 ;
        RECT 5.665 2923.915 5.835 2924.085 ;
        RECT 6.125 2923.915 6.295 2924.085 ;
        RECT 6.585 2923.915 6.755 2924.085 ;
        RECT 2910.105 2923.915 2910.275 2924.085 ;
        RECT 2912.865 2923.915 2913.035 2924.085 ;
        RECT 2913.325 2923.915 2913.495 2924.085 ;
        RECT 2913.785 2923.915 2913.955 2924.085 ;
        RECT 5.665 2918.475 5.835 2918.645 ;
        RECT 6.125 2918.475 6.295 2918.645 ;
        RECT 6.585 2918.475 6.755 2918.645 ;
        RECT 2910.105 2918.475 2910.275 2918.645 ;
        RECT 2912.865 2918.475 2913.035 2918.645 ;
        RECT 2913.325 2918.475 2913.495 2918.645 ;
        RECT 2913.785 2918.475 2913.955 2918.645 ;
        RECT 5.665 2913.035 5.835 2913.205 ;
        RECT 6.125 2913.035 6.295 2913.205 ;
        RECT 6.585 2913.035 6.755 2913.205 ;
        RECT 2910.105 2913.035 2910.275 2913.205 ;
        RECT 2910.565 2913.035 2910.735 2913.205 ;
        RECT 2911.025 2913.035 2911.195 2913.205 ;
        RECT 2911.485 2913.035 2911.655 2913.205 ;
        RECT 2912.865 2913.035 2913.035 2913.205 ;
        RECT 2913.325 2913.035 2913.495 2913.205 ;
        RECT 2913.785 2913.035 2913.955 2913.205 ;
        RECT 5.665 2907.595 5.835 2907.765 ;
        RECT 6.125 2907.595 6.295 2907.765 ;
        RECT 6.585 2907.595 6.755 2907.765 ;
        RECT 2910.105 2907.595 2910.275 2907.765 ;
        RECT 2912.865 2907.595 2913.035 2907.765 ;
        RECT 2913.325 2907.595 2913.495 2907.765 ;
        RECT 2913.785 2907.595 2913.955 2907.765 ;
        RECT 5.665 2902.155 5.835 2902.325 ;
        RECT 6.125 2902.155 6.295 2902.325 ;
        RECT 6.585 2902.155 6.755 2902.325 ;
        RECT 2910.105 2902.155 2910.275 2902.325 ;
        RECT 2912.865 2902.155 2913.035 2902.325 ;
        RECT 2913.325 2902.155 2913.495 2902.325 ;
        RECT 2913.785 2902.155 2913.955 2902.325 ;
        RECT 5.665 2896.715 5.835 2896.885 ;
        RECT 6.125 2896.715 6.295 2896.885 ;
        RECT 6.585 2896.715 6.755 2896.885 ;
        RECT 2910.105 2896.715 2910.275 2896.885 ;
        RECT 2912.865 2896.715 2913.035 2896.885 ;
        RECT 2913.325 2896.715 2913.495 2896.885 ;
        RECT 2913.785 2896.715 2913.955 2896.885 ;
        RECT 5.665 2891.275 5.835 2891.445 ;
        RECT 6.125 2891.275 6.295 2891.445 ;
        RECT 6.585 2891.275 6.755 2891.445 ;
        RECT 2910.105 2891.275 2910.275 2891.445 ;
        RECT 2912.865 2891.275 2913.035 2891.445 ;
        RECT 2913.325 2891.275 2913.495 2891.445 ;
        RECT 2913.785 2891.275 2913.955 2891.445 ;
        RECT 5.665 2885.835 5.835 2886.005 ;
        RECT 6.125 2885.835 6.295 2886.005 ;
        RECT 6.585 2885.835 6.755 2886.005 ;
        RECT 8.885 2885.835 9.055 2886.005 ;
        RECT 9.345 2885.835 9.515 2886.005 ;
        RECT 9.805 2885.835 9.975 2886.005 ;
        RECT 2910.105 2885.835 2910.275 2886.005 ;
        RECT 2912.865 2885.835 2913.035 2886.005 ;
        RECT 2913.325 2885.835 2913.495 2886.005 ;
        RECT 2913.785 2885.835 2913.955 2886.005 ;
        RECT 5.665 2880.395 5.835 2880.565 ;
        RECT 6.125 2880.395 6.295 2880.565 ;
        RECT 6.585 2880.395 6.755 2880.565 ;
        RECT 2910.105 2880.395 2910.275 2880.565 ;
        RECT 2912.865 2880.395 2913.035 2880.565 ;
        RECT 2913.325 2880.395 2913.495 2880.565 ;
        RECT 2913.785 2880.395 2913.955 2880.565 ;
        RECT 5.665 2874.955 5.835 2875.125 ;
        RECT 6.125 2874.955 6.295 2875.125 ;
        RECT 6.585 2874.955 6.755 2875.125 ;
        RECT 2910.105 2874.955 2910.275 2875.125 ;
        RECT 2912.865 2874.955 2913.035 2875.125 ;
        RECT 2913.325 2874.955 2913.495 2875.125 ;
        RECT 2913.785 2874.955 2913.955 2875.125 ;
        RECT 5.665 2869.515 5.835 2869.685 ;
        RECT 6.125 2869.515 6.295 2869.685 ;
        RECT 6.585 2869.515 6.755 2869.685 ;
        RECT 8.885 2869.515 9.055 2869.685 ;
        RECT 9.345 2869.515 9.515 2869.685 ;
        RECT 9.805 2869.515 9.975 2869.685 ;
        RECT 2910.105 2869.515 2910.275 2869.685 ;
        RECT 2912.865 2869.515 2913.035 2869.685 ;
        RECT 2913.325 2869.515 2913.495 2869.685 ;
        RECT 2913.785 2869.515 2913.955 2869.685 ;
        RECT 5.665 2864.075 5.835 2864.245 ;
        RECT 6.125 2864.075 6.295 2864.245 ;
        RECT 6.585 2864.075 6.755 2864.245 ;
        RECT 2910.105 2864.075 2910.275 2864.245 ;
        RECT 2912.865 2864.075 2913.035 2864.245 ;
        RECT 2913.325 2864.075 2913.495 2864.245 ;
        RECT 2913.785 2864.075 2913.955 2864.245 ;
        RECT 5.665 2858.635 5.835 2858.805 ;
        RECT 6.125 2858.635 6.295 2858.805 ;
        RECT 6.585 2858.635 6.755 2858.805 ;
        RECT 2910.105 2858.635 2910.275 2858.805 ;
        RECT 2912.865 2858.635 2913.035 2858.805 ;
        RECT 2913.325 2858.635 2913.495 2858.805 ;
        RECT 2913.785 2858.635 2913.955 2858.805 ;
        RECT 5.665 2853.195 5.835 2853.365 ;
        RECT 6.125 2853.195 6.295 2853.365 ;
        RECT 6.585 2853.195 6.755 2853.365 ;
        RECT 2910.105 2853.195 2910.275 2853.365 ;
        RECT 2912.865 2853.195 2913.035 2853.365 ;
        RECT 2913.325 2853.195 2913.495 2853.365 ;
        RECT 2913.785 2853.195 2913.955 2853.365 ;
        RECT 5.665 2847.755 5.835 2847.925 ;
        RECT 6.125 2847.755 6.295 2847.925 ;
        RECT 6.585 2847.755 6.755 2847.925 ;
        RECT 2910.105 2847.755 2910.275 2847.925 ;
        RECT 2912.865 2847.755 2913.035 2847.925 ;
        RECT 2913.325 2847.755 2913.495 2847.925 ;
        RECT 2913.785 2847.755 2913.955 2847.925 ;
        RECT 5.665 2842.315 5.835 2842.485 ;
        RECT 6.125 2842.315 6.295 2842.485 ;
        RECT 6.585 2842.315 6.755 2842.485 ;
        RECT 2910.105 2842.315 2910.275 2842.485 ;
        RECT 2912.865 2842.315 2913.035 2842.485 ;
        RECT 2913.325 2842.315 2913.495 2842.485 ;
        RECT 2913.785 2842.315 2913.955 2842.485 ;
        RECT 5.665 2836.875 5.835 2837.045 ;
        RECT 6.125 2836.875 6.295 2837.045 ;
        RECT 6.585 2836.875 6.755 2837.045 ;
        RECT 2910.105 2836.875 2910.275 2837.045 ;
        RECT 2912.865 2836.875 2913.035 2837.045 ;
        RECT 2913.325 2836.875 2913.495 2837.045 ;
        RECT 2913.785 2836.875 2913.955 2837.045 ;
        RECT 5.665 2831.435 5.835 2831.605 ;
        RECT 6.125 2831.435 6.295 2831.605 ;
        RECT 6.585 2831.435 6.755 2831.605 ;
        RECT 2910.105 2831.435 2910.275 2831.605 ;
        RECT 2912.865 2831.435 2913.035 2831.605 ;
        RECT 2913.325 2831.435 2913.495 2831.605 ;
        RECT 2913.785 2831.435 2913.955 2831.605 ;
        RECT 5.665 2825.995 5.835 2826.165 ;
        RECT 6.125 2825.995 6.295 2826.165 ;
        RECT 6.585 2825.995 6.755 2826.165 ;
        RECT 2910.105 2825.995 2910.275 2826.165 ;
        RECT 2912.865 2825.995 2913.035 2826.165 ;
        RECT 2913.325 2825.995 2913.495 2826.165 ;
        RECT 2913.785 2825.995 2913.955 2826.165 ;
        RECT 5.665 2820.555 5.835 2820.725 ;
        RECT 6.125 2820.555 6.295 2820.725 ;
        RECT 6.585 2820.555 6.755 2820.725 ;
        RECT 2910.105 2820.555 2910.275 2820.725 ;
        RECT 2912.865 2820.555 2913.035 2820.725 ;
        RECT 2913.325 2820.555 2913.495 2820.725 ;
        RECT 2913.785 2820.555 2913.955 2820.725 ;
        RECT 5.665 2815.115 5.835 2815.285 ;
        RECT 6.125 2815.115 6.295 2815.285 ;
        RECT 6.585 2815.115 6.755 2815.285 ;
        RECT 2910.105 2815.115 2910.275 2815.285 ;
        RECT 2912.865 2815.115 2913.035 2815.285 ;
        RECT 2913.325 2815.115 2913.495 2815.285 ;
        RECT 2913.785 2815.115 2913.955 2815.285 ;
        RECT 5.665 2809.675 5.835 2809.845 ;
        RECT 6.125 2809.675 6.295 2809.845 ;
        RECT 6.585 2809.675 6.755 2809.845 ;
        RECT 2910.105 2809.675 2910.275 2809.845 ;
        RECT 2912.865 2809.675 2913.035 2809.845 ;
        RECT 2913.325 2809.675 2913.495 2809.845 ;
        RECT 2913.785 2809.675 2913.955 2809.845 ;
        RECT 5.665 2804.235 5.835 2804.405 ;
        RECT 6.125 2804.235 6.295 2804.405 ;
        RECT 6.585 2804.235 6.755 2804.405 ;
        RECT 2910.105 2804.235 2910.275 2804.405 ;
        RECT 2912.865 2804.235 2913.035 2804.405 ;
        RECT 2913.325 2804.235 2913.495 2804.405 ;
        RECT 2913.785 2804.235 2913.955 2804.405 ;
        RECT 5.665 2798.795 5.835 2798.965 ;
        RECT 6.125 2798.795 6.295 2798.965 ;
        RECT 6.585 2798.795 6.755 2798.965 ;
        RECT 2910.105 2798.795 2910.275 2798.965 ;
        RECT 2912.865 2798.795 2913.035 2798.965 ;
        RECT 2913.325 2798.795 2913.495 2798.965 ;
        RECT 2913.785 2798.795 2913.955 2798.965 ;
        RECT 5.665 2793.355 5.835 2793.525 ;
        RECT 6.125 2793.355 6.295 2793.525 ;
        RECT 6.585 2793.355 6.755 2793.525 ;
        RECT 2910.105 2793.355 2910.275 2793.525 ;
        RECT 2912.865 2793.355 2913.035 2793.525 ;
        RECT 2913.325 2793.355 2913.495 2793.525 ;
        RECT 2913.785 2793.355 2913.955 2793.525 ;
        RECT 5.665 2787.915 5.835 2788.085 ;
        RECT 6.125 2787.915 6.295 2788.085 ;
        RECT 6.585 2787.915 6.755 2788.085 ;
        RECT 2910.105 2787.915 2910.275 2788.085 ;
        RECT 2912.865 2787.915 2913.035 2788.085 ;
        RECT 2913.325 2787.915 2913.495 2788.085 ;
        RECT 2913.785 2787.915 2913.955 2788.085 ;
        RECT 5.665 2782.475 5.835 2782.645 ;
        RECT 6.125 2782.475 6.295 2782.645 ;
        RECT 6.585 2782.475 6.755 2782.645 ;
        RECT 2910.105 2782.475 2910.275 2782.645 ;
        RECT 2912.865 2782.475 2913.035 2782.645 ;
        RECT 2913.325 2782.475 2913.495 2782.645 ;
        RECT 2913.785 2782.475 2913.955 2782.645 ;
        RECT 5.665 2777.035 5.835 2777.205 ;
        RECT 6.125 2777.035 6.295 2777.205 ;
        RECT 6.585 2777.035 6.755 2777.205 ;
        RECT 2909.185 2777.035 2909.355 2777.205 ;
        RECT 2909.645 2777.035 2909.815 2777.205 ;
        RECT 2910.105 2777.035 2910.275 2777.205 ;
        RECT 2912.865 2777.035 2913.035 2777.205 ;
        RECT 2913.325 2777.035 2913.495 2777.205 ;
        RECT 2913.785 2777.035 2913.955 2777.205 ;
        RECT 5.665 2771.595 5.835 2771.765 ;
        RECT 6.125 2771.595 6.295 2771.765 ;
        RECT 6.585 2771.595 6.755 2771.765 ;
        RECT 2910.105 2771.595 2910.275 2771.765 ;
        RECT 2912.865 2771.595 2913.035 2771.765 ;
        RECT 2913.325 2771.595 2913.495 2771.765 ;
        RECT 2913.785 2771.595 2913.955 2771.765 ;
        RECT 5.665 2766.155 5.835 2766.325 ;
        RECT 6.125 2766.155 6.295 2766.325 ;
        RECT 6.585 2766.155 6.755 2766.325 ;
        RECT 2910.105 2766.155 2910.275 2766.325 ;
        RECT 2912.865 2766.155 2913.035 2766.325 ;
        RECT 2913.325 2766.155 2913.495 2766.325 ;
        RECT 2913.785 2766.155 2913.955 2766.325 ;
        RECT 5.665 2760.715 5.835 2760.885 ;
        RECT 6.125 2760.715 6.295 2760.885 ;
        RECT 6.585 2760.715 6.755 2760.885 ;
        RECT 2910.105 2760.715 2910.275 2760.885 ;
        RECT 2912.865 2760.715 2913.035 2760.885 ;
        RECT 2913.325 2760.715 2913.495 2760.885 ;
        RECT 2913.785 2760.715 2913.955 2760.885 ;
        RECT 5.665 2755.275 5.835 2755.445 ;
        RECT 6.125 2755.275 6.295 2755.445 ;
        RECT 6.585 2755.275 6.755 2755.445 ;
        RECT 2910.105 2755.275 2910.275 2755.445 ;
        RECT 2912.865 2755.275 2913.035 2755.445 ;
        RECT 2913.325 2755.275 2913.495 2755.445 ;
        RECT 2913.785 2755.275 2913.955 2755.445 ;
        RECT 5.665 2749.835 5.835 2750.005 ;
        RECT 6.125 2749.835 6.295 2750.005 ;
        RECT 6.585 2749.835 6.755 2750.005 ;
        RECT 2910.105 2749.835 2910.275 2750.005 ;
        RECT 2912.865 2749.835 2913.035 2750.005 ;
        RECT 2913.325 2749.835 2913.495 2750.005 ;
        RECT 2913.785 2749.835 2913.955 2750.005 ;
        RECT 5.665 2744.395 5.835 2744.565 ;
        RECT 6.125 2744.395 6.295 2744.565 ;
        RECT 6.585 2744.395 6.755 2744.565 ;
        RECT 2910.105 2744.395 2910.275 2744.565 ;
        RECT 2912.865 2744.395 2913.035 2744.565 ;
        RECT 2913.325 2744.395 2913.495 2744.565 ;
        RECT 2913.785 2744.395 2913.955 2744.565 ;
        RECT 5.665 2738.955 5.835 2739.125 ;
        RECT 6.125 2738.955 6.295 2739.125 ;
        RECT 6.585 2738.955 6.755 2739.125 ;
        RECT 2910.105 2738.955 2910.275 2739.125 ;
        RECT 2912.865 2738.955 2913.035 2739.125 ;
        RECT 2913.325 2738.955 2913.495 2739.125 ;
        RECT 2913.785 2738.955 2913.955 2739.125 ;
        RECT 5.665 2733.515 5.835 2733.685 ;
        RECT 6.125 2733.515 6.295 2733.685 ;
        RECT 6.585 2733.515 6.755 2733.685 ;
        RECT 2910.105 2733.515 2910.275 2733.685 ;
        RECT 2912.865 2733.515 2913.035 2733.685 ;
        RECT 2913.325 2733.515 2913.495 2733.685 ;
        RECT 2913.785 2733.515 2913.955 2733.685 ;
        RECT 5.665 2728.075 5.835 2728.245 ;
        RECT 6.125 2728.075 6.295 2728.245 ;
        RECT 6.585 2728.075 6.755 2728.245 ;
        RECT 2910.105 2728.075 2910.275 2728.245 ;
        RECT 2912.865 2728.075 2913.035 2728.245 ;
        RECT 2913.325 2728.075 2913.495 2728.245 ;
        RECT 2913.785 2728.075 2913.955 2728.245 ;
        RECT 5.665 2722.635 5.835 2722.805 ;
        RECT 6.125 2722.635 6.295 2722.805 ;
        RECT 6.585 2722.635 6.755 2722.805 ;
        RECT 2910.105 2722.635 2910.275 2722.805 ;
        RECT 2912.865 2722.635 2913.035 2722.805 ;
        RECT 2913.325 2722.635 2913.495 2722.805 ;
        RECT 2913.785 2722.635 2913.955 2722.805 ;
        RECT 5.665 2717.195 5.835 2717.365 ;
        RECT 6.125 2717.195 6.295 2717.365 ;
        RECT 6.585 2717.195 6.755 2717.365 ;
        RECT 2910.105 2717.195 2910.275 2717.365 ;
        RECT 2912.865 2717.195 2913.035 2717.365 ;
        RECT 2913.325 2717.195 2913.495 2717.365 ;
        RECT 2913.785 2717.195 2913.955 2717.365 ;
        RECT 5.665 2711.755 5.835 2711.925 ;
        RECT 6.125 2711.755 6.295 2711.925 ;
        RECT 6.585 2711.755 6.755 2711.925 ;
        RECT 2910.105 2711.755 2910.275 2711.925 ;
        RECT 2912.865 2711.755 2913.035 2711.925 ;
        RECT 2913.325 2711.755 2913.495 2711.925 ;
        RECT 2913.785 2711.755 2913.955 2711.925 ;
        RECT 5.665 2706.315 5.835 2706.485 ;
        RECT 6.125 2706.315 6.295 2706.485 ;
        RECT 6.585 2706.315 6.755 2706.485 ;
        RECT 2910.105 2706.315 2910.275 2706.485 ;
        RECT 2912.865 2706.315 2913.035 2706.485 ;
        RECT 2913.325 2706.315 2913.495 2706.485 ;
        RECT 2913.785 2706.315 2913.955 2706.485 ;
        RECT 5.665 2700.875 5.835 2701.045 ;
        RECT 6.125 2700.875 6.295 2701.045 ;
        RECT 6.585 2700.875 6.755 2701.045 ;
        RECT 2910.105 2700.875 2910.275 2701.045 ;
        RECT 2912.865 2700.875 2913.035 2701.045 ;
        RECT 2913.325 2700.875 2913.495 2701.045 ;
        RECT 2913.785 2700.875 2913.955 2701.045 ;
        RECT 5.665 2695.435 5.835 2695.605 ;
        RECT 6.125 2695.435 6.295 2695.605 ;
        RECT 6.585 2695.435 6.755 2695.605 ;
        RECT 2910.105 2695.435 2910.275 2695.605 ;
        RECT 2912.865 2695.435 2913.035 2695.605 ;
        RECT 2913.325 2695.435 2913.495 2695.605 ;
        RECT 2913.785 2695.435 2913.955 2695.605 ;
        RECT 5.665 2689.995 5.835 2690.165 ;
        RECT 6.125 2689.995 6.295 2690.165 ;
        RECT 6.585 2689.995 6.755 2690.165 ;
        RECT 2906.425 2689.995 2906.595 2690.165 ;
        RECT 2912.865 2689.995 2913.035 2690.165 ;
        RECT 2913.325 2689.995 2913.495 2690.165 ;
        RECT 2913.785 2689.995 2913.955 2690.165 ;
        RECT 5.665 2684.555 5.835 2684.725 ;
        RECT 6.125 2684.555 6.295 2684.725 ;
        RECT 6.585 2684.555 6.755 2684.725 ;
        RECT 2906.425 2684.555 2906.595 2684.725 ;
        RECT 2912.865 2684.555 2913.035 2684.725 ;
        RECT 2913.325 2684.555 2913.495 2684.725 ;
        RECT 2913.785 2684.555 2913.955 2684.725 ;
        RECT 5.665 2679.115 5.835 2679.285 ;
        RECT 6.125 2679.115 6.295 2679.285 ;
        RECT 6.585 2679.115 6.755 2679.285 ;
        RECT 2906.425 2679.115 2906.595 2679.285 ;
        RECT 2912.865 2679.115 2913.035 2679.285 ;
        RECT 2913.325 2679.115 2913.495 2679.285 ;
        RECT 2913.785 2679.115 2913.955 2679.285 ;
        RECT 5.665 2673.675 5.835 2673.845 ;
        RECT 6.125 2673.675 6.295 2673.845 ;
        RECT 6.585 2673.675 6.755 2673.845 ;
        RECT 2906.425 2673.675 2906.595 2673.845 ;
        RECT 2912.865 2673.675 2913.035 2673.845 ;
        RECT 2913.325 2673.675 2913.495 2673.845 ;
        RECT 2913.785 2673.675 2913.955 2673.845 ;
        RECT 5.665 2668.235 5.835 2668.405 ;
        RECT 6.125 2668.235 6.295 2668.405 ;
        RECT 6.585 2668.235 6.755 2668.405 ;
        RECT 2906.425 2668.235 2906.595 2668.405 ;
        RECT 2912.865 2668.235 2913.035 2668.405 ;
        RECT 2913.325 2668.235 2913.495 2668.405 ;
        RECT 2913.785 2668.235 2913.955 2668.405 ;
        RECT 5.665 2662.795 5.835 2662.965 ;
        RECT 6.125 2662.795 6.295 2662.965 ;
        RECT 6.585 2662.795 6.755 2662.965 ;
        RECT 2906.425 2662.795 2906.595 2662.965 ;
        RECT 2912.865 2662.795 2913.035 2662.965 ;
        RECT 2913.325 2662.795 2913.495 2662.965 ;
        RECT 2913.785 2662.795 2913.955 2662.965 ;
        RECT 5.665 2657.355 5.835 2657.525 ;
        RECT 6.125 2657.355 6.295 2657.525 ;
        RECT 6.585 2657.355 6.755 2657.525 ;
        RECT 2906.425 2657.355 2906.595 2657.525 ;
        RECT 2912.865 2657.355 2913.035 2657.525 ;
        RECT 2913.325 2657.355 2913.495 2657.525 ;
        RECT 2913.785 2657.355 2913.955 2657.525 ;
        RECT 5.665 2651.915 5.835 2652.085 ;
        RECT 6.125 2651.915 6.295 2652.085 ;
        RECT 6.585 2651.915 6.755 2652.085 ;
        RECT 2906.425 2651.915 2906.595 2652.085 ;
        RECT 2912.865 2651.915 2913.035 2652.085 ;
        RECT 2913.325 2651.915 2913.495 2652.085 ;
        RECT 2913.785 2651.915 2913.955 2652.085 ;
        RECT 5.665 2646.475 5.835 2646.645 ;
        RECT 6.125 2646.475 6.295 2646.645 ;
        RECT 6.585 2646.475 6.755 2646.645 ;
        RECT 2906.425 2646.475 2906.595 2646.645 ;
        RECT 2912.865 2646.475 2913.035 2646.645 ;
        RECT 2913.325 2646.475 2913.495 2646.645 ;
        RECT 2913.785 2646.475 2913.955 2646.645 ;
        RECT 5.665 2641.035 5.835 2641.205 ;
        RECT 6.125 2641.035 6.295 2641.205 ;
        RECT 6.585 2641.035 6.755 2641.205 ;
        RECT 2906.425 2641.035 2906.595 2641.205 ;
        RECT 2912.865 2641.035 2913.035 2641.205 ;
        RECT 2913.325 2641.035 2913.495 2641.205 ;
        RECT 2913.785 2641.035 2913.955 2641.205 ;
        RECT 5.665 2635.595 5.835 2635.765 ;
        RECT 6.125 2635.595 6.295 2635.765 ;
        RECT 6.585 2635.595 6.755 2635.765 ;
        RECT 2906.425 2635.595 2906.595 2635.765 ;
        RECT 2912.865 2635.595 2913.035 2635.765 ;
        RECT 2913.325 2635.595 2913.495 2635.765 ;
        RECT 2913.785 2635.595 2913.955 2635.765 ;
        RECT 5.665 2630.155 5.835 2630.325 ;
        RECT 6.125 2630.155 6.295 2630.325 ;
        RECT 6.585 2630.155 6.755 2630.325 ;
        RECT 2906.425 2630.155 2906.595 2630.325 ;
        RECT 2909.185 2630.155 2909.355 2630.325 ;
        RECT 2909.645 2630.155 2909.815 2630.325 ;
        RECT 2910.105 2630.155 2910.275 2630.325 ;
        RECT 2912.865 2630.155 2913.035 2630.325 ;
        RECT 2913.325 2630.155 2913.495 2630.325 ;
        RECT 2913.785 2630.155 2913.955 2630.325 ;
        RECT 5.665 2624.715 5.835 2624.885 ;
        RECT 6.125 2624.715 6.295 2624.885 ;
        RECT 6.585 2624.715 6.755 2624.885 ;
        RECT 2906.425 2624.715 2906.595 2624.885 ;
        RECT 2912.865 2624.715 2913.035 2624.885 ;
        RECT 2913.325 2624.715 2913.495 2624.885 ;
        RECT 2913.785 2624.715 2913.955 2624.885 ;
        RECT 5.665 2619.275 5.835 2619.445 ;
        RECT 6.125 2619.275 6.295 2619.445 ;
        RECT 6.585 2619.275 6.755 2619.445 ;
        RECT 2906.425 2619.275 2906.595 2619.445 ;
        RECT 2912.865 2619.275 2913.035 2619.445 ;
        RECT 2913.325 2619.275 2913.495 2619.445 ;
        RECT 2913.785 2619.275 2913.955 2619.445 ;
        RECT 5.665 2613.835 5.835 2614.005 ;
        RECT 6.125 2613.835 6.295 2614.005 ;
        RECT 6.585 2613.835 6.755 2614.005 ;
        RECT 2906.425 2613.835 2906.595 2614.005 ;
        RECT 2912.865 2613.835 2913.035 2614.005 ;
        RECT 2913.325 2613.835 2913.495 2614.005 ;
        RECT 2913.785 2613.835 2913.955 2614.005 ;
        RECT 5.665 2608.395 5.835 2608.565 ;
        RECT 6.125 2608.395 6.295 2608.565 ;
        RECT 6.585 2608.395 6.755 2608.565 ;
        RECT 2906.425 2608.395 2906.595 2608.565 ;
        RECT 2912.865 2608.395 2913.035 2608.565 ;
        RECT 2913.325 2608.395 2913.495 2608.565 ;
        RECT 2913.785 2608.395 2913.955 2608.565 ;
        RECT 5.665 2602.955 5.835 2603.125 ;
        RECT 6.125 2602.955 6.295 2603.125 ;
        RECT 6.585 2602.955 6.755 2603.125 ;
        RECT 2906.425 2602.955 2906.595 2603.125 ;
        RECT 2909.185 2602.955 2909.355 2603.125 ;
        RECT 2909.645 2602.955 2909.815 2603.125 ;
        RECT 2910.105 2602.955 2910.275 2603.125 ;
        RECT 2912.865 2602.955 2913.035 2603.125 ;
        RECT 2913.325 2602.955 2913.495 2603.125 ;
        RECT 2913.785 2602.955 2913.955 2603.125 ;
        RECT 5.665 2597.515 5.835 2597.685 ;
        RECT 6.125 2597.515 6.295 2597.685 ;
        RECT 6.585 2597.515 6.755 2597.685 ;
        RECT 2906.425 2597.515 2906.595 2597.685 ;
        RECT 2912.865 2597.515 2913.035 2597.685 ;
        RECT 2913.325 2597.515 2913.495 2597.685 ;
        RECT 2913.785 2597.515 2913.955 2597.685 ;
        RECT 5.665 2592.075 5.835 2592.245 ;
        RECT 6.125 2592.075 6.295 2592.245 ;
        RECT 6.585 2592.075 6.755 2592.245 ;
        RECT 2906.425 2592.075 2906.595 2592.245 ;
        RECT 2912.865 2592.075 2913.035 2592.245 ;
        RECT 2913.325 2592.075 2913.495 2592.245 ;
        RECT 2913.785 2592.075 2913.955 2592.245 ;
        RECT 5.665 2586.635 5.835 2586.805 ;
        RECT 6.125 2586.635 6.295 2586.805 ;
        RECT 6.585 2586.635 6.755 2586.805 ;
        RECT 2906.425 2586.635 2906.595 2586.805 ;
        RECT 2912.865 2586.635 2913.035 2586.805 ;
        RECT 2913.325 2586.635 2913.495 2586.805 ;
        RECT 2913.785 2586.635 2913.955 2586.805 ;
        RECT 5.665 2581.195 5.835 2581.365 ;
        RECT 6.125 2581.195 6.295 2581.365 ;
        RECT 6.585 2581.195 6.755 2581.365 ;
        RECT 2906.425 2581.195 2906.595 2581.365 ;
        RECT 2912.865 2581.195 2913.035 2581.365 ;
        RECT 2913.325 2581.195 2913.495 2581.365 ;
        RECT 2913.785 2581.195 2913.955 2581.365 ;
        RECT 5.665 2575.755 5.835 2575.925 ;
        RECT 6.125 2575.755 6.295 2575.925 ;
        RECT 6.585 2575.755 6.755 2575.925 ;
        RECT 2906.425 2575.755 2906.595 2575.925 ;
        RECT 2912.865 2575.755 2913.035 2575.925 ;
        RECT 2913.325 2575.755 2913.495 2575.925 ;
        RECT 2913.785 2575.755 2913.955 2575.925 ;
        RECT 5.665 2570.315 5.835 2570.485 ;
        RECT 6.125 2570.315 6.295 2570.485 ;
        RECT 6.585 2570.315 6.755 2570.485 ;
        RECT 2906.425 2570.315 2906.595 2570.485 ;
        RECT 2912.865 2570.315 2913.035 2570.485 ;
        RECT 2913.325 2570.315 2913.495 2570.485 ;
        RECT 2913.785 2570.315 2913.955 2570.485 ;
        RECT 5.665 2564.875 5.835 2565.045 ;
        RECT 6.125 2564.875 6.295 2565.045 ;
        RECT 6.585 2564.875 6.755 2565.045 ;
        RECT 2906.425 2564.875 2906.595 2565.045 ;
        RECT 2912.865 2564.875 2913.035 2565.045 ;
        RECT 2913.325 2564.875 2913.495 2565.045 ;
        RECT 2913.785 2564.875 2913.955 2565.045 ;
        RECT 5.665 2559.435 5.835 2559.605 ;
        RECT 6.125 2559.435 6.295 2559.605 ;
        RECT 6.585 2559.435 6.755 2559.605 ;
        RECT 2906.425 2559.435 2906.595 2559.605 ;
        RECT 2912.865 2559.435 2913.035 2559.605 ;
        RECT 2913.325 2559.435 2913.495 2559.605 ;
        RECT 2913.785 2559.435 2913.955 2559.605 ;
        RECT 5.665 2553.995 5.835 2554.165 ;
        RECT 6.125 2553.995 6.295 2554.165 ;
        RECT 6.585 2553.995 6.755 2554.165 ;
        RECT 2906.425 2553.995 2906.595 2554.165 ;
        RECT 2912.865 2553.995 2913.035 2554.165 ;
        RECT 2913.325 2553.995 2913.495 2554.165 ;
        RECT 2913.785 2553.995 2913.955 2554.165 ;
        RECT 5.665 2548.555 5.835 2548.725 ;
        RECT 6.125 2548.555 6.295 2548.725 ;
        RECT 6.585 2548.555 6.755 2548.725 ;
        RECT 2906.425 2548.555 2906.595 2548.725 ;
        RECT 2912.865 2548.555 2913.035 2548.725 ;
        RECT 2913.325 2548.555 2913.495 2548.725 ;
        RECT 2913.785 2548.555 2913.955 2548.725 ;
        RECT 5.665 2543.115 5.835 2543.285 ;
        RECT 6.125 2543.115 6.295 2543.285 ;
        RECT 6.585 2543.115 6.755 2543.285 ;
        RECT 2906.425 2543.115 2906.595 2543.285 ;
        RECT 2912.865 2543.115 2913.035 2543.285 ;
        RECT 2913.325 2543.115 2913.495 2543.285 ;
        RECT 2913.785 2543.115 2913.955 2543.285 ;
        RECT 5.665 2537.675 5.835 2537.845 ;
        RECT 6.125 2537.675 6.295 2537.845 ;
        RECT 6.585 2537.675 6.755 2537.845 ;
        RECT 2906.425 2537.675 2906.595 2537.845 ;
        RECT 2912.865 2537.675 2913.035 2537.845 ;
        RECT 2913.325 2537.675 2913.495 2537.845 ;
        RECT 2913.785 2537.675 2913.955 2537.845 ;
        RECT 5.665 2532.235 5.835 2532.405 ;
        RECT 6.125 2532.235 6.295 2532.405 ;
        RECT 6.585 2532.235 6.755 2532.405 ;
        RECT 2906.425 2532.235 2906.595 2532.405 ;
        RECT 2912.865 2532.235 2913.035 2532.405 ;
        RECT 2913.325 2532.235 2913.495 2532.405 ;
        RECT 2913.785 2532.235 2913.955 2532.405 ;
        RECT 5.665 2526.795 5.835 2526.965 ;
        RECT 6.125 2526.795 6.295 2526.965 ;
        RECT 6.585 2526.795 6.755 2526.965 ;
        RECT 2906.425 2526.795 2906.595 2526.965 ;
        RECT 2912.865 2526.795 2913.035 2526.965 ;
        RECT 2913.325 2526.795 2913.495 2526.965 ;
        RECT 2913.785 2526.795 2913.955 2526.965 ;
        RECT 5.665 2521.355 5.835 2521.525 ;
        RECT 6.125 2521.355 6.295 2521.525 ;
        RECT 6.585 2521.355 6.755 2521.525 ;
        RECT 2906.425 2521.355 2906.595 2521.525 ;
        RECT 2912.865 2521.355 2913.035 2521.525 ;
        RECT 2913.325 2521.355 2913.495 2521.525 ;
        RECT 2913.785 2521.355 2913.955 2521.525 ;
        RECT 5.665 2515.915 5.835 2516.085 ;
        RECT 6.125 2515.915 6.295 2516.085 ;
        RECT 6.585 2515.915 6.755 2516.085 ;
        RECT 2906.425 2515.915 2906.595 2516.085 ;
        RECT 2912.865 2515.915 2913.035 2516.085 ;
        RECT 2913.325 2515.915 2913.495 2516.085 ;
        RECT 2913.785 2515.915 2913.955 2516.085 ;
        RECT 5.665 2510.475 5.835 2510.645 ;
        RECT 6.125 2510.475 6.295 2510.645 ;
        RECT 6.585 2510.475 6.755 2510.645 ;
        RECT 2906.425 2510.475 2906.595 2510.645 ;
        RECT 2912.865 2510.475 2913.035 2510.645 ;
        RECT 2913.325 2510.475 2913.495 2510.645 ;
        RECT 2913.785 2510.475 2913.955 2510.645 ;
        RECT 5.665 2505.035 5.835 2505.205 ;
        RECT 6.125 2505.035 6.295 2505.205 ;
        RECT 6.585 2505.035 6.755 2505.205 ;
        RECT 2906.425 2505.035 2906.595 2505.205 ;
        RECT 2912.865 2505.035 2913.035 2505.205 ;
        RECT 2913.325 2505.035 2913.495 2505.205 ;
        RECT 2913.785 2505.035 2913.955 2505.205 ;
        RECT 5.665 2499.595 5.835 2499.765 ;
        RECT 6.125 2499.595 6.295 2499.765 ;
        RECT 6.585 2499.595 6.755 2499.765 ;
        RECT 8.885 2499.595 9.055 2499.765 ;
        RECT 9.345 2499.595 9.515 2499.765 ;
        RECT 9.805 2499.595 9.975 2499.765 ;
        RECT 2906.425 2499.595 2906.595 2499.765 ;
        RECT 2912.865 2499.595 2913.035 2499.765 ;
        RECT 2913.325 2499.595 2913.495 2499.765 ;
        RECT 2913.785 2499.595 2913.955 2499.765 ;
        RECT 5.665 2494.155 5.835 2494.325 ;
        RECT 6.125 2494.155 6.295 2494.325 ;
        RECT 6.585 2494.155 6.755 2494.325 ;
        RECT 2906.425 2494.155 2906.595 2494.325 ;
        RECT 2912.865 2494.155 2913.035 2494.325 ;
        RECT 2913.325 2494.155 2913.495 2494.325 ;
        RECT 2913.785 2494.155 2913.955 2494.325 ;
        RECT 5.665 2488.715 5.835 2488.885 ;
        RECT 6.125 2488.715 6.295 2488.885 ;
        RECT 6.585 2488.715 6.755 2488.885 ;
        RECT 2906.425 2488.715 2906.595 2488.885 ;
        RECT 2912.865 2488.715 2913.035 2488.885 ;
        RECT 2913.325 2488.715 2913.495 2488.885 ;
        RECT 2913.785 2488.715 2913.955 2488.885 ;
        RECT 5.665 2483.275 5.835 2483.445 ;
        RECT 6.125 2483.275 6.295 2483.445 ;
        RECT 6.585 2483.275 6.755 2483.445 ;
        RECT 2906.425 2483.275 2906.595 2483.445 ;
        RECT 2912.865 2483.275 2913.035 2483.445 ;
        RECT 2913.325 2483.275 2913.495 2483.445 ;
        RECT 2913.785 2483.275 2913.955 2483.445 ;
        RECT 5.665 2477.835 5.835 2478.005 ;
        RECT 6.125 2477.835 6.295 2478.005 ;
        RECT 6.585 2477.835 6.755 2478.005 ;
        RECT 2906.425 2477.835 2906.595 2478.005 ;
        RECT 2912.865 2477.835 2913.035 2478.005 ;
        RECT 2913.325 2477.835 2913.495 2478.005 ;
        RECT 2913.785 2477.835 2913.955 2478.005 ;
        RECT 5.665 2472.395 5.835 2472.565 ;
        RECT 6.125 2472.395 6.295 2472.565 ;
        RECT 6.585 2472.395 6.755 2472.565 ;
        RECT 2906.425 2472.395 2906.595 2472.565 ;
        RECT 2912.865 2472.395 2913.035 2472.565 ;
        RECT 2913.325 2472.395 2913.495 2472.565 ;
        RECT 2913.785 2472.395 2913.955 2472.565 ;
        RECT 5.665 2466.955 5.835 2467.125 ;
        RECT 6.125 2466.955 6.295 2467.125 ;
        RECT 6.585 2466.955 6.755 2467.125 ;
        RECT 2906.425 2466.955 2906.595 2467.125 ;
        RECT 2912.865 2466.955 2913.035 2467.125 ;
        RECT 2913.325 2466.955 2913.495 2467.125 ;
        RECT 2913.785 2466.955 2913.955 2467.125 ;
        RECT 5.665 2461.515 5.835 2461.685 ;
        RECT 6.125 2461.515 6.295 2461.685 ;
        RECT 6.585 2461.515 6.755 2461.685 ;
        RECT 2906.425 2461.515 2906.595 2461.685 ;
        RECT 2909.185 2461.515 2909.355 2461.685 ;
        RECT 2909.645 2461.515 2909.815 2461.685 ;
        RECT 2910.105 2461.515 2910.275 2461.685 ;
        RECT 2912.865 2461.515 2913.035 2461.685 ;
        RECT 2913.325 2461.515 2913.495 2461.685 ;
        RECT 2913.785 2461.515 2913.955 2461.685 ;
        RECT 5.665 2456.075 5.835 2456.245 ;
        RECT 6.125 2456.075 6.295 2456.245 ;
        RECT 6.585 2456.075 6.755 2456.245 ;
        RECT 2906.425 2456.075 2906.595 2456.245 ;
        RECT 2912.865 2456.075 2913.035 2456.245 ;
        RECT 2913.325 2456.075 2913.495 2456.245 ;
        RECT 2913.785 2456.075 2913.955 2456.245 ;
        RECT 5.665 2450.635 5.835 2450.805 ;
        RECT 6.125 2450.635 6.295 2450.805 ;
        RECT 6.585 2450.635 6.755 2450.805 ;
        RECT 2906.425 2450.635 2906.595 2450.805 ;
        RECT 2912.865 2450.635 2913.035 2450.805 ;
        RECT 2913.325 2450.635 2913.495 2450.805 ;
        RECT 2913.785 2450.635 2913.955 2450.805 ;
        RECT 5.665 2445.195 5.835 2445.365 ;
        RECT 6.125 2445.195 6.295 2445.365 ;
        RECT 6.585 2445.195 6.755 2445.365 ;
        RECT 2906.425 2445.195 2906.595 2445.365 ;
        RECT 2912.865 2445.195 2913.035 2445.365 ;
        RECT 2913.325 2445.195 2913.495 2445.365 ;
        RECT 2913.785 2445.195 2913.955 2445.365 ;
        RECT 5.665 2439.755 5.835 2439.925 ;
        RECT 6.125 2439.755 6.295 2439.925 ;
        RECT 6.585 2439.755 6.755 2439.925 ;
        RECT 2906.425 2439.755 2906.595 2439.925 ;
        RECT 2912.865 2439.755 2913.035 2439.925 ;
        RECT 2913.325 2439.755 2913.495 2439.925 ;
        RECT 2913.785 2439.755 2913.955 2439.925 ;
        RECT 5.665 2434.315 5.835 2434.485 ;
        RECT 6.125 2434.315 6.295 2434.485 ;
        RECT 6.585 2434.315 6.755 2434.485 ;
        RECT 2906.425 2434.315 2906.595 2434.485 ;
        RECT 2909.185 2434.315 2909.355 2434.485 ;
        RECT 2909.645 2434.315 2909.815 2434.485 ;
        RECT 2910.105 2434.315 2910.275 2434.485 ;
        RECT 2912.865 2434.315 2913.035 2434.485 ;
        RECT 2913.325 2434.315 2913.495 2434.485 ;
        RECT 2913.785 2434.315 2913.955 2434.485 ;
        RECT 5.665 2428.875 5.835 2429.045 ;
        RECT 6.125 2428.875 6.295 2429.045 ;
        RECT 6.585 2428.875 6.755 2429.045 ;
        RECT 2906.425 2428.875 2906.595 2429.045 ;
        RECT 2912.865 2428.875 2913.035 2429.045 ;
        RECT 2913.325 2428.875 2913.495 2429.045 ;
        RECT 2913.785 2428.875 2913.955 2429.045 ;
        RECT 5.665 2423.435 5.835 2423.605 ;
        RECT 6.125 2423.435 6.295 2423.605 ;
        RECT 6.585 2423.435 6.755 2423.605 ;
        RECT 2906.425 2423.435 2906.595 2423.605 ;
        RECT 2912.865 2423.435 2913.035 2423.605 ;
        RECT 2913.325 2423.435 2913.495 2423.605 ;
        RECT 2913.785 2423.435 2913.955 2423.605 ;
        RECT 5.665 2417.995 5.835 2418.165 ;
        RECT 6.125 2417.995 6.295 2418.165 ;
        RECT 6.585 2417.995 6.755 2418.165 ;
        RECT 2906.425 2417.995 2906.595 2418.165 ;
        RECT 2912.865 2417.995 2913.035 2418.165 ;
        RECT 2913.325 2417.995 2913.495 2418.165 ;
        RECT 2913.785 2417.995 2913.955 2418.165 ;
        RECT 5.665 2412.555 5.835 2412.725 ;
        RECT 6.125 2412.555 6.295 2412.725 ;
        RECT 6.585 2412.555 6.755 2412.725 ;
        RECT 2906.425 2412.555 2906.595 2412.725 ;
        RECT 2912.865 2412.555 2913.035 2412.725 ;
        RECT 2913.325 2412.555 2913.495 2412.725 ;
        RECT 2913.785 2412.555 2913.955 2412.725 ;
        RECT 5.665 2407.115 5.835 2407.285 ;
        RECT 6.125 2407.115 6.295 2407.285 ;
        RECT 6.585 2407.115 6.755 2407.285 ;
        RECT 2906.425 2407.115 2906.595 2407.285 ;
        RECT 2912.865 2407.115 2913.035 2407.285 ;
        RECT 2913.325 2407.115 2913.495 2407.285 ;
        RECT 2913.785 2407.115 2913.955 2407.285 ;
        RECT 5.665 2401.675 5.835 2401.845 ;
        RECT 6.125 2401.675 6.295 2401.845 ;
        RECT 6.585 2401.675 6.755 2401.845 ;
        RECT 2906.425 2401.675 2906.595 2401.845 ;
        RECT 2912.865 2401.675 2913.035 2401.845 ;
        RECT 2913.325 2401.675 2913.495 2401.845 ;
        RECT 2913.785 2401.675 2913.955 2401.845 ;
        RECT 5.665 2396.235 5.835 2396.405 ;
        RECT 6.125 2396.235 6.295 2396.405 ;
        RECT 6.585 2396.235 6.755 2396.405 ;
        RECT 2906.425 2396.235 2906.595 2396.405 ;
        RECT 2912.865 2396.235 2913.035 2396.405 ;
        RECT 2913.325 2396.235 2913.495 2396.405 ;
        RECT 2913.785 2396.235 2913.955 2396.405 ;
        RECT 5.665 2390.795 5.835 2390.965 ;
        RECT 6.125 2390.795 6.295 2390.965 ;
        RECT 6.585 2390.795 6.755 2390.965 ;
        RECT 2906.425 2390.795 2906.595 2390.965 ;
        RECT 2912.865 2390.795 2913.035 2390.965 ;
        RECT 2913.325 2390.795 2913.495 2390.965 ;
        RECT 2913.785 2390.795 2913.955 2390.965 ;
        RECT 5.665 2385.355 5.835 2385.525 ;
        RECT 6.125 2385.355 6.295 2385.525 ;
        RECT 6.585 2385.355 6.755 2385.525 ;
        RECT 2906.425 2385.355 2906.595 2385.525 ;
        RECT 2909.185 2385.355 2909.355 2385.525 ;
        RECT 2909.645 2385.355 2909.815 2385.525 ;
        RECT 2910.105 2385.355 2910.275 2385.525 ;
        RECT 2912.865 2385.355 2913.035 2385.525 ;
        RECT 2913.325 2385.355 2913.495 2385.525 ;
        RECT 2913.785 2385.355 2913.955 2385.525 ;
        RECT 5.665 2379.915 5.835 2380.085 ;
        RECT 6.125 2379.915 6.295 2380.085 ;
        RECT 6.585 2379.915 6.755 2380.085 ;
        RECT 8.885 2379.915 9.055 2380.085 ;
        RECT 9.345 2379.915 9.515 2380.085 ;
        RECT 9.805 2379.915 9.975 2380.085 ;
        RECT 2906.425 2379.915 2906.595 2380.085 ;
        RECT 2912.865 2379.915 2913.035 2380.085 ;
        RECT 2913.325 2379.915 2913.495 2380.085 ;
        RECT 2913.785 2379.915 2913.955 2380.085 ;
        RECT 5.665 2374.475 5.835 2374.645 ;
        RECT 6.125 2374.475 6.295 2374.645 ;
        RECT 6.585 2374.475 6.755 2374.645 ;
        RECT 2906.425 2374.475 2906.595 2374.645 ;
        RECT 2912.865 2374.475 2913.035 2374.645 ;
        RECT 2913.325 2374.475 2913.495 2374.645 ;
        RECT 2913.785 2374.475 2913.955 2374.645 ;
        RECT 5.665 2369.035 5.835 2369.205 ;
        RECT 6.125 2369.035 6.295 2369.205 ;
        RECT 6.585 2369.035 6.755 2369.205 ;
        RECT 2906.425 2369.035 2906.595 2369.205 ;
        RECT 2912.865 2369.035 2913.035 2369.205 ;
        RECT 2913.325 2369.035 2913.495 2369.205 ;
        RECT 2913.785 2369.035 2913.955 2369.205 ;
        RECT 5.665 2363.595 5.835 2363.765 ;
        RECT 6.125 2363.595 6.295 2363.765 ;
        RECT 6.585 2363.595 6.755 2363.765 ;
        RECT 2906.425 2363.595 2906.595 2363.765 ;
        RECT 2912.865 2363.595 2913.035 2363.765 ;
        RECT 2913.325 2363.595 2913.495 2363.765 ;
        RECT 2913.785 2363.595 2913.955 2363.765 ;
        RECT 5.665 2358.155 5.835 2358.325 ;
        RECT 6.125 2358.155 6.295 2358.325 ;
        RECT 6.585 2358.155 6.755 2358.325 ;
        RECT 2906.425 2358.155 2906.595 2358.325 ;
        RECT 2912.865 2358.155 2913.035 2358.325 ;
        RECT 2913.325 2358.155 2913.495 2358.325 ;
        RECT 2913.785 2358.155 2913.955 2358.325 ;
        RECT 5.665 2352.715 5.835 2352.885 ;
        RECT 6.125 2352.715 6.295 2352.885 ;
        RECT 6.585 2352.715 6.755 2352.885 ;
        RECT 2906.425 2352.715 2906.595 2352.885 ;
        RECT 2912.865 2352.715 2913.035 2352.885 ;
        RECT 2913.325 2352.715 2913.495 2352.885 ;
        RECT 2913.785 2352.715 2913.955 2352.885 ;
        RECT 5.665 2347.275 5.835 2347.445 ;
        RECT 6.125 2347.275 6.295 2347.445 ;
        RECT 6.585 2347.275 6.755 2347.445 ;
        RECT 2906.425 2347.275 2906.595 2347.445 ;
        RECT 2912.865 2347.275 2913.035 2347.445 ;
        RECT 2913.325 2347.275 2913.495 2347.445 ;
        RECT 2913.785 2347.275 2913.955 2347.445 ;
        RECT 5.665 2341.835 5.835 2342.005 ;
        RECT 6.125 2341.835 6.295 2342.005 ;
        RECT 6.585 2341.835 6.755 2342.005 ;
        RECT 2906.425 2341.835 2906.595 2342.005 ;
        RECT 2912.865 2341.835 2913.035 2342.005 ;
        RECT 2913.325 2341.835 2913.495 2342.005 ;
        RECT 2913.785 2341.835 2913.955 2342.005 ;
        RECT 5.665 2336.395 5.835 2336.565 ;
        RECT 6.125 2336.395 6.295 2336.565 ;
        RECT 6.585 2336.395 6.755 2336.565 ;
        RECT 2906.425 2336.395 2906.595 2336.565 ;
        RECT 2912.865 2336.395 2913.035 2336.565 ;
        RECT 2913.325 2336.395 2913.495 2336.565 ;
        RECT 2913.785 2336.395 2913.955 2336.565 ;
        RECT 5.665 2330.955 5.835 2331.125 ;
        RECT 6.125 2330.955 6.295 2331.125 ;
        RECT 6.585 2330.955 6.755 2331.125 ;
        RECT 2906.425 2330.955 2906.595 2331.125 ;
        RECT 2912.865 2330.955 2913.035 2331.125 ;
        RECT 2913.325 2330.955 2913.495 2331.125 ;
        RECT 2913.785 2330.955 2913.955 2331.125 ;
        RECT 5.665 2325.515 5.835 2325.685 ;
        RECT 6.125 2325.515 6.295 2325.685 ;
        RECT 6.585 2325.515 6.755 2325.685 ;
        RECT 2906.425 2325.515 2906.595 2325.685 ;
        RECT 2912.865 2325.515 2913.035 2325.685 ;
        RECT 2913.325 2325.515 2913.495 2325.685 ;
        RECT 2913.785 2325.515 2913.955 2325.685 ;
        RECT 5.665 2320.075 5.835 2320.245 ;
        RECT 6.125 2320.075 6.295 2320.245 ;
        RECT 6.585 2320.075 6.755 2320.245 ;
        RECT 2906.425 2320.075 2906.595 2320.245 ;
        RECT 2912.865 2320.075 2913.035 2320.245 ;
        RECT 2913.325 2320.075 2913.495 2320.245 ;
        RECT 2913.785 2320.075 2913.955 2320.245 ;
        RECT 5.665 2314.635 5.835 2314.805 ;
        RECT 6.125 2314.635 6.295 2314.805 ;
        RECT 6.585 2314.635 6.755 2314.805 ;
        RECT 2906.425 2314.635 2906.595 2314.805 ;
        RECT 2912.865 2314.635 2913.035 2314.805 ;
        RECT 2913.325 2314.635 2913.495 2314.805 ;
        RECT 2913.785 2314.635 2913.955 2314.805 ;
        RECT 5.665 2309.195 5.835 2309.365 ;
        RECT 6.125 2309.195 6.295 2309.365 ;
        RECT 6.585 2309.195 6.755 2309.365 ;
        RECT 2906.425 2309.195 2906.595 2309.365 ;
        RECT 2912.865 2309.195 2913.035 2309.365 ;
        RECT 2913.325 2309.195 2913.495 2309.365 ;
        RECT 2913.785 2309.195 2913.955 2309.365 ;
        RECT 5.665 2303.755 5.835 2303.925 ;
        RECT 6.125 2303.755 6.295 2303.925 ;
        RECT 6.585 2303.755 6.755 2303.925 ;
        RECT 2906.425 2303.755 2906.595 2303.925 ;
        RECT 2912.865 2303.755 2913.035 2303.925 ;
        RECT 2913.325 2303.755 2913.495 2303.925 ;
        RECT 2913.785 2303.755 2913.955 2303.925 ;
        RECT 5.665 2298.315 5.835 2298.485 ;
        RECT 6.125 2298.315 6.295 2298.485 ;
        RECT 6.585 2298.315 6.755 2298.485 ;
        RECT 2906.425 2298.315 2906.595 2298.485 ;
        RECT 2912.865 2298.315 2913.035 2298.485 ;
        RECT 2913.325 2298.315 2913.495 2298.485 ;
        RECT 2913.785 2298.315 2913.955 2298.485 ;
        RECT 5.665 2292.875 5.835 2293.045 ;
        RECT 6.125 2292.875 6.295 2293.045 ;
        RECT 6.585 2292.875 6.755 2293.045 ;
        RECT 2906.425 2292.875 2906.595 2293.045 ;
        RECT 2912.865 2292.875 2913.035 2293.045 ;
        RECT 2913.325 2292.875 2913.495 2293.045 ;
        RECT 2913.785 2292.875 2913.955 2293.045 ;
        RECT 5.665 2287.435 5.835 2287.605 ;
        RECT 6.125 2287.435 6.295 2287.605 ;
        RECT 6.585 2287.435 6.755 2287.605 ;
        RECT 2906.425 2287.435 2906.595 2287.605 ;
        RECT 2912.865 2287.435 2913.035 2287.605 ;
        RECT 2913.325 2287.435 2913.495 2287.605 ;
        RECT 2913.785 2287.435 2913.955 2287.605 ;
        RECT 5.665 2281.995 5.835 2282.165 ;
        RECT 6.125 2281.995 6.295 2282.165 ;
        RECT 6.585 2281.995 6.755 2282.165 ;
        RECT 2906.425 2281.995 2906.595 2282.165 ;
        RECT 2912.865 2281.995 2913.035 2282.165 ;
        RECT 2913.325 2281.995 2913.495 2282.165 ;
        RECT 2913.785 2281.995 2913.955 2282.165 ;
        RECT 5.665 2276.555 5.835 2276.725 ;
        RECT 6.125 2276.555 6.295 2276.725 ;
        RECT 6.585 2276.555 6.755 2276.725 ;
        RECT 2906.425 2276.555 2906.595 2276.725 ;
        RECT 2912.865 2276.555 2913.035 2276.725 ;
        RECT 2913.325 2276.555 2913.495 2276.725 ;
        RECT 2913.785 2276.555 2913.955 2276.725 ;
        RECT 5.665 2271.115 5.835 2271.285 ;
        RECT 6.125 2271.115 6.295 2271.285 ;
        RECT 6.585 2271.115 6.755 2271.285 ;
        RECT 2906.425 2271.115 2906.595 2271.285 ;
        RECT 2912.865 2271.115 2913.035 2271.285 ;
        RECT 2913.325 2271.115 2913.495 2271.285 ;
        RECT 2913.785 2271.115 2913.955 2271.285 ;
        RECT 5.665 2265.675 5.835 2265.845 ;
        RECT 6.125 2265.675 6.295 2265.845 ;
        RECT 6.585 2265.675 6.755 2265.845 ;
        RECT 2906.425 2265.675 2906.595 2265.845 ;
        RECT 2909.185 2265.675 2909.355 2265.845 ;
        RECT 2909.645 2265.675 2909.815 2265.845 ;
        RECT 2910.105 2265.675 2910.275 2265.845 ;
        RECT 2912.865 2265.675 2913.035 2265.845 ;
        RECT 2913.325 2265.675 2913.495 2265.845 ;
        RECT 2913.785 2265.675 2913.955 2265.845 ;
        RECT 5.665 2260.235 5.835 2260.405 ;
        RECT 6.125 2260.235 6.295 2260.405 ;
        RECT 6.585 2260.235 6.755 2260.405 ;
        RECT 2906.425 2260.235 2906.595 2260.405 ;
        RECT 2912.865 2260.235 2913.035 2260.405 ;
        RECT 2913.325 2260.235 2913.495 2260.405 ;
        RECT 2913.785 2260.235 2913.955 2260.405 ;
        RECT 5.665 2254.795 5.835 2254.965 ;
        RECT 6.125 2254.795 6.295 2254.965 ;
        RECT 6.585 2254.795 6.755 2254.965 ;
        RECT 2906.425 2254.795 2906.595 2254.965 ;
        RECT 2912.865 2254.795 2913.035 2254.965 ;
        RECT 2913.325 2254.795 2913.495 2254.965 ;
        RECT 2913.785 2254.795 2913.955 2254.965 ;
        RECT 5.665 2249.355 5.835 2249.525 ;
        RECT 6.125 2249.355 6.295 2249.525 ;
        RECT 6.585 2249.355 6.755 2249.525 ;
        RECT 2906.425 2249.355 2906.595 2249.525 ;
        RECT 2912.865 2249.355 2913.035 2249.525 ;
        RECT 2913.325 2249.355 2913.495 2249.525 ;
        RECT 2913.785 2249.355 2913.955 2249.525 ;
        RECT 5.665 2243.915 5.835 2244.085 ;
        RECT 6.125 2243.915 6.295 2244.085 ;
        RECT 6.585 2243.915 6.755 2244.085 ;
        RECT 2906.425 2243.915 2906.595 2244.085 ;
        RECT 2912.865 2243.915 2913.035 2244.085 ;
        RECT 2913.325 2243.915 2913.495 2244.085 ;
        RECT 2913.785 2243.915 2913.955 2244.085 ;
        RECT 5.665 2238.475 5.835 2238.645 ;
        RECT 6.125 2238.475 6.295 2238.645 ;
        RECT 6.585 2238.475 6.755 2238.645 ;
        RECT 2906.425 2238.475 2906.595 2238.645 ;
        RECT 2912.865 2238.475 2913.035 2238.645 ;
        RECT 2913.325 2238.475 2913.495 2238.645 ;
        RECT 2913.785 2238.475 2913.955 2238.645 ;
        RECT 5.665 2233.035 5.835 2233.205 ;
        RECT 6.125 2233.035 6.295 2233.205 ;
        RECT 6.585 2233.035 6.755 2233.205 ;
        RECT 2906.425 2233.035 2906.595 2233.205 ;
        RECT 2912.865 2233.035 2913.035 2233.205 ;
        RECT 2913.325 2233.035 2913.495 2233.205 ;
        RECT 2913.785 2233.035 2913.955 2233.205 ;
        RECT 5.665 2227.595 5.835 2227.765 ;
        RECT 6.125 2227.595 6.295 2227.765 ;
        RECT 6.585 2227.595 6.755 2227.765 ;
        RECT 2906.425 2227.595 2906.595 2227.765 ;
        RECT 2912.865 2227.595 2913.035 2227.765 ;
        RECT 2913.325 2227.595 2913.495 2227.765 ;
        RECT 2913.785 2227.595 2913.955 2227.765 ;
        RECT 5.665 2222.155 5.835 2222.325 ;
        RECT 6.125 2222.155 6.295 2222.325 ;
        RECT 6.585 2222.155 6.755 2222.325 ;
        RECT 2906.425 2222.155 2906.595 2222.325 ;
        RECT 2912.865 2222.155 2913.035 2222.325 ;
        RECT 2913.325 2222.155 2913.495 2222.325 ;
        RECT 2913.785 2222.155 2913.955 2222.325 ;
        RECT 5.665 2216.715 5.835 2216.885 ;
        RECT 6.125 2216.715 6.295 2216.885 ;
        RECT 6.585 2216.715 6.755 2216.885 ;
        RECT 2906.425 2216.715 2906.595 2216.885 ;
        RECT 2912.865 2216.715 2913.035 2216.885 ;
        RECT 2913.325 2216.715 2913.495 2216.885 ;
        RECT 2913.785 2216.715 2913.955 2216.885 ;
        RECT 5.665 2211.275 5.835 2211.445 ;
        RECT 6.125 2211.275 6.295 2211.445 ;
        RECT 6.585 2211.275 6.755 2211.445 ;
        RECT 2906.425 2211.275 2906.595 2211.445 ;
        RECT 2912.865 2211.275 2913.035 2211.445 ;
        RECT 2913.325 2211.275 2913.495 2211.445 ;
        RECT 2913.785 2211.275 2913.955 2211.445 ;
        RECT 5.665 2205.835 5.835 2206.005 ;
        RECT 6.125 2205.835 6.295 2206.005 ;
        RECT 6.585 2205.835 6.755 2206.005 ;
        RECT 2906.425 2205.835 2906.595 2206.005 ;
        RECT 2912.865 2205.835 2913.035 2206.005 ;
        RECT 2913.325 2205.835 2913.495 2206.005 ;
        RECT 2913.785 2205.835 2913.955 2206.005 ;
        RECT 5.665 2200.395 5.835 2200.565 ;
        RECT 6.125 2200.395 6.295 2200.565 ;
        RECT 6.585 2200.395 6.755 2200.565 ;
        RECT 2906.425 2200.395 2906.595 2200.565 ;
        RECT 2912.865 2200.395 2913.035 2200.565 ;
        RECT 2913.325 2200.395 2913.495 2200.565 ;
        RECT 2913.785 2200.395 2913.955 2200.565 ;
        RECT 5.665 2194.955 5.835 2195.125 ;
        RECT 6.125 2194.955 6.295 2195.125 ;
        RECT 6.585 2194.955 6.755 2195.125 ;
        RECT 2906.425 2194.955 2906.595 2195.125 ;
        RECT 2912.865 2194.955 2913.035 2195.125 ;
        RECT 2913.325 2194.955 2913.495 2195.125 ;
        RECT 2913.785 2194.955 2913.955 2195.125 ;
        RECT 5.665 2189.515 5.835 2189.685 ;
        RECT 6.125 2189.515 6.295 2189.685 ;
        RECT 6.585 2189.515 6.755 2189.685 ;
        RECT 2906.425 2189.515 2906.595 2189.685 ;
        RECT 2912.865 2189.515 2913.035 2189.685 ;
        RECT 2913.325 2189.515 2913.495 2189.685 ;
        RECT 2913.785 2189.515 2913.955 2189.685 ;
        RECT 5.665 2184.075 5.835 2184.245 ;
        RECT 6.125 2184.075 6.295 2184.245 ;
        RECT 6.585 2184.075 6.755 2184.245 ;
        RECT 2906.425 2184.075 2906.595 2184.245 ;
        RECT 2912.865 2184.075 2913.035 2184.245 ;
        RECT 2913.325 2184.075 2913.495 2184.245 ;
        RECT 2913.785 2184.075 2913.955 2184.245 ;
        RECT 5.665 2178.635 5.835 2178.805 ;
        RECT 6.125 2178.635 6.295 2178.805 ;
        RECT 6.585 2178.635 6.755 2178.805 ;
        RECT 2906.425 2178.635 2906.595 2178.805 ;
        RECT 2912.865 2178.635 2913.035 2178.805 ;
        RECT 2913.325 2178.635 2913.495 2178.805 ;
        RECT 2913.785 2178.635 2913.955 2178.805 ;
        RECT 5.665 2173.195 5.835 2173.365 ;
        RECT 6.125 2173.195 6.295 2173.365 ;
        RECT 6.585 2173.195 6.755 2173.365 ;
        RECT 2906.425 2173.195 2906.595 2173.365 ;
        RECT 2912.865 2173.195 2913.035 2173.365 ;
        RECT 2913.325 2173.195 2913.495 2173.365 ;
        RECT 2913.785 2173.195 2913.955 2173.365 ;
        RECT 5.665 2167.755 5.835 2167.925 ;
        RECT 6.125 2167.755 6.295 2167.925 ;
        RECT 6.585 2167.755 6.755 2167.925 ;
        RECT 2906.425 2167.755 2906.595 2167.925 ;
        RECT 2912.865 2167.755 2913.035 2167.925 ;
        RECT 2913.325 2167.755 2913.495 2167.925 ;
        RECT 2913.785 2167.755 2913.955 2167.925 ;
        RECT 5.665 2162.315 5.835 2162.485 ;
        RECT 6.125 2162.315 6.295 2162.485 ;
        RECT 6.585 2162.315 6.755 2162.485 ;
        RECT 2906.425 2162.315 2906.595 2162.485 ;
        RECT 2912.865 2162.315 2913.035 2162.485 ;
        RECT 2913.325 2162.315 2913.495 2162.485 ;
        RECT 2913.785 2162.315 2913.955 2162.485 ;
        RECT 5.665 2156.875 5.835 2157.045 ;
        RECT 6.125 2156.875 6.295 2157.045 ;
        RECT 6.585 2156.875 6.755 2157.045 ;
        RECT 2906.425 2156.875 2906.595 2157.045 ;
        RECT 2912.865 2156.875 2913.035 2157.045 ;
        RECT 2913.325 2156.875 2913.495 2157.045 ;
        RECT 2913.785 2156.875 2913.955 2157.045 ;
        RECT 5.665 2151.435 5.835 2151.605 ;
        RECT 6.125 2151.435 6.295 2151.605 ;
        RECT 6.585 2151.435 6.755 2151.605 ;
        RECT 2906.425 2151.435 2906.595 2151.605 ;
        RECT 2912.865 2151.435 2913.035 2151.605 ;
        RECT 2913.325 2151.435 2913.495 2151.605 ;
        RECT 2913.785 2151.435 2913.955 2151.605 ;
        RECT 5.665 2145.995 5.835 2146.165 ;
        RECT 6.125 2145.995 6.295 2146.165 ;
        RECT 6.585 2145.995 6.755 2146.165 ;
        RECT 2906.425 2145.995 2906.595 2146.165 ;
        RECT 2912.865 2145.995 2913.035 2146.165 ;
        RECT 2913.325 2145.995 2913.495 2146.165 ;
        RECT 2913.785 2145.995 2913.955 2146.165 ;
        RECT 5.665 2140.555 5.835 2140.725 ;
        RECT 6.125 2140.555 6.295 2140.725 ;
        RECT 6.585 2140.555 6.755 2140.725 ;
        RECT 2906.425 2140.555 2906.595 2140.725 ;
        RECT 2912.865 2140.555 2913.035 2140.725 ;
        RECT 2913.325 2140.555 2913.495 2140.725 ;
        RECT 2913.785 2140.555 2913.955 2140.725 ;
        RECT 5.665 2135.115 5.835 2135.285 ;
        RECT 6.125 2135.115 6.295 2135.285 ;
        RECT 6.585 2135.115 6.755 2135.285 ;
        RECT 2906.425 2135.115 2906.595 2135.285 ;
        RECT 2912.865 2135.115 2913.035 2135.285 ;
        RECT 2913.325 2135.115 2913.495 2135.285 ;
        RECT 2913.785 2135.115 2913.955 2135.285 ;
        RECT 5.665 2129.675 5.835 2129.845 ;
        RECT 6.125 2129.675 6.295 2129.845 ;
        RECT 6.585 2129.675 6.755 2129.845 ;
        RECT 2906.425 2129.675 2906.595 2129.845 ;
        RECT 2912.865 2129.675 2913.035 2129.845 ;
        RECT 2913.325 2129.675 2913.495 2129.845 ;
        RECT 2913.785 2129.675 2913.955 2129.845 ;
        RECT 5.665 2124.235 5.835 2124.405 ;
        RECT 6.125 2124.235 6.295 2124.405 ;
        RECT 6.585 2124.235 6.755 2124.405 ;
        RECT 2906.425 2124.235 2906.595 2124.405 ;
        RECT 2912.865 2124.235 2913.035 2124.405 ;
        RECT 2913.325 2124.235 2913.495 2124.405 ;
        RECT 2913.785 2124.235 2913.955 2124.405 ;
        RECT 5.665 2118.795 5.835 2118.965 ;
        RECT 6.125 2118.795 6.295 2118.965 ;
        RECT 6.585 2118.795 6.755 2118.965 ;
        RECT 2906.425 2118.795 2906.595 2118.965 ;
        RECT 2909.185 2118.795 2909.355 2118.965 ;
        RECT 2909.645 2118.795 2909.815 2118.965 ;
        RECT 2910.105 2118.795 2910.275 2118.965 ;
        RECT 2912.865 2118.795 2913.035 2118.965 ;
        RECT 2913.325 2118.795 2913.495 2118.965 ;
        RECT 2913.785 2118.795 2913.955 2118.965 ;
        RECT 5.665 2113.355 5.835 2113.525 ;
        RECT 6.125 2113.355 6.295 2113.525 ;
        RECT 6.585 2113.355 6.755 2113.525 ;
        RECT 2906.425 2113.355 2906.595 2113.525 ;
        RECT 2912.865 2113.355 2913.035 2113.525 ;
        RECT 2913.325 2113.355 2913.495 2113.525 ;
        RECT 2913.785 2113.355 2913.955 2113.525 ;
        RECT 5.665 2107.915 5.835 2108.085 ;
        RECT 6.125 2107.915 6.295 2108.085 ;
        RECT 6.585 2107.915 6.755 2108.085 ;
        RECT 2906.425 2107.915 2906.595 2108.085 ;
        RECT 2912.865 2107.915 2913.035 2108.085 ;
        RECT 2913.325 2107.915 2913.495 2108.085 ;
        RECT 2913.785 2107.915 2913.955 2108.085 ;
        RECT 5.665 2102.475 5.835 2102.645 ;
        RECT 6.125 2102.475 6.295 2102.645 ;
        RECT 6.585 2102.475 6.755 2102.645 ;
        RECT 2906.425 2102.475 2906.595 2102.645 ;
        RECT 2912.865 2102.475 2913.035 2102.645 ;
        RECT 2913.325 2102.475 2913.495 2102.645 ;
        RECT 2913.785 2102.475 2913.955 2102.645 ;
        RECT 5.665 2097.035 5.835 2097.205 ;
        RECT 6.125 2097.035 6.295 2097.205 ;
        RECT 6.585 2097.035 6.755 2097.205 ;
        RECT 2906.425 2097.035 2906.595 2097.205 ;
        RECT 2912.865 2097.035 2913.035 2097.205 ;
        RECT 2913.325 2097.035 2913.495 2097.205 ;
        RECT 2913.785 2097.035 2913.955 2097.205 ;
        RECT 5.665 2091.595 5.835 2091.765 ;
        RECT 6.125 2091.595 6.295 2091.765 ;
        RECT 6.585 2091.595 6.755 2091.765 ;
        RECT 2906.425 2091.595 2906.595 2091.765 ;
        RECT 2912.865 2091.595 2913.035 2091.765 ;
        RECT 2913.325 2091.595 2913.495 2091.765 ;
        RECT 2913.785 2091.595 2913.955 2091.765 ;
        RECT 5.665 2086.155 5.835 2086.325 ;
        RECT 6.125 2086.155 6.295 2086.325 ;
        RECT 6.585 2086.155 6.755 2086.325 ;
        RECT 2906.425 2086.155 2906.595 2086.325 ;
        RECT 2912.865 2086.155 2913.035 2086.325 ;
        RECT 2913.325 2086.155 2913.495 2086.325 ;
        RECT 2913.785 2086.155 2913.955 2086.325 ;
        RECT 5.665 2080.715 5.835 2080.885 ;
        RECT 6.125 2080.715 6.295 2080.885 ;
        RECT 6.585 2080.715 6.755 2080.885 ;
        RECT 2906.425 2080.715 2906.595 2080.885 ;
        RECT 2912.865 2080.715 2913.035 2080.885 ;
        RECT 2913.325 2080.715 2913.495 2080.885 ;
        RECT 2913.785 2080.715 2913.955 2080.885 ;
        RECT 5.665 2075.275 5.835 2075.445 ;
        RECT 6.125 2075.275 6.295 2075.445 ;
        RECT 6.585 2075.275 6.755 2075.445 ;
        RECT 2906.425 2075.275 2906.595 2075.445 ;
        RECT 2912.865 2075.275 2913.035 2075.445 ;
        RECT 2913.325 2075.275 2913.495 2075.445 ;
        RECT 2913.785 2075.275 2913.955 2075.445 ;
        RECT 5.665 2069.835 5.835 2070.005 ;
        RECT 6.125 2069.835 6.295 2070.005 ;
        RECT 6.585 2069.835 6.755 2070.005 ;
        RECT 2906.425 2069.835 2906.595 2070.005 ;
        RECT 2912.865 2069.835 2913.035 2070.005 ;
        RECT 2913.325 2069.835 2913.495 2070.005 ;
        RECT 2913.785 2069.835 2913.955 2070.005 ;
        RECT 5.665 2064.395 5.835 2064.565 ;
        RECT 6.125 2064.395 6.295 2064.565 ;
        RECT 6.585 2064.395 6.755 2064.565 ;
        RECT 2906.425 2064.395 2906.595 2064.565 ;
        RECT 2912.865 2064.395 2913.035 2064.565 ;
        RECT 2913.325 2064.395 2913.495 2064.565 ;
        RECT 2913.785 2064.395 2913.955 2064.565 ;
        RECT 5.665 2058.955 5.835 2059.125 ;
        RECT 6.125 2058.955 6.295 2059.125 ;
        RECT 6.585 2058.955 6.755 2059.125 ;
        RECT 2906.425 2058.955 2906.595 2059.125 ;
        RECT 2912.865 2058.955 2913.035 2059.125 ;
        RECT 2913.325 2058.955 2913.495 2059.125 ;
        RECT 2913.785 2058.955 2913.955 2059.125 ;
        RECT 5.665 2053.515 5.835 2053.685 ;
        RECT 6.125 2053.515 6.295 2053.685 ;
        RECT 6.585 2053.515 6.755 2053.685 ;
        RECT 2906.425 2053.515 2906.595 2053.685 ;
        RECT 2912.865 2053.515 2913.035 2053.685 ;
        RECT 2913.325 2053.515 2913.495 2053.685 ;
        RECT 2913.785 2053.515 2913.955 2053.685 ;
        RECT 5.665 2048.075 5.835 2048.245 ;
        RECT 6.125 2048.075 6.295 2048.245 ;
        RECT 6.585 2048.075 6.755 2048.245 ;
        RECT 2906.425 2048.075 2906.595 2048.245 ;
        RECT 2912.865 2048.075 2913.035 2048.245 ;
        RECT 2913.325 2048.075 2913.495 2048.245 ;
        RECT 2913.785 2048.075 2913.955 2048.245 ;
        RECT 5.665 2042.635 5.835 2042.805 ;
        RECT 6.125 2042.635 6.295 2042.805 ;
        RECT 6.585 2042.635 6.755 2042.805 ;
        RECT 2906.425 2042.635 2906.595 2042.805 ;
        RECT 2912.865 2042.635 2913.035 2042.805 ;
        RECT 2913.325 2042.635 2913.495 2042.805 ;
        RECT 2913.785 2042.635 2913.955 2042.805 ;
        RECT 5.665 2037.195 5.835 2037.365 ;
        RECT 6.125 2037.195 6.295 2037.365 ;
        RECT 6.585 2037.195 6.755 2037.365 ;
        RECT 2906.425 2037.195 2906.595 2037.365 ;
        RECT 2912.865 2037.195 2913.035 2037.365 ;
        RECT 2913.325 2037.195 2913.495 2037.365 ;
        RECT 2913.785 2037.195 2913.955 2037.365 ;
        RECT 5.665 2031.755 5.835 2031.925 ;
        RECT 6.125 2031.755 6.295 2031.925 ;
        RECT 6.585 2031.755 6.755 2031.925 ;
        RECT 2906.425 2031.755 2906.595 2031.925 ;
        RECT 2912.865 2031.755 2913.035 2031.925 ;
        RECT 2913.325 2031.755 2913.495 2031.925 ;
        RECT 2913.785 2031.755 2913.955 2031.925 ;
        RECT 5.665 2026.315 5.835 2026.485 ;
        RECT 6.125 2026.315 6.295 2026.485 ;
        RECT 6.585 2026.315 6.755 2026.485 ;
        RECT 2906.425 2026.315 2906.595 2026.485 ;
        RECT 2912.865 2026.315 2913.035 2026.485 ;
        RECT 2913.325 2026.315 2913.495 2026.485 ;
        RECT 2913.785 2026.315 2913.955 2026.485 ;
        RECT 5.665 2020.875 5.835 2021.045 ;
        RECT 6.125 2020.875 6.295 2021.045 ;
        RECT 6.585 2020.875 6.755 2021.045 ;
        RECT 2906.425 2020.875 2906.595 2021.045 ;
        RECT 2912.865 2020.875 2913.035 2021.045 ;
        RECT 2913.325 2020.875 2913.495 2021.045 ;
        RECT 2913.785 2020.875 2913.955 2021.045 ;
        RECT 5.665 2015.435 5.835 2015.605 ;
        RECT 6.125 2015.435 6.295 2015.605 ;
        RECT 6.585 2015.435 6.755 2015.605 ;
        RECT 2906.425 2015.435 2906.595 2015.605 ;
        RECT 2912.865 2015.435 2913.035 2015.605 ;
        RECT 2913.325 2015.435 2913.495 2015.605 ;
        RECT 2913.785 2015.435 2913.955 2015.605 ;
        RECT 5.665 2009.995 5.835 2010.165 ;
        RECT 6.125 2009.995 6.295 2010.165 ;
        RECT 6.585 2009.995 6.755 2010.165 ;
        RECT 2906.425 2009.995 2906.595 2010.165 ;
        RECT 2912.865 2009.995 2913.035 2010.165 ;
        RECT 2913.325 2009.995 2913.495 2010.165 ;
        RECT 2913.785 2009.995 2913.955 2010.165 ;
        RECT 5.665 2004.555 5.835 2004.725 ;
        RECT 6.125 2004.555 6.295 2004.725 ;
        RECT 6.585 2004.555 6.755 2004.725 ;
        RECT 2906.425 2004.555 2906.595 2004.725 ;
        RECT 2912.865 2004.555 2913.035 2004.725 ;
        RECT 2913.325 2004.555 2913.495 2004.725 ;
        RECT 2913.785 2004.555 2913.955 2004.725 ;
        RECT 5.665 1999.115 5.835 1999.285 ;
        RECT 6.125 1999.115 6.295 1999.285 ;
        RECT 6.585 1999.115 6.755 1999.285 ;
        RECT 2906.425 1999.115 2906.595 1999.285 ;
        RECT 2912.865 1999.115 2913.035 1999.285 ;
        RECT 2913.325 1999.115 2913.495 1999.285 ;
        RECT 2913.785 1999.115 2913.955 1999.285 ;
        RECT 5.665 1993.675 5.835 1993.845 ;
        RECT 6.125 1993.675 6.295 1993.845 ;
        RECT 6.585 1993.675 6.755 1993.845 ;
        RECT 2906.425 1993.675 2906.595 1993.845 ;
        RECT 2912.865 1993.675 2913.035 1993.845 ;
        RECT 2913.325 1993.675 2913.495 1993.845 ;
        RECT 2913.785 1993.675 2913.955 1993.845 ;
        RECT 5.665 1988.235 5.835 1988.405 ;
        RECT 6.125 1988.235 6.295 1988.405 ;
        RECT 6.585 1988.235 6.755 1988.405 ;
        RECT 2906.425 1988.235 2906.595 1988.405 ;
        RECT 2912.865 1988.235 2913.035 1988.405 ;
        RECT 2913.325 1988.235 2913.495 1988.405 ;
        RECT 2913.785 1988.235 2913.955 1988.405 ;
        RECT 5.665 1982.795 5.835 1982.965 ;
        RECT 6.125 1982.795 6.295 1982.965 ;
        RECT 6.585 1982.795 6.755 1982.965 ;
        RECT 8.885 1982.795 9.055 1982.965 ;
        RECT 9.345 1982.795 9.515 1982.965 ;
        RECT 9.805 1982.795 9.975 1982.965 ;
        RECT 2906.425 1982.795 2906.595 1982.965 ;
        RECT 2912.865 1982.795 2913.035 1982.965 ;
        RECT 2913.325 1982.795 2913.495 1982.965 ;
        RECT 2913.785 1982.795 2913.955 1982.965 ;
        RECT 5.665 1977.355 5.835 1977.525 ;
        RECT 6.125 1977.355 6.295 1977.525 ;
        RECT 6.585 1977.355 6.755 1977.525 ;
        RECT 2906.425 1977.355 2906.595 1977.525 ;
        RECT 2912.865 1977.355 2913.035 1977.525 ;
        RECT 2913.325 1977.355 2913.495 1977.525 ;
        RECT 2913.785 1977.355 2913.955 1977.525 ;
        RECT 5.665 1971.915 5.835 1972.085 ;
        RECT 6.125 1971.915 6.295 1972.085 ;
        RECT 6.585 1971.915 6.755 1972.085 ;
        RECT 2906.425 1971.915 2906.595 1972.085 ;
        RECT 2912.865 1971.915 2913.035 1972.085 ;
        RECT 2913.325 1971.915 2913.495 1972.085 ;
        RECT 2913.785 1971.915 2913.955 1972.085 ;
        RECT 5.665 1966.475 5.835 1966.645 ;
        RECT 6.125 1966.475 6.295 1966.645 ;
        RECT 6.585 1966.475 6.755 1966.645 ;
        RECT 2906.425 1966.475 2906.595 1966.645 ;
        RECT 2912.865 1966.475 2913.035 1966.645 ;
        RECT 2913.325 1966.475 2913.495 1966.645 ;
        RECT 2913.785 1966.475 2913.955 1966.645 ;
        RECT 5.665 1961.035 5.835 1961.205 ;
        RECT 6.125 1961.035 6.295 1961.205 ;
        RECT 6.585 1961.035 6.755 1961.205 ;
        RECT 2906.425 1961.035 2906.595 1961.205 ;
        RECT 2912.865 1961.035 2913.035 1961.205 ;
        RECT 2913.325 1961.035 2913.495 1961.205 ;
        RECT 2913.785 1961.035 2913.955 1961.205 ;
        RECT 5.665 1955.595 5.835 1955.765 ;
        RECT 6.125 1955.595 6.295 1955.765 ;
        RECT 6.585 1955.595 6.755 1955.765 ;
        RECT 8.885 1955.595 9.055 1955.765 ;
        RECT 9.345 1955.595 9.515 1955.765 ;
        RECT 9.805 1955.595 9.975 1955.765 ;
        RECT 2906.425 1955.595 2906.595 1955.765 ;
        RECT 2912.865 1955.595 2913.035 1955.765 ;
        RECT 2913.325 1955.595 2913.495 1955.765 ;
        RECT 2913.785 1955.595 2913.955 1955.765 ;
        RECT 5.665 1950.155 5.835 1950.325 ;
        RECT 6.125 1950.155 6.295 1950.325 ;
        RECT 6.585 1950.155 6.755 1950.325 ;
        RECT 2906.425 1950.155 2906.595 1950.325 ;
        RECT 2912.865 1950.155 2913.035 1950.325 ;
        RECT 2913.325 1950.155 2913.495 1950.325 ;
        RECT 2913.785 1950.155 2913.955 1950.325 ;
        RECT 5.665 1944.715 5.835 1944.885 ;
        RECT 6.125 1944.715 6.295 1944.885 ;
        RECT 6.585 1944.715 6.755 1944.885 ;
        RECT 2906.425 1944.715 2906.595 1944.885 ;
        RECT 2912.865 1944.715 2913.035 1944.885 ;
        RECT 2913.325 1944.715 2913.495 1944.885 ;
        RECT 2913.785 1944.715 2913.955 1944.885 ;
        RECT 5.665 1939.275 5.835 1939.445 ;
        RECT 6.125 1939.275 6.295 1939.445 ;
        RECT 6.585 1939.275 6.755 1939.445 ;
        RECT 2906.425 1939.275 2906.595 1939.445 ;
        RECT 2912.865 1939.275 2913.035 1939.445 ;
        RECT 2913.325 1939.275 2913.495 1939.445 ;
        RECT 2913.785 1939.275 2913.955 1939.445 ;
        RECT 5.665 1933.835 5.835 1934.005 ;
        RECT 6.125 1933.835 6.295 1934.005 ;
        RECT 6.585 1933.835 6.755 1934.005 ;
        RECT 2906.425 1933.835 2906.595 1934.005 ;
        RECT 2909.185 1933.835 2909.355 1934.005 ;
        RECT 2909.645 1933.835 2909.815 1934.005 ;
        RECT 2910.105 1933.835 2910.275 1934.005 ;
        RECT 2912.865 1933.835 2913.035 1934.005 ;
        RECT 2913.325 1933.835 2913.495 1934.005 ;
        RECT 2913.785 1933.835 2913.955 1934.005 ;
        RECT 5.665 1928.395 5.835 1928.565 ;
        RECT 6.125 1928.395 6.295 1928.565 ;
        RECT 6.585 1928.395 6.755 1928.565 ;
        RECT 2906.425 1928.395 2906.595 1928.565 ;
        RECT 2912.865 1928.395 2913.035 1928.565 ;
        RECT 2913.325 1928.395 2913.495 1928.565 ;
        RECT 2913.785 1928.395 2913.955 1928.565 ;
        RECT 5.665 1922.955 5.835 1923.125 ;
        RECT 6.125 1922.955 6.295 1923.125 ;
        RECT 6.585 1922.955 6.755 1923.125 ;
        RECT 2906.425 1922.955 2906.595 1923.125 ;
        RECT 2912.865 1922.955 2913.035 1923.125 ;
        RECT 2913.325 1922.955 2913.495 1923.125 ;
        RECT 2913.785 1922.955 2913.955 1923.125 ;
        RECT 5.665 1917.515 5.835 1917.685 ;
        RECT 6.125 1917.515 6.295 1917.685 ;
        RECT 6.585 1917.515 6.755 1917.685 ;
        RECT 2906.425 1917.515 2906.595 1917.685 ;
        RECT 2912.865 1917.515 2913.035 1917.685 ;
        RECT 2913.325 1917.515 2913.495 1917.685 ;
        RECT 2913.785 1917.515 2913.955 1917.685 ;
        RECT 5.665 1912.075 5.835 1912.245 ;
        RECT 6.125 1912.075 6.295 1912.245 ;
        RECT 6.585 1912.075 6.755 1912.245 ;
        RECT 2906.425 1912.075 2906.595 1912.245 ;
        RECT 2912.865 1912.075 2913.035 1912.245 ;
        RECT 2913.325 1912.075 2913.495 1912.245 ;
        RECT 2913.785 1912.075 2913.955 1912.245 ;
        RECT 5.665 1906.635 5.835 1906.805 ;
        RECT 6.125 1906.635 6.295 1906.805 ;
        RECT 6.585 1906.635 6.755 1906.805 ;
        RECT 2906.425 1906.635 2906.595 1906.805 ;
        RECT 2912.865 1906.635 2913.035 1906.805 ;
        RECT 2913.325 1906.635 2913.495 1906.805 ;
        RECT 2913.785 1906.635 2913.955 1906.805 ;
        RECT 5.665 1901.195 5.835 1901.365 ;
        RECT 6.125 1901.195 6.295 1901.365 ;
        RECT 6.585 1901.195 6.755 1901.365 ;
        RECT 2906.425 1901.195 2906.595 1901.365 ;
        RECT 2912.865 1901.195 2913.035 1901.365 ;
        RECT 2913.325 1901.195 2913.495 1901.365 ;
        RECT 2913.785 1901.195 2913.955 1901.365 ;
        RECT 5.665 1895.755 5.835 1895.925 ;
        RECT 6.125 1895.755 6.295 1895.925 ;
        RECT 6.585 1895.755 6.755 1895.925 ;
        RECT 2906.425 1895.755 2906.595 1895.925 ;
        RECT 2912.865 1895.755 2913.035 1895.925 ;
        RECT 2913.325 1895.755 2913.495 1895.925 ;
        RECT 2913.785 1895.755 2913.955 1895.925 ;
        RECT 5.665 1890.315 5.835 1890.485 ;
        RECT 6.125 1890.315 6.295 1890.485 ;
        RECT 6.585 1890.315 6.755 1890.485 ;
        RECT 2906.425 1890.315 2906.595 1890.485 ;
        RECT 2912.865 1890.315 2913.035 1890.485 ;
        RECT 2913.325 1890.315 2913.495 1890.485 ;
        RECT 2913.785 1890.315 2913.955 1890.485 ;
        RECT 5.665 1884.875 5.835 1885.045 ;
        RECT 6.125 1884.875 6.295 1885.045 ;
        RECT 6.585 1884.875 6.755 1885.045 ;
        RECT 2906.425 1884.875 2906.595 1885.045 ;
        RECT 2912.865 1884.875 2913.035 1885.045 ;
        RECT 2913.325 1884.875 2913.495 1885.045 ;
        RECT 2913.785 1884.875 2913.955 1885.045 ;
        RECT 5.665 1879.435 5.835 1879.605 ;
        RECT 6.125 1879.435 6.295 1879.605 ;
        RECT 6.585 1879.435 6.755 1879.605 ;
        RECT 2906.425 1879.435 2906.595 1879.605 ;
        RECT 2912.865 1879.435 2913.035 1879.605 ;
        RECT 2913.325 1879.435 2913.495 1879.605 ;
        RECT 2913.785 1879.435 2913.955 1879.605 ;
        RECT 5.665 1873.995 5.835 1874.165 ;
        RECT 6.125 1873.995 6.295 1874.165 ;
        RECT 6.585 1873.995 6.755 1874.165 ;
        RECT 2906.425 1873.995 2906.595 1874.165 ;
        RECT 2912.865 1873.995 2913.035 1874.165 ;
        RECT 2913.325 1873.995 2913.495 1874.165 ;
        RECT 2913.785 1873.995 2913.955 1874.165 ;
        RECT 5.665 1868.555 5.835 1868.725 ;
        RECT 6.125 1868.555 6.295 1868.725 ;
        RECT 6.585 1868.555 6.755 1868.725 ;
        RECT 2906.425 1868.555 2906.595 1868.725 ;
        RECT 2912.865 1868.555 2913.035 1868.725 ;
        RECT 2913.325 1868.555 2913.495 1868.725 ;
        RECT 2913.785 1868.555 2913.955 1868.725 ;
        RECT 5.665 1863.115 5.835 1863.285 ;
        RECT 6.125 1863.115 6.295 1863.285 ;
        RECT 6.585 1863.115 6.755 1863.285 ;
        RECT 2906.425 1863.115 2906.595 1863.285 ;
        RECT 2912.865 1863.115 2913.035 1863.285 ;
        RECT 2913.325 1863.115 2913.495 1863.285 ;
        RECT 2913.785 1863.115 2913.955 1863.285 ;
        RECT 5.665 1857.675 5.835 1857.845 ;
        RECT 6.125 1857.675 6.295 1857.845 ;
        RECT 6.585 1857.675 6.755 1857.845 ;
        RECT 2906.425 1857.675 2906.595 1857.845 ;
        RECT 2912.865 1857.675 2913.035 1857.845 ;
        RECT 2913.325 1857.675 2913.495 1857.845 ;
        RECT 2913.785 1857.675 2913.955 1857.845 ;
        RECT 5.665 1852.235 5.835 1852.405 ;
        RECT 6.125 1852.235 6.295 1852.405 ;
        RECT 6.585 1852.235 6.755 1852.405 ;
        RECT 2906.425 1852.235 2906.595 1852.405 ;
        RECT 2912.865 1852.235 2913.035 1852.405 ;
        RECT 2913.325 1852.235 2913.495 1852.405 ;
        RECT 2913.785 1852.235 2913.955 1852.405 ;
        RECT 5.665 1846.795 5.835 1846.965 ;
        RECT 6.125 1846.795 6.295 1846.965 ;
        RECT 6.585 1846.795 6.755 1846.965 ;
        RECT 2906.425 1846.795 2906.595 1846.965 ;
        RECT 2912.865 1846.795 2913.035 1846.965 ;
        RECT 2913.325 1846.795 2913.495 1846.965 ;
        RECT 2913.785 1846.795 2913.955 1846.965 ;
        RECT 5.665 1841.355 5.835 1841.525 ;
        RECT 6.125 1841.355 6.295 1841.525 ;
        RECT 6.585 1841.355 6.755 1841.525 ;
        RECT 2906.425 1841.355 2906.595 1841.525 ;
        RECT 2912.865 1841.355 2913.035 1841.525 ;
        RECT 2913.325 1841.355 2913.495 1841.525 ;
        RECT 2913.785 1841.355 2913.955 1841.525 ;
        RECT 5.665 1835.915 5.835 1836.085 ;
        RECT 6.125 1835.915 6.295 1836.085 ;
        RECT 6.585 1835.915 6.755 1836.085 ;
        RECT 2906.425 1835.915 2906.595 1836.085 ;
        RECT 2912.865 1835.915 2913.035 1836.085 ;
        RECT 2913.325 1835.915 2913.495 1836.085 ;
        RECT 2913.785 1835.915 2913.955 1836.085 ;
        RECT 5.665 1830.475 5.835 1830.645 ;
        RECT 6.125 1830.475 6.295 1830.645 ;
        RECT 6.585 1830.475 6.755 1830.645 ;
        RECT 2906.425 1830.475 2906.595 1830.645 ;
        RECT 2912.865 1830.475 2913.035 1830.645 ;
        RECT 2913.325 1830.475 2913.495 1830.645 ;
        RECT 2913.785 1830.475 2913.955 1830.645 ;
        RECT 5.665 1825.035 5.835 1825.205 ;
        RECT 6.125 1825.035 6.295 1825.205 ;
        RECT 6.585 1825.035 6.755 1825.205 ;
        RECT 2906.425 1825.035 2906.595 1825.205 ;
        RECT 2912.865 1825.035 2913.035 1825.205 ;
        RECT 2913.325 1825.035 2913.495 1825.205 ;
        RECT 2913.785 1825.035 2913.955 1825.205 ;
        RECT 5.665 1819.595 5.835 1819.765 ;
        RECT 6.125 1819.595 6.295 1819.765 ;
        RECT 6.585 1819.595 6.755 1819.765 ;
        RECT 2906.425 1819.595 2906.595 1819.765 ;
        RECT 2912.865 1819.595 2913.035 1819.765 ;
        RECT 2913.325 1819.595 2913.495 1819.765 ;
        RECT 2913.785 1819.595 2913.955 1819.765 ;
        RECT 5.665 1814.155 5.835 1814.325 ;
        RECT 6.125 1814.155 6.295 1814.325 ;
        RECT 6.585 1814.155 6.755 1814.325 ;
        RECT 2906.425 1814.155 2906.595 1814.325 ;
        RECT 2912.865 1814.155 2913.035 1814.325 ;
        RECT 2913.325 1814.155 2913.495 1814.325 ;
        RECT 2913.785 1814.155 2913.955 1814.325 ;
        RECT 5.665 1808.715 5.835 1808.885 ;
        RECT 6.125 1808.715 6.295 1808.885 ;
        RECT 6.585 1808.715 6.755 1808.885 ;
        RECT 2906.425 1808.715 2906.595 1808.885 ;
        RECT 2912.865 1808.715 2913.035 1808.885 ;
        RECT 2913.325 1808.715 2913.495 1808.885 ;
        RECT 2913.785 1808.715 2913.955 1808.885 ;
        RECT 5.665 1803.275 5.835 1803.445 ;
        RECT 6.125 1803.275 6.295 1803.445 ;
        RECT 6.585 1803.275 6.755 1803.445 ;
        RECT 2906.425 1803.275 2906.595 1803.445 ;
        RECT 2912.865 1803.275 2913.035 1803.445 ;
        RECT 2913.325 1803.275 2913.495 1803.445 ;
        RECT 2913.785 1803.275 2913.955 1803.445 ;
        RECT 5.665 1797.835 5.835 1798.005 ;
        RECT 6.125 1797.835 6.295 1798.005 ;
        RECT 6.585 1797.835 6.755 1798.005 ;
        RECT 2906.425 1797.835 2906.595 1798.005 ;
        RECT 2912.865 1797.835 2913.035 1798.005 ;
        RECT 2913.325 1797.835 2913.495 1798.005 ;
        RECT 2913.785 1797.835 2913.955 1798.005 ;
        RECT 5.665 1792.395 5.835 1792.565 ;
        RECT 6.125 1792.395 6.295 1792.565 ;
        RECT 6.585 1792.395 6.755 1792.565 ;
        RECT 2906.425 1792.395 2906.595 1792.565 ;
        RECT 2912.865 1792.395 2913.035 1792.565 ;
        RECT 2913.325 1792.395 2913.495 1792.565 ;
        RECT 2913.785 1792.395 2913.955 1792.565 ;
        RECT 5.665 1786.955 5.835 1787.125 ;
        RECT 6.125 1786.955 6.295 1787.125 ;
        RECT 6.585 1786.955 6.755 1787.125 ;
        RECT 2906.425 1786.955 2906.595 1787.125 ;
        RECT 2912.865 1786.955 2913.035 1787.125 ;
        RECT 2913.325 1786.955 2913.495 1787.125 ;
        RECT 2913.785 1786.955 2913.955 1787.125 ;
        RECT 5.665 1781.515 5.835 1781.685 ;
        RECT 6.125 1781.515 6.295 1781.685 ;
        RECT 6.585 1781.515 6.755 1781.685 ;
        RECT 2906.425 1781.515 2906.595 1781.685 ;
        RECT 2912.865 1781.515 2913.035 1781.685 ;
        RECT 2913.325 1781.515 2913.495 1781.685 ;
        RECT 2913.785 1781.515 2913.955 1781.685 ;
        RECT 5.665 1776.075 5.835 1776.245 ;
        RECT 6.125 1776.075 6.295 1776.245 ;
        RECT 6.585 1776.075 6.755 1776.245 ;
        RECT 8.885 1776.075 9.055 1776.245 ;
        RECT 9.345 1776.075 9.515 1776.245 ;
        RECT 9.805 1776.075 9.975 1776.245 ;
        RECT 2906.425 1776.075 2906.595 1776.245 ;
        RECT 2912.865 1776.075 2913.035 1776.245 ;
        RECT 2913.325 1776.075 2913.495 1776.245 ;
        RECT 2913.785 1776.075 2913.955 1776.245 ;
        RECT 5.665 1770.635 5.835 1770.805 ;
        RECT 6.125 1770.635 6.295 1770.805 ;
        RECT 6.585 1770.635 6.755 1770.805 ;
        RECT 2906.425 1770.635 2906.595 1770.805 ;
        RECT 2912.865 1770.635 2913.035 1770.805 ;
        RECT 2913.325 1770.635 2913.495 1770.805 ;
        RECT 2913.785 1770.635 2913.955 1770.805 ;
        RECT 5.665 1765.195 5.835 1765.365 ;
        RECT 6.125 1765.195 6.295 1765.365 ;
        RECT 6.585 1765.195 6.755 1765.365 ;
        RECT 2906.425 1765.195 2906.595 1765.365 ;
        RECT 2912.865 1765.195 2913.035 1765.365 ;
        RECT 2913.325 1765.195 2913.495 1765.365 ;
        RECT 2913.785 1765.195 2913.955 1765.365 ;
        RECT 5.665 1759.755 5.835 1759.925 ;
        RECT 6.125 1759.755 6.295 1759.925 ;
        RECT 6.585 1759.755 6.755 1759.925 ;
        RECT 2906.425 1759.755 2906.595 1759.925 ;
        RECT 2912.865 1759.755 2913.035 1759.925 ;
        RECT 2913.325 1759.755 2913.495 1759.925 ;
        RECT 2913.785 1759.755 2913.955 1759.925 ;
        RECT 5.665 1754.315 5.835 1754.485 ;
        RECT 6.125 1754.315 6.295 1754.485 ;
        RECT 6.585 1754.315 6.755 1754.485 ;
        RECT 2906.425 1754.315 2906.595 1754.485 ;
        RECT 2912.865 1754.315 2913.035 1754.485 ;
        RECT 2913.325 1754.315 2913.495 1754.485 ;
        RECT 2913.785 1754.315 2913.955 1754.485 ;
        RECT 5.665 1748.875 5.835 1749.045 ;
        RECT 6.125 1748.875 6.295 1749.045 ;
        RECT 6.585 1748.875 6.755 1749.045 ;
        RECT 2906.425 1748.875 2906.595 1749.045 ;
        RECT 2912.865 1748.875 2913.035 1749.045 ;
        RECT 2913.325 1748.875 2913.495 1749.045 ;
        RECT 2913.785 1748.875 2913.955 1749.045 ;
        RECT 5.665 1743.435 5.835 1743.605 ;
        RECT 6.125 1743.435 6.295 1743.605 ;
        RECT 6.585 1743.435 6.755 1743.605 ;
        RECT 2906.425 1743.435 2906.595 1743.605 ;
        RECT 2912.865 1743.435 2913.035 1743.605 ;
        RECT 2913.325 1743.435 2913.495 1743.605 ;
        RECT 2913.785 1743.435 2913.955 1743.605 ;
        RECT 5.665 1737.995 5.835 1738.165 ;
        RECT 6.125 1737.995 6.295 1738.165 ;
        RECT 6.585 1737.995 6.755 1738.165 ;
        RECT 2906.425 1737.995 2906.595 1738.165 ;
        RECT 2912.865 1737.995 2913.035 1738.165 ;
        RECT 2913.325 1737.995 2913.495 1738.165 ;
        RECT 2913.785 1737.995 2913.955 1738.165 ;
        RECT 5.665 1732.555 5.835 1732.725 ;
        RECT 6.125 1732.555 6.295 1732.725 ;
        RECT 6.585 1732.555 6.755 1732.725 ;
        RECT 2906.425 1732.555 2906.595 1732.725 ;
        RECT 2912.865 1732.555 2913.035 1732.725 ;
        RECT 2913.325 1732.555 2913.495 1732.725 ;
        RECT 2913.785 1732.555 2913.955 1732.725 ;
        RECT 5.665 1727.115 5.835 1727.285 ;
        RECT 6.125 1727.115 6.295 1727.285 ;
        RECT 6.585 1727.115 6.755 1727.285 ;
        RECT 2906.425 1727.115 2906.595 1727.285 ;
        RECT 2912.865 1727.115 2913.035 1727.285 ;
        RECT 2913.325 1727.115 2913.495 1727.285 ;
        RECT 2913.785 1727.115 2913.955 1727.285 ;
        RECT 5.665 1721.675 5.835 1721.845 ;
        RECT 6.125 1721.675 6.295 1721.845 ;
        RECT 6.585 1721.675 6.755 1721.845 ;
        RECT 2906.425 1721.675 2906.595 1721.845 ;
        RECT 2912.865 1721.675 2913.035 1721.845 ;
        RECT 2913.325 1721.675 2913.495 1721.845 ;
        RECT 2913.785 1721.675 2913.955 1721.845 ;
        RECT 5.665 1716.235 5.835 1716.405 ;
        RECT 6.125 1716.235 6.295 1716.405 ;
        RECT 6.585 1716.235 6.755 1716.405 ;
        RECT 2906.425 1716.235 2906.595 1716.405 ;
        RECT 2912.865 1716.235 2913.035 1716.405 ;
        RECT 2913.325 1716.235 2913.495 1716.405 ;
        RECT 2913.785 1716.235 2913.955 1716.405 ;
        RECT 5.665 1710.795 5.835 1710.965 ;
        RECT 6.125 1710.795 6.295 1710.965 ;
        RECT 6.585 1710.795 6.755 1710.965 ;
        RECT 2906.425 1710.795 2906.595 1710.965 ;
        RECT 2912.865 1710.795 2913.035 1710.965 ;
        RECT 2913.325 1710.795 2913.495 1710.965 ;
        RECT 2913.785 1710.795 2913.955 1710.965 ;
        RECT 5.665 1705.355 5.835 1705.525 ;
        RECT 6.125 1705.355 6.295 1705.525 ;
        RECT 6.585 1705.355 6.755 1705.525 ;
        RECT 8.885 1705.355 9.055 1705.525 ;
        RECT 9.345 1705.355 9.515 1705.525 ;
        RECT 9.805 1705.355 9.975 1705.525 ;
        RECT 2906.425 1705.355 2906.595 1705.525 ;
        RECT 2912.865 1705.355 2913.035 1705.525 ;
        RECT 2913.325 1705.355 2913.495 1705.525 ;
        RECT 2913.785 1705.355 2913.955 1705.525 ;
        RECT 5.665 1699.915 5.835 1700.085 ;
        RECT 6.125 1699.915 6.295 1700.085 ;
        RECT 6.585 1699.915 6.755 1700.085 ;
        RECT 2906.425 1699.915 2906.595 1700.085 ;
        RECT 2912.865 1699.915 2913.035 1700.085 ;
        RECT 2913.325 1699.915 2913.495 1700.085 ;
        RECT 2913.785 1699.915 2913.955 1700.085 ;
        RECT 5.665 1694.475 5.835 1694.645 ;
        RECT 6.125 1694.475 6.295 1694.645 ;
        RECT 6.585 1694.475 6.755 1694.645 ;
        RECT 2906.425 1694.475 2906.595 1694.645 ;
        RECT 2912.865 1694.475 2913.035 1694.645 ;
        RECT 2913.325 1694.475 2913.495 1694.645 ;
        RECT 2913.785 1694.475 2913.955 1694.645 ;
        RECT 5.665 1689.035 5.835 1689.205 ;
        RECT 6.125 1689.035 6.295 1689.205 ;
        RECT 6.585 1689.035 6.755 1689.205 ;
        RECT 2906.425 1689.035 2906.595 1689.205 ;
        RECT 2912.865 1689.035 2913.035 1689.205 ;
        RECT 2913.325 1689.035 2913.495 1689.205 ;
        RECT 2913.785 1689.035 2913.955 1689.205 ;
        RECT 5.665 1683.595 5.835 1683.765 ;
        RECT 6.125 1683.595 6.295 1683.765 ;
        RECT 6.585 1683.595 6.755 1683.765 ;
        RECT 2906.425 1683.595 2906.595 1683.765 ;
        RECT 2912.865 1683.595 2913.035 1683.765 ;
        RECT 2913.325 1683.595 2913.495 1683.765 ;
        RECT 2913.785 1683.595 2913.955 1683.765 ;
        RECT 5.665 1678.155 5.835 1678.325 ;
        RECT 6.125 1678.155 6.295 1678.325 ;
        RECT 6.585 1678.155 6.755 1678.325 ;
        RECT 2906.425 1678.155 2906.595 1678.325 ;
        RECT 2912.865 1678.155 2913.035 1678.325 ;
        RECT 2913.325 1678.155 2913.495 1678.325 ;
        RECT 2913.785 1678.155 2913.955 1678.325 ;
        RECT 5.665 1672.715 5.835 1672.885 ;
        RECT 6.125 1672.715 6.295 1672.885 ;
        RECT 6.585 1672.715 6.755 1672.885 ;
        RECT 2906.425 1672.715 2906.595 1672.885 ;
        RECT 2909.185 1672.715 2909.355 1672.885 ;
        RECT 2909.645 1672.715 2909.815 1672.885 ;
        RECT 2910.105 1672.715 2910.275 1672.885 ;
        RECT 2912.865 1672.715 2913.035 1672.885 ;
        RECT 2913.325 1672.715 2913.495 1672.885 ;
        RECT 2913.785 1672.715 2913.955 1672.885 ;
        RECT 5.665 1667.275 5.835 1667.445 ;
        RECT 6.125 1667.275 6.295 1667.445 ;
        RECT 6.585 1667.275 6.755 1667.445 ;
        RECT 2906.425 1667.275 2906.595 1667.445 ;
        RECT 2912.865 1667.275 2913.035 1667.445 ;
        RECT 2913.325 1667.275 2913.495 1667.445 ;
        RECT 2913.785 1667.275 2913.955 1667.445 ;
        RECT 5.665 1661.835 5.835 1662.005 ;
        RECT 6.125 1661.835 6.295 1662.005 ;
        RECT 6.585 1661.835 6.755 1662.005 ;
        RECT 2906.425 1661.835 2906.595 1662.005 ;
        RECT 2912.865 1661.835 2913.035 1662.005 ;
        RECT 2913.325 1661.835 2913.495 1662.005 ;
        RECT 2913.785 1661.835 2913.955 1662.005 ;
        RECT 5.665 1656.395 5.835 1656.565 ;
        RECT 6.125 1656.395 6.295 1656.565 ;
        RECT 6.585 1656.395 6.755 1656.565 ;
        RECT 2906.425 1656.395 2906.595 1656.565 ;
        RECT 2912.865 1656.395 2913.035 1656.565 ;
        RECT 2913.325 1656.395 2913.495 1656.565 ;
        RECT 2913.785 1656.395 2913.955 1656.565 ;
        RECT 5.665 1650.955 5.835 1651.125 ;
        RECT 6.125 1650.955 6.295 1651.125 ;
        RECT 6.585 1650.955 6.755 1651.125 ;
        RECT 2906.425 1650.955 2906.595 1651.125 ;
        RECT 2912.865 1650.955 2913.035 1651.125 ;
        RECT 2913.325 1650.955 2913.495 1651.125 ;
        RECT 2913.785 1650.955 2913.955 1651.125 ;
        RECT 5.665 1645.515 5.835 1645.685 ;
        RECT 6.125 1645.515 6.295 1645.685 ;
        RECT 6.585 1645.515 6.755 1645.685 ;
        RECT 2906.425 1645.515 2906.595 1645.685 ;
        RECT 2912.865 1645.515 2913.035 1645.685 ;
        RECT 2913.325 1645.515 2913.495 1645.685 ;
        RECT 2913.785 1645.515 2913.955 1645.685 ;
        RECT 5.665 1640.075 5.835 1640.245 ;
        RECT 6.125 1640.075 6.295 1640.245 ;
        RECT 6.585 1640.075 6.755 1640.245 ;
        RECT 2906.425 1640.075 2906.595 1640.245 ;
        RECT 2912.865 1640.075 2913.035 1640.245 ;
        RECT 2913.325 1640.075 2913.495 1640.245 ;
        RECT 2913.785 1640.075 2913.955 1640.245 ;
        RECT 5.665 1634.635 5.835 1634.805 ;
        RECT 6.125 1634.635 6.295 1634.805 ;
        RECT 6.585 1634.635 6.755 1634.805 ;
        RECT 2906.425 1634.635 2906.595 1634.805 ;
        RECT 2912.865 1634.635 2913.035 1634.805 ;
        RECT 2913.325 1634.635 2913.495 1634.805 ;
        RECT 2913.785 1634.635 2913.955 1634.805 ;
        RECT 5.665 1629.195 5.835 1629.365 ;
        RECT 6.125 1629.195 6.295 1629.365 ;
        RECT 6.585 1629.195 6.755 1629.365 ;
        RECT 2906.425 1629.195 2906.595 1629.365 ;
        RECT 2912.865 1629.195 2913.035 1629.365 ;
        RECT 2913.325 1629.195 2913.495 1629.365 ;
        RECT 2913.785 1629.195 2913.955 1629.365 ;
        RECT 5.665 1623.755 5.835 1623.925 ;
        RECT 6.125 1623.755 6.295 1623.925 ;
        RECT 6.585 1623.755 6.755 1623.925 ;
        RECT 2906.425 1623.755 2906.595 1623.925 ;
        RECT 2912.865 1623.755 2913.035 1623.925 ;
        RECT 2913.325 1623.755 2913.495 1623.925 ;
        RECT 2913.785 1623.755 2913.955 1623.925 ;
        RECT 5.665 1618.315 5.835 1618.485 ;
        RECT 6.125 1618.315 6.295 1618.485 ;
        RECT 6.585 1618.315 6.755 1618.485 ;
        RECT 2906.425 1618.315 2906.595 1618.485 ;
        RECT 2912.865 1618.315 2913.035 1618.485 ;
        RECT 2913.325 1618.315 2913.495 1618.485 ;
        RECT 2913.785 1618.315 2913.955 1618.485 ;
        RECT 5.665 1612.875 5.835 1613.045 ;
        RECT 6.125 1612.875 6.295 1613.045 ;
        RECT 6.585 1612.875 6.755 1613.045 ;
        RECT 2906.425 1612.875 2906.595 1613.045 ;
        RECT 2912.865 1612.875 2913.035 1613.045 ;
        RECT 2913.325 1612.875 2913.495 1613.045 ;
        RECT 2913.785 1612.875 2913.955 1613.045 ;
        RECT 5.665 1607.435 5.835 1607.605 ;
        RECT 6.125 1607.435 6.295 1607.605 ;
        RECT 6.585 1607.435 6.755 1607.605 ;
        RECT 2906.425 1607.435 2906.595 1607.605 ;
        RECT 2912.865 1607.435 2913.035 1607.605 ;
        RECT 2913.325 1607.435 2913.495 1607.605 ;
        RECT 2913.785 1607.435 2913.955 1607.605 ;
        RECT 5.665 1601.995 5.835 1602.165 ;
        RECT 6.125 1601.995 6.295 1602.165 ;
        RECT 6.585 1601.995 6.755 1602.165 ;
        RECT 2906.425 1601.995 2906.595 1602.165 ;
        RECT 2912.865 1601.995 2913.035 1602.165 ;
        RECT 2913.325 1601.995 2913.495 1602.165 ;
        RECT 2913.785 1601.995 2913.955 1602.165 ;
        RECT 5.665 1596.555 5.835 1596.725 ;
        RECT 6.125 1596.555 6.295 1596.725 ;
        RECT 6.585 1596.555 6.755 1596.725 ;
        RECT 2906.425 1596.555 2906.595 1596.725 ;
        RECT 2912.865 1596.555 2913.035 1596.725 ;
        RECT 2913.325 1596.555 2913.495 1596.725 ;
        RECT 2913.785 1596.555 2913.955 1596.725 ;
        RECT 5.665 1591.115 5.835 1591.285 ;
        RECT 6.125 1591.115 6.295 1591.285 ;
        RECT 6.585 1591.115 6.755 1591.285 ;
        RECT 2906.425 1591.115 2906.595 1591.285 ;
        RECT 2912.865 1591.115 2913.035 1591.285 ;
        RECT 2913.325 1591.115 2913.495 1591.285 ;
        RECT 2913.785 1591.115 2913.955 1591.285 ;
        RECT 5.665 1585.675 5.835 1585.845 ;
        RECT 6.125 1585.675 6.295 1585.845 ;
        RECT 6.585 1585.675 6.755 1585.845 ;
        RECT 2906.425 1585.675 2906.595 1585.845 ;
        RECT 2912.865 1585.675 2913.035 1585.845 ;
        RECT 2913.325 1585.675 2913.495 1585.845 ;
        RECT 2913.785 1585.675 2913.955 1585.845 ;
        RECT 5.665 1580.235 5.835 1580.405 ;
        RECT 6.125 1580.235 6.295 1580.405 ;
        RECT 6.585 1580.235 6.755 1580.405 ;
        RECT 8.885 1580.235 9.055 1580.405 ;
        RECT 9.345 1580.235 9.515 1580.405 ;
        RECT 9.805 1580.235 9.975 1580.405 ;
        RECT 2906.425 1580.235 2906.595 1580.405 ;
        RECT 2912.865 1580.235 2913.035 1580.405 ;
        RECT 2913.325 1580.235 2913.495 1580.405 ;
        RECT 2913.785 1580.235 2913.955 1580.405 ;
        RECT 5.665 1574.795 5.835 1574.965 ;
        RECT 6.125 1574.795 6.295 1574.965 ;
        RECT 6.585 1574.795 6.755 1574.965 ;
        RECT 2906.425 1574.795 2906.595 1574.965 ;
        RECT 2912.865 1574.795 2913.035 1574.965 ;
        RECT 2913.325 1574.795 2913.495 1574.965 ;
        RECT 2913.785 1574.795 2913.955 1574.965 ;
        RECT 5.665 1569.355 5.835 1569.525 ;
        RECT 6.125 1569.355 6.295 1569.525 ;
        RECT 6.585 1569.355 6.755 1569.525 ;
        RECT 2906.425 1569.355 2906.595 1569.525 ;
        RECT 2912.865 1569.355 2913.035 1569.525 ;
        RECT 2913.325 1569.355 2913.495 1569.525 ;
        RECT 2913.785 1569.355 2913.955 1569.525 ;
        RECT 5.665 1563.915 5.835 1564.085 ;
        RECT 6.125 1563.915 6.295 1564.085 ;
        RECT 6.585 1563.915 6.755 1564.085 ;
        RECT 2906.425 1563.915 2906.595 1564.085 ;
        RECT 2912.865 1563.915 2913.035 1564.085 ;
        RECT 2913.325 1563.915 2913.495 1564.085 ;
        RECT 2913.785 1563.915 2913.955 1564.085 ;
        RECT 5.665 1558.475 5.835 1558.645 ;
        RECT 6.125 1558.475 6.295 1558.645 ;
        RECT 6.585 1558.475 6.755 1558.645 ;
        RECT 2906.425 1558.475 2906.595 1558.645 ;
        RECT 2912.865 1558.475 2913.035 1558.645 ;
        RECT 2913.325 1558.475 2913.495 1558.645 ;
        RECT 2913.785 1558.475 2913.955 1558.645 ;
        RECT 5.665 1553.035 5.835 1553.205 ;
        RECT 6.125 1553.035 6.295 1553.205 ;
        RECT 6.585 1553.035 6.755 1553.205 ;
        RECT 2906.425 1553.035 2906.595 1553.205 ;
        RECT 2912.865 1553.035 2913.035 1553.205 ;
        RECT 2913.325 1553.035 2913.495 1553.205 ;
        RECT 2913.785 1553.035 2913.955 1553.205 ;
        RECT 5.665 1547.595 5.835 1547.765 ;
        RECT 6.125 1547.595 6.295 1547.765 ;
        RECT 6.585 1547.595 6.755 1547.765 ;
        RECT 2906.425 1547.595 2906.595 1547.765 ;
        RECT 2912.865 1547.595 2913.035 1547.765 ;
        RECT 2913.325 1547.595 2913.495 1547.765 ;
        RECT 2913.785 1547.595 2913.955 1547.765 ;
        RECT 5.665 1542.155 5.835 1542.325 ;
        RECT 6.125 1542.155 6.295 1542.325 ;
        RECT 6.585 1542.155 6.755 1542.325 ;
        RECT 2906.425 1542.155 2906.595 1542.325 ;
        RECT 2912.865 1542.155 2913.035 1542.325 ;
        RECT 2913.325 1542.155 2913.495 1542.325 ;
        RECT 2913.785 1542.155 2913.955 1542.325 ;
        RECT 5.665 1536.715 5.835 1536.885 ;
        RECT 6.125 1536.715 6.295 1536.885 ;
        RECT 6.585 1536.715 6.755 1536.885 ;
        RECT 2906.425 1536.715 2906.595 1536.885 ;
        RECT 2912.865 1536.715 2913.035 1536.885 ;
        RECT 2913.325 1536.715 2913.495 1536.885 ;
        RECT 2913.785 1536.715 2913.955 1536.885 ;
        RECT 5.665 1531.275 5.835 1531.445 ;
        RECT 6.125 1531.275 6.295 1531.445 ;
        RECT 6.585 1531.275 6.755 1531.445 ;
        RECT 2906.425 1531.275 2906.595 1531.445 ;
        RECT 2912.865 1531.275 2913.035 1531.445 ;
        RECT 2913.325 1531.275 2913.495 1531.445 ;
        RECT 2913.785 1531.275 2913.955 1531.445 ;
        RECT 5.665 1525.835 5.835 1526.005 ;
        RECT 6.125 1525.835 6.295 1526.005 ;
        RECT 6.585 1525.835 6.755 1526.005 ;
        RECT 2906.425 1525.835 2906.595 1526.005 ;
        RECT 2909.185 1525.835 2909.355 1526.005 ;
        RECT 2909.645 1525.835 2909.815 1526.005 ;
        RECT 2910.105 1525.835 2910.275 1526.005 ;
        RECT 2912.865 1525.835 2913.035 1526.005 ;
        RECT 2913.325 1525.835 2913.495 1526.005 ;
        RECT 2913.785 1525.835 2913.955 1526.005 ;
        RECT 5.665 1520.395 5.835 1520.565 ;
        RECT 6.125 1520.395 6.295 1520.565 ;
        RECT 6.585 1520.395 6.755 1520.565 ;
        RECT 2906.425 1520.395 2906.595 1520.565 ;
        RECT 2912.865 1520.395 2913.035 1520.565 ;
        RECT 2913.325 1520.395 2913.495 1520.565 ;
        RECT 2913.785 1520.395 2913.955 1520.565 ;
        RECT 5.665 1514.955 5.835 1515.125 ;
        RECT 6.125 1514.955 6.295 1515.125 ;
        RECT 6.585 1514.955 6.755 1515.125 ;
        RECT 2906.425 1514.955 2906.595 1515.125 ;
        RECT 2909.185 1514.955 2909.355 1515.125 ;
        RECT 2909.645 1514.955 2909.815 1515.125 ;
        RECT 2910.105 1514.955 2910.275 1515.125 ;
        RECT 2912.865 1514.955 2913.035 1515.125 ;
        RECT 2913.325 1514.955 2913.495 1515.125 ;
        RECT 2913.785 1514.955 2913.955 1515.125 ;
        RECT 5.665 1509.515 5.835 1509.685 ;
        RECT 6.125 1509.515 6.295 1509.685 ;
        RECT 6.585 1509.515 6.755 1509.685 ;
        RECT 2906.425 1509.515 2906.595 1509.685 ;
        RECT 2912.865 1509.515 2913.035 1509.685 ;
        RECT 2913.325 1509.515 2913.495 1509.685 ;
        RECT 2913.785 1509.515 2913.955 1509.685 ;
        RECT 5.665 1504.075 5.835 1504.245 ;
        RECT 6.125 1504.075 6.295 1504.245 ;
        RECT 6.585 1504.075 6.755 1504.245 ;
        RECT 2906.425 1504.075 2906.595 1504.245 ;
        RECT 2912.865 1504.075 2913.035 1504.245 ;
        RECT 2913.325 1504.075 2913.495 1504.245 ;
        RECT 2913.785 1504.075 2913.955 1504.245 ;
        RECT 5.665 1498.635 5.835 1498.805 ;
        RECT 6.125 1498.635 6.295 1498.805 ;
        RECT 6.585 1498.635 6.755 1498.805 ;
        RECT 2906.425 1498.635 2906.595 1498.805 ;
        RECT 2912.865 1498.635 2913.035 1498.805 ;
        RECT 2913.325 1498.635 2913.495 1498.805 ;
        RECT 2913.785 1498.635 2913.955 1498.805 ;
        RECT 5.665 1493.195 5.835 1493.365 ;
        RECT 6.125 1493.195 6.295 1493.365 ;
        RECT 6.585 1493.195 6.755 1493.365 ;
        RECT 2906.425 1493.195 2906.595 1493.365 ;
        RECT 2912.865 1493.195 2913.035 1493.365 ;
        RECT 2913.325 1493.195 2913.495 1493.365 ;
        RECT 2913.785 1493.195 2913.955 1493.365 ;
        RECT 5.665 1487.755 5.835 1487.925 ;
        RECT 6.125 1487.755 6.295 1487.925 ;
        RECT 6.585 1487.755 6.755 1487.925 ;
        RECT 2906.425 1487.755 2906.595 1487.925 ;
        RECT 2912.865 1487.755 2913.035 1487.925 ;
        RECT 2913.325 1487.755 2913.495 1487.925 ;
        RECT 2913.785 1487.755 2913.955 1487.925 ;
        RECT 5.665 1482.315 5.835 1482.485 ;
        RECT 6.125 1482.315 6.295 1482.485 ;
        RECT 6.585 1482.315 6.755 1482.485 ;
        RECT 2906.425 1482.315 2906.595 1482.485 ;
        RECT 2912.865 1482.315 2913.035 1482.485 ;
        RECT 2913.325 1482.315 2913.495 1482.485 ;
        RECT 2913.785 1482.315 2913.955 1482.485 ;
        RECT 5.665 1476.875 5.835 1477.045 ;
        RECT 6.125 1476.875 6.295 1477.045 ;
        RECT 6.585 1476.875 6.755 1477.045 ;
        RECT 2906.425 1476.875 2906.595 1477.045 ;
        RECT 2912.865 1476.875 2913.035 1477.045 ;
        RECT 2913.325 1476.875 2913.495 1477.045 ;
        RECT 2913.785 1476.875 2913.955 1477.045 ;
        RECT 5.665 1471.435 5.835 1471.605 ;
        RECT 6.125 1471.435 6.295 1471.605 ;
        RECT 6.585 1471.435 6.755 1471.605 ;
        RECT 2906.425 1471.435 2906.595 1471.605 ;
        RECT 2909.185 1471.435 2909.355 1471.605 ;
        RECT 2909.645 1471.435 2909.815 1471.605 ;
        RECT 2910.105 1471.435 2910.275 1471.605 ;
        RECT 2912.865 1471.435 2913.035 1471.605 ;
        RECT 2913.325 1471.435 2913.495 1471.605 ;
        RECT 2913.785 1471.435 2913.955 1471.605 ;
        RECT 5.665 1465.995 5.835 1466.165 ;
        RECT 6.125 1465.995 6.295 1466.165 ;
        RECT 6.585 1465.995 6.755 1466.165 ;
        RECT 2906.425 1465.995 2906.595 1466.165 ;
        RECT 2912.865 1465.995 2913.035 1466.165 ;
        RECT 2913.325 1465.995 2913.495 1466.165 ;
        RECT 2913.785 1465.995 2913.955 1466.165 ;
        RECT 5.665 1460.555 5.835 1460.725 ;
        RECT 6.125 1460.555 6.295 1460.725 ;
        RECT 6.585 1460.555 6.755 1460.725 ;
        RECT 2906.425 1460.555 2906.595 1460.725 ;
        RECT 2912.865 1460.555 2913.035 1460.725 ;
        RECT 2913.325 1460.555 2913.495 1460.725 ;
        RECT 2913.785 1460.555 2913.955 1460.725 ;
        RECT 5.665 1455.115 5.835 1455.285 ;
        RECT 6.125 1455.115 6.295 1455.285 ;
        RECT 6.585 1455.115 6.755 1455.285 ;
        RECT 2906.425 1455.115 2906.595 1455.285 ;
        RECT 2912.865 1455.115 2913.035 1455.285 ;
        RECT 2913.325 1455.115 2913.495 1455.285 ;
        RECT 2913.785 1455.115 2913.955 1455.285 ;
        RECT 5.665 1449.675 5.835 1449.845 ;
        RECT 6.125 1449.675 6.295 1449.845 ;
        RECT 6.585 1449.675 6.755 1449.845 ;
        RECT 2906.425 1449.675 2906.595 1449.845 ;
        RECT 2912.865 1449.675 2913.035 1449.845 ;
        RECT 2913.325 1449.675 2913.495 1449.845 ;
        RECT 2913.785 1449.675 2913.955 1449.845 ;
        RECT 5.665 1444.235 5.835 1444.405 ;
        RECT 6.125 1444.235 6.295 1444.405 ;
        RECT 6.585 1444.235 6.755 1444.405 ;
        RECT 2906.425 1444.235 2906.595 1444.405 ;
        RECT 2912.865 1444.235 2913.035 1444.405 ;
        RECT 2913.325 1444.235 2913.495 1444.405 ;
        RECT 2913.785 1444.235 2913.955 1444.405 ;
        RECT 5.665 1438.795 5.835 1438.965 ;
        RECT 6.125 1438.795 6.295 1438.965 ;
        RECT 6.585 1438.795 6.755 1438.965 ;
        RECT 2906.425 1438.795 2906.595 1438.965 ;
        RECT 2912.865 1438.795 2913.035 1438.965 ;
        RECT 2913.325 1438.795 2913.495 1438.965 ;
        RECT 2913.785 1438.795 2913.955 1438.965 ;
        RECT 5.665 1433.355 5.835 1433.525 ;
        RECT 6.125 1433.355 6.295 1433.525 ;
        RECT 6.585 1433.355 6.755 1433.525 ;
        RECT 2906.425 1433.355 2906.595 1433.525 ;
        RECT 2912.865 1433.355 2913.035 1433.525 ;
        RECT 2913.325 1433.355 2913.495 1433.525 ;
        RECT 2913.785 1433.355 2913.955 1433.525 ;
        RECT 5.665 1427.915 5.835 1428.085 ;
        RECT 6.125 1427.915 6.295 1428.085 ;
        RECT 6.585 1427.915 6.755 1428.085 ;
        RECT 2906.425 1427.915 2906.595 1428.085 ;
        RECT 2912.865 1427.915 2913.035 1428.085 ;
        RECT 2913.325 1427.915 2913.495 1428.085 ;
        RECT 2913.785 1427.915 2913.955 1428.085 ;
        RECT 5.665 1422.475 5.835 1422.645 ;
        RECT 6.125 1422.475 6.295 1422.645 ;
        RECT 6.585 1422.475 6.755 1422.645 ;
        RECT 2906.425 1422.475 2906.595 1422.645 ;
        RECT 2912.865 1422.475 2913.035 1422.645 ;
        RECT 2913.325 1422.475 2913.495 1422.645 ;
        RECT 2913.785 1422.475 2913.955 1422.645 ;
        RECT 5.665 1417.035 5.835 1417.205 ;
        RECT 6.125 1417.035 6.295 1417.205 ;
        RECT 6.585 1417.035 6.755 1417.205 ;
        RECT 2906.425 1417.035 2906.595 1417.205 ;
        RECT 2912.865 1417.035 2913.035 1417.205 ;
        RECT 2913.325 1417.035 2913.495 1417.205 ;
        RECT 2913.785 1417.035 2913.955 1417.205 ;
        RECT 5.665 1411.595 5.835 1411.765 ;
        RECT 6.125 1411.595 6.295 1411.765 ;
        RECT 6.585 1411.595 6.755 1411.765 ;
        RECT 2906.425 1411.595 2906.595 1411.765 ;
        RECT 2912.865 1411.595 2913.035 1411.765 ;
        RECT 2913.325 1411.595 2913.495 1411.765 ;
        RECT 2913.785 1411.595 2913.955 1411.765 ;
        RECT 5.665 1406.155 5.835 1406.325 ;
        RECT 6.125 1406.155 6.295 1406.325 ;
        RECT 6.585 1406.155 6.755 1406.325 ;
        RECT 2906.425 1406.155 2906.595 1406.325 ;
        RECT 2912.865 1406.155 2913.035 1406.325 ;
        RECT 2913.325 1406.155 2913.495 1406.325 ;
        RECT 2913.785 1406.155 2913.955 1406.325 ;
        RECT 5.665 1400.715 5.835 1400.885 ;
        RECT 6.125 1400.715 6.295 1400.885 ;
        RECT 6.585 1400.715 6.755 1400.885 ;
        RECT 2906.425 1400.715 2906.595 1400.885 ;
        RECT 2912.865 1400.715 2913.035 1400.885 ;
        RECT 2913.325 1400.715 2913.495 1400.885 ;
        RECT 2913.785 1400.715 2913.955 1400.885 ;
        RECT 5.665 1395.275 5.835 1395.445 ;
        RECT 6.125 1395.275 6.295 1395.445 ;
        RECT 6.585 1395.275 6.755 1395.445 ;
        RECT 2906.425 1395.275 2906.595 1395.445 ;
        RECT 2912.865 1395.275 2913.035 1395.445 ;
        RECT 2913.325 1395.275 2913.495 1395.445 ;
        RECT 2913.785 1395.275 2913.955 1395.445 ;
        RECT 5.665 1389.835 5.835 1390.005 ;
        RECT 6.125 1389.835 6.295 1390.005 ;
        RECT 6.585 1389.835 6.755 1390.005 ;
        RECT 2906.425 1389.835 2906.595 1390.005 ;
        RECT 2912.865 1389.835 2913.035 1390.005 ;
        RECT 2913.325 1389.835 2913.495 1390.005 ;
        RECT 2913.785 1389.835 2913.955 1390.005 ;
        RECT 5.665 1384.395 5.835 1384.565 ;
        RECT 6.125 1384.395 6.295 1384.565 ;
        RECT 6.585 1384.395 6.755 1384.565 ;
        RECT 2906.425 1384.395 2906.595 1384.565 ;
        RECT 2912.865 1384.395 2913.035 1384.565 ;
        RECT 2913.325 1384.395 2913.495 1384.565 ;
        RECT 2913.785 1384.395 2913.955 1384.565 ;
        RECT 5.665 1378.955 5.835 1379.125 ;
        RECT 6.125 1378.955 6.295 1379.125 ;
        RECT 6.585 1378.955 6.755 1379.125 ;
        RECT 2906.425 1378.955 2906.595 1379.125 ;
        RECT 2912.865 1378.955 2913.035 1379.125 ;
        RECT 2913.325 1378.955 2913.495 1379.125 ;
        RECT 2913.785 1378.955 2913.955 1379.125 ;
        RECT 5.665 1373.515 5.835 1373.685 ;
        RECT 6.125 1373.515 6.295 1373.685 ;
        RECT 6.585 1373.515 6.755 1373.685 ;
        RECT 2906.425 1373.515 2906.595 1373.685 ;
        RECT 2912.865 1373.515 2913.035 1373.685 ;
        RECT 2913.325 1373.515 2913.495 1373.685 ;
        RECT 2913.785 1373.515 2913.955 1373.685 ;
        RECT 5.665 1368.075 5.835 1368.245 ;
        RECT 6.125 1368.075 6.295 1368.245 ;
        RECT 6.585 1368.075 6.755 1368.245 ;
        RECT 2906.425 1368.075 2906.595 1368.245 ;
        RECT 2912.865 1368.075 2913.035 1368.245 ;
        RECT 2913.325 1368.075 2913.495 1368.245 ;
        RECT 2913.785 1368.075 2913.955 1368.245 ;
        RECT 5.665 1362.635 5.835 1362.805 ;
        RECT 6.125 1362.635 6.295 1362.805 ;
        RECT 6.585 1362.635 6.755 1362.805 ;
        RECT 2906.425 1362.635 2906.595 1362.805 ;
        RECT 2912.865 1362.635 2913.035 1362.805 ;
        RECT 2913.325 1362.635 2913.495 1362.805 ;
        RECT 2913.785 1362.635 2913.955 1362.805 ;
        RECT 5.665 1357.195 5.835 1357.365 ;
        RECT 6.125 1357.195 6.295 1357.365 ;
        RECT 6.585 1357.195 6.755 1357.365 ;
        RECT 2906.425 1357.195 2906.595 1357.365 ;
        RECT 2912.865 1357.195 2913.035 1357.365 ;
        RECT 2913.325 1357.195 2913.495 1357.365 ;
        RECT 2913.785 1357.195 2913.955 1357.365 ;
        RECT 5.665 1351.755 5.835 1351.925 ;
        RECT 6.125 1351.755 6.295 1351.925 ;
        RECT 6.585 1351.755 6.755 1351.925 ;
        RECT 2906.425 1351.755 2906.595 1351.925 ;
        RECT 2912.865 1351.755 2913.035 1351.925 ;
        RECT 2913.325 1351.755 2913.495 1351.925 ;
        RECT 2913.785 1351.755 2913.955 1351.925 ;
        RECT 5.665 1346.315 5.835 1346.485 ;
        RECT 6.125 1346.315 6.295 1346.485 ;
        RECT 6.585 1346.315 6.755 1346.485 ;
        RECT 2906.425 1346.315 2906.595 1346.485 ;
        RECT 2912.865 1346.315 2913.035 1346.485 ;
        RECT 2913.325 1346.315 2913.495 1346.485 ;
        RECT 2913.785 1346.315 2913.955 1346.485 ;
        RECT 5.665 1340.875 5.835 1341.045 ;
        RECT 6.125 1340.875 6.295 1341.045 ;
        RECT 6.585 1340.875 6.755 1341.045 ;
        RECT 2906.425 1340.875 2906.595 1341.045 ;
        RECT 2912.865 1340.875 2913.035 1341.045 ;
        RECT 2913.325 1340.875 2913.495 1341.045 ;
        RECT 2913.785 1340.875 2913.955 1341.045 ;
        RECT 5.665 1335.435 5.835 1335.605 ;
        RECT 6.125 1335.435 6.295 1335.605 ;
        RECT 6.585 1335.435 6.755 1335.605 ;
        RECT 2906.425 1335.435 2906.595 1335.605 ;
        RECT 2912.865 1335.435 2913.035 1335.605 ;
        RECT 2913.325 1335.435 2913.495 1335.605 ;
        RECT 2913.785 1335.435 2913.955 1335.605 ;
        RECT 5.665 1329.995 5.835 1330.165 ;
        RECT 6.125 1329.995 6.295 1330.165 ;
        RECT 6.585 1329.995 6.755 1330.165 ;
        RECT 8.885 1329.995 9.055 1330.165 ;
        RECT 9.345 1329.995 9.515 1330.165 ;
        RECT 9.805 1329.995 9.975 1330.165 ;
        RECT 2906.425 1329.995 2906.595 1330.165 ;
        RECT 2912.865 1329.995 2913.035 1330.165 ;
        RECT 2913.325 1329.995 2913.495 1330.165 ;
        RECT 2913.785 1329.995 2913.955 1330.165 ;
        RECT 5.665 1324.555 5.835 1324.725 ;
        RECT 6.125 1324.555 6.295 1324.725 ;
        RECT 6.585 1324.555 6.755 1324.725 ;
        RECT 2906.425 1324.555 2906.595 1324.725 ;
        RECT 2912.865 1324.555 2913.035 1324.725 ;
        RECT 2913.325 1324.555 2913.495 1324.725 ;
        RECT 2913.785 1324.555 2913.955 1324.725 ;
        RECT 5.665 1319.115 5.835 1319.285 ;
        RECT 6.125 1319.115 6.295 1319.285 ;
        RECT 6.585 1319.115 6.755 1319.285 ;
        RECT 2906.425 1319.115 2906.595 1319.285 ;
        RECT 2912.865 1319.115 2913.035 1319.285 ;
        RECT 2913.325 1319.115 2913.495 1319.285 ;
        RECT 2913.785 1319.115 2913.955 1319.285 ;
        RECT 5.665 1313.675 5.835 1313.845 ;
        RECT 6.125 1313.675 6.295 1313.845 ;
        RECT 6.585 1313.675 6.755 1313.845 ;
        RECT 2906.425 1313.675 2906.595 1313.845 ;
        RECT 2912.865 1313.675 2913.035 1313.845 ;
        RECT 2913.325 1313.675 2913.495 1313.845 ;
        RECT 2913.785 1313.675 2913.955 1313.845 ;
        RECT 5.665 1308.235 5.835 1308.405 ;
        RECT 6.125 1308.235 6.295 1308.405 ;
        RECT 6.585 1308.235 6.755 1308.405 ;
        RECT 2906.425 1308.235 2906.595 1308.405 ;
        RECT 2912.865 1308.235 2913.035 1308.405 ;
        RECT 2913.325 1308.235 2913.495 1308.405 ;
        RECT 2913.785 1308.235 2913.955 1308.405 ;
        RECT 5.665 1302.795 5.835 1302.965 ;
        RECT 6.125 1302.795 6.295 1302.965 ;
        RECT 6.585 1302.795 6.755 1302.965 ;
        RECT 2906.425 1302.795 2906.595 1302.965 ;
        RECT 2909.185 1302.795 2909.355 1302.965 ;
        RECT 2909.645 1302.795 2909.815 1302.965 ;
        RECT 2910.105 1302.795 2910.275 1302.965 ;
        RECT 2912.865 1302.795 2913.035 1302.965 ;
        RECT 2913.325 1302.795 2913.495 1302.965 ;
        RECT 2913.785 1302.795 2913.955 1302.965 ;
        RECT 5.665 1297.355 5.835 1297.525 ;
        RECT 6.125 1297.355 6.295 1297.525 ;
        RECT 6.585 1297.355 6.755 1297.525 ;
        RECT 2906.425 1297.355 2906.595 1297.525 ;
        RECT 2912.865 1297.355 2913.035 1297.525 ;
        RECT 2913.325 1297.355 2913.495 1297.525 ;
        RECT 2913.785 1297.355 2913.955 1297.525 ;
        RECT 5.665 1291.915 5.835 1292.085 ;
        RECT 6.125 1291.915 6.295 1292.085 ;
        RECT 6.585 1291.915 6.755 1292.085 ;
        RECT 2906.425 1291.915 2906.595 1292.085 ;
        RECT 2912.865 1291.915 2913.035 1292.085 ;
        RECT 2913.325 1291.915 2913.495 1292.085 ;
        RECT 2913.785 1291.915 2913.955 1292.085 ;
        RECT 5.665 1286.475 5.835 1286.645 ;
        RECT 6.125 1286.475 6.295 1286.645 ;
        RECT 6.585 1286.475 6.755 1286.645 ;
        RECT 8.885 1286.475 9.055 1286.645 ;
        RECT 9.345 1286.475 9.515 1286.645 ;
        RECT 9.805 1286.475 9.975 1286.645 ;
        RECT 2906.425 1286.475 2906.595 1286.645 ;
        RECT 2912.865 1286.475 2913.035 1286.645 ;
        RECT 2913.325 1286.475 2913.495 1286.645 ;
        RECT 2913.785 1286.475 2913.955 1286.645 ;
        RECT 5.665 1281.035 5.835 1281.205 ;
        RECT 6.125 1281.035 6.295 1281.205 ;
        RECT 6.585 1281.035 6.755 1281.205 ;
        RECT 2906.425 1281.035 2906.595 1281.205 ;
        RECT 2912.865 1281.035 2913.035 1281.205 ;
        RECT 2913.325 1281.035 2913.495 1281.205 ;
        RECT 2913.785 1281.035 2913.955 1281.205 ;
        RECT 5.665 1275.595 5.835 1275.765 ;
        RECT 6.125 1275.595 6.295 1275.765 ;
        RECT 6.585 1275.595 6.755 1275.765 ;
        RECT 8.885 1275.595 9.055 1275.765 ;
        RECT 9.345 1275.595 9.515 1275.765 ;
        RECT 9.805 1275.595 9.975 1275.765 ;
        RECT 2906.425 1275.595 2906.595 1275.765 ;
        RECT 2912.865 1275.595 2913.035 1275.765 ;
        RECT 2913.325 1275.595 2913.495 1275.765 ;
        RECT 2913.785 1275.595 2913.955 1275.765 ;
        RECT 5.665 1270.155 5.835 1270.325 ;
        RECT 6.125 1270.155 6.295 1270.325 ;
        RECT 6.585 1270.155 6.755 1270.325 ;
        RECT 2906.425 1270.155 2906.595 1270.325 ;
        RECT 2912.865 1270.155 2913.035 1270.325 ;
        RECT 2913.325 1270.155 2913.495 1270.325 ;
        RECT 2913.785 1270.155 2913.955 1270.325 ;
        RECT 5.665 1264.715 5.835 1264.885 ;
        RECT 6.125 1264.715 6.295 1264.885 ;
        RECT 6.585 1264.715 6.755 1264.885 ;
        RECT 2906.425 1264.715 2906.595 1264.885 ;
        RECT 2909.185 1264.715 2909.355 1264.885 ;
        RECT 2909.645 1264.715 2909.815 1264.885 ;
        RECT 2910.105 1264.715 2910.275 1264.885 ;
        RECT 2912.865 1264.715 2913.035 1264.885 ;
        RECT 2913.325 1264.715 2913.495 1264.885 ;
        RECT 2913.785 1264.715 2913.955 1264.885 ;
        RECT 5.665 1259.275 5.835 1259.445 ;
        RECT 6.125 1259.275 6.295 1259.445 ;
        RECT 6.585 1259.275 6.755 1259.445 ;
        RECT 2906.425 1259.275 2906.595 1259.445 ;
        RECT 2912.865 1259.275 2913.035 1259.445 ;
        RECT 2913.325 1259.275 2913.495 1259.445 ;
        RECT 2913.785 1259.275 2913.955 1259.445 ;
        RECT 5.665 1253.835 5.835 1254.005 ;
        RECT 6.125 1253.835 6.295 1254.005 ;
        RECT 6.585 1253.835 6.755 1254.005 ;
        RECT 2906.425 1253.835 2906.595 1254.005 ;
        RECT 2912.865 1253.835 2913.035 1254.005 ;
        RECT 2913.325 1253.835 2913.495 1254.005 ;
        RECT 2913.785 1253.835 2913.955 1254.005 ;
        RECT 5.665 1248.395 5.835 1248.565 ;
        RECT 6.125 1248.395 6.295 1248.565 ;
        RECT 6.585 1248.395 6.755 1248.565 ;
        RECT 2906.425 1248.395 2906.595 1248.565 ;
        RECT 2912.865 1248.395 2913.035 1248.565 ;
        RECT 2913.325 1248.395 2913.495 1248.565 ;
        RECT 2913.785 1248.395 2913.955 1248.565 ;
        RECT 5.665 1242.955 5.835 1243.125 ;
        RECT 6.125 1242.955 6.295 1243.125 ;
        RECT 6.585 1242.955 6.755 1243.125 ;
        RECT 2912.865 1242.955 2913.035 1243.125 ;
        RECT 2913.325 1242.955 2913.495 1243.125 ;
        RECT 2913.785 1242.955 2913.955 1243.125 ;
        RECT 5.665 1237.515 5.835 1237.685 ;
        RECT 6.125 1237.515 6.295 1237.685 ;
        RECT 6.585 1237.515 6.755 1237.685 ;
        RECT 2910.105 1237.515 2910.275 1237.685 ;
        RECT 2912.865 1237.515 2913.035 1237.685 ;
        RECT 2913.325 1237.515 2913.495 1237.685 ;
        RECT 2913.785 1237.515 2913.955 1237.685 ;
        RECT 5.665 1232.075 5.835 1232.245 ;
        RECT 6.125 1232.075 6.295 1232.245 ;
        RECT 6.585 1232.075 6.755 1232.245 ;
        RECT 2910.105 1232.075 2910.275 1232.245 ;
        RECT 2912.865 1232.075 2913.035 1232.245 ;
        RECT 2913.325 1232.075 2913.495 1232.245 ;
        RECT 2913.785 1232.075 2913.955 1232.245 ;
        RECT 5.665 1226.635 5.835 1226.805 ;
        RECT 6.125 1226.635 6.295 1226.805 ;
        RECT 6.585 1226.635 6.755 1226.805 ;
        RECT 2910.105 1226.635 2910.275 1226.805 ;
        RECT 2912.865 1226.635 2913.035 1226.805 ;
        RECT 2913.325 1226.635 2913.495 1226.805 ;
        RECT 2913.785 1226.635 2913.955 1226.805 ;
        RECT 5.665 1221.195 5.835 1221.365 ;
        RECT 6.125 1221.195 6.295 1221.365 ;
        RECT 6.585 1221.195 6.755 1221.365 ;
        RECT 2910.105 1221.195 2910.275 1221.365 ;
        RECT 2912.865 1221.195 2913.035 1221.365 ;
        RECT 2913.325 1221.195 2913.495 1221.365 ;
        RECT 2913.785 1221.195 2913.955 1221.365 ;
        RECT 5.665 1215.755 5.835 1215.925 ;
        RECT 6.125 1215.755 6.295 1215.925 ;
        RECT 6.585 1215.755 6.755 1215.925 ;
        RECT 8.885 1215.755 9.055 1215.925 ;
        RECT 9.345 1215.755 9.515 1215.925 ;
        RECT 9.805 1215.755 9.975 1215.925 ;
        RECT 2910.105 1215.755 2910.275 1215.925 ;
        RECT 2912.865 1215.755 2913.035 1215.925 ;
        RECT 2913.325 1215.755 2913.495 1215.925 ;
        RECT 2913.785 1215.755 2913.955 1215.925 ;
        RECT 5.665 1210.315 5.835 1210.485 ;
        RECT 6.125 1210.315 6.295 1210.485 ;
        RECT 6.585 1210.315 6.755 1210.485 ;
        RECT 2910.105 1210.315 2910.275 1210.485 ;
        RECT 2912.865 1210.315 2913.035 1210.485 ;
        RECT 2913.325 1210.315 2913.495 1210.485 ;
        RECT 2913.785 1210.315 2913.955 1210.485 ;
        RECT 5.665 1204.875 5.835 1205.045 ;
        RECT 6.125 1204.875 6.295 1205.045 ;
        RECT 6.585 1204.875 6.755 1205.045 ;
        RECT 2910.105 1204.875 2910.275 1205.045 ;
        RECT 2912.865 1204.875 2913.035 1205.045 ;
        RECT 2913.325 1204.875 2913.495 1205.045 ;
        RECT 2913.785 1204.875 2913.955 1205.045 ;
        RECT 5.665 1199.435 5.835 1199.605 ;
        RECT 6.125 1199.435 6.295 1199.605 ;
        RECT 6.585 1199.435 6.755 1199.605 ;
        RECT 2910.105 1199.435 2910.275 1199.605 ;
        RECT 2912.865 1199.435 2913.035 1199.605 ;
        RECT 2913.325 1199.435 2913.495 1199.605 ;
        RECT 2913.785 1199.435 2913.955 1199.605 ;
        RECT 5.665 1193.995 5.835 1194.165 ;
        RECT 6.125 1193.995 6.295 1194.165 ;
        RECT 6.585 1193.995 6.755 1194.165 ;
        RECT 2910.105 1193.995 2910.275 1194.165 ;
        RECT 2912.865 1193.995 2913.035 1194.165 ;
        RECT 2913.325 1193.995 2913.495 1194.165 ;
        RECT 2913.785 1193.995 2913.955 1194.165 ;
        RECT 5.665 1188.555 5.835 1188.725 ;
        RECT 6.125 1188.555 6.295 1188.725 ;
        RECT 6.585 1188.555 6.755 1188.725 ;
        RECT 2910.105 1188.555 2910.275 1188.725 ;
        RECT 2912.865 1188.555 2913.035 1188.725 ;
        RECT 2913.325 1188.555 2913.495 1188.725 ;
        RECT 2913.785 1188.555 2913.955 1188.725 ;
        RECT 5.665 1183.115 5.835 1183.285 ;
        RECT 6.125 1183.115 6.295 1183.285 ;
        RECT 6.585 1183.115 6.755 1183.285 ;
        RECT 2910.105 1183.115 2910.275 1183.285 ;
        RECT 2912.865 1183.115 2913.035 1183.285 ;
        RECT 2913.325 1183.115 2913.495 1183.285 ;
        RECT 2913.785 1183.115 2913.955 1183.285 ;
        RECT 5.665 1177.675 5.835 1177.845 ;
        RECT 6.125 1177.675 6.295 1177.845 ;
        RECT 6.585 1177.675 6.755 1177.845 ;
        RECT 2910.105 1177.675 2910.275 1177.845 ;
        RECT 2912.865 1177.675 2913.035 1177.845 ;
        RECT 2913.325 1177.675 2913.495 1177.845 ;
        RECT 2913.785 1177.675 2913.955 1177.845 ;
        RECT 5.665 1172.235 5.835 1172.405 ;
        RECT 6.125 1172.235 6.295 1172.405 ;
        RECT 6.585 1172.235 6.755 1172.405 ;
        RECT 2910.105 1172.235 2910.275 1172.405 ;
        RECT 2912.865 1172.235 2913.035 1172.405 ;
        RECT 2913.325 1172.235 2913.495 1172.405 ;
        RECT 2913.785 1172.235 2913.955 1172.405 ;
        RECT 5.665 1166.795 5.835 1166.965 ;
        RECT 6.125 1166.795 6.295 1166.965 ;
        RECT 6.585 1166.795 6.755 1166.965 ;
        RECT 2910.105 1166.795 2910.275 1166.965 ;
        RECT 2912.865 1166.795 2913.035 1166.965 ;
        RECT 2913.325 1166.795 2913.495 1166.965 ;
        RECT 2913.785 1166.795 2913.955 1166.965 ;
        RECT 5.665 1161.355 5.835 1161.525 ;
        RECT 6.125 1161.355 6.295 1161.525 ;
        RECT 6.585 1161.355 6.755 1161.525 ;
        RECT 2910.105 1161.355 2910.275 1161.525 ;
        RECT 2912.865 1161.355 2913.035 1161.525 ;
        RECT 2913.325 1161.355 2913.495 1161.525 ;
        RECT 2913.785 1161.355 2913.955 1161.525 ;
        RECT 5.665 1155.915 5.835 1156.085 ;
        RECT 6.125 1155.915 6.295 1156.085 ;
        RECT 6.585 1155.915 6.755 1156.085 ;
        RECT 2910.105 1155.915 2910.275 1156.085 ;
        RECT 2912.865 1155.915 2913.035 1156.085 ;
        RECT 2913.325 1155.915 2913.495 1156.085 ;
        RECT 2913.785 1155.915 2913.955 1156.085 ;
        RECT 5.665 1150.475 5.835 1150.645 ;
        RECT 6.125 1150.475 6.295 1150.645 ;
        RECT 6.585 1150.475 6.755 1150.645 ;
        RECT 2910.105 1150.475 2910.275 1150.645 ;
        RECT 2912.865 1150.475 2913.035 1150.645 ;
        RECT 2913.325 1150.475 2913.495 1150.645 ;
        RECT 2913.785 1150.475 2913.955 1150.645 ;
        RECT 5.665 1145.035 5.835 1145.205 ;
        RECT 6.125 1145.035 6.295 1145.205 ;
        RECT 6.585 1145.035 6.755 1145.205 ;
        RECT 2910.105 1145.035 2910.275 1145.205 ;
        RECT 2912.865 1145.035 2913.035 1145.205 ;
        RECT 2913.325 1145.035 2913.495 1145.205 ;
        RECT 2913.785 1145.035 2913.955 1145.205 ;
        RECT 5.665 1139.595 5.835 1139.765 ;
        RECT 6.125 1139.595 6.295 1139.765 ;
        RECT 6.585 1139.595 6.755 1139.765 ;
        RECT 2910.105 1139.595 2910.275 1139.765 ;
        RECT 2912.865 1139.595 2913.035 1139.765 ;
        RECT 2913.325 1139.595 2913.495 1139.765 ;
        RECT 2913.785 1139.595 2913.955 1139.765 ;
        RECT 5.665 1134.155 5.835 1134.325 ;
        RECT 6.125 1134.155 6.295 1134.325 ;
        RECT 6.585 1134.155 6.755 1134.325 ;
        RECT 2910.105 1134.155 2910.275 1134.325 ;
        RECT 2912.865 1134.155 2913.035 1134.325 ;
        RECT 2913.325 1134.155 2913.495 1134.325 ;
        RECT 2913.785 1134.155 2913.955 1134.325 ;
        RECT 5.665 1128.715 5.835 1128.885 ;
        RECT 6.125 1128.715 6.295 1128.885 ;
        RECT 6.585 1128.715 6.755 1128.885 ;
        RECT 2910.105 1128.715 2910.275 1128.885 ;
        RECT 2912.865 1128.715 2913.035 1128.885 ;
        RECT 2913.325 1128.715 2913.495 1128.885 ;
        RECT 2913.785 1128.715 2913.955 1128.885 ;
        RECT 5.665 1123.275 5.835 1123.445 ;
        RECT 6.125 1123.275 6.295 1123.445 ;
        RECT 6.585 1123.275 6.755 1123.445 ;
        RECT 2910.105 1123.275 2910.275 1123.445 ;
        RECT 2912.865 1123.275 2913.035 1123.445 ;
        RECT 2913.325 1123.275 2913.495 1123.445 ;
        RECT 2913.785 1123.275 2913.955 1123.445 ;
        RECT 5.665 1117.835 5.835 1118.005 ;
        RECT 6.125 1117.835 6.295 1118.005 ;
        RECT 6.585 1117.835 6.755 1118.005 ;
        RECT 2910.105 1117.835 2910.275 1118.005 ;
        RECT 2912.865 1117.835 2913.035 1118.005 ;
        RECT 2913.325 1117.835 2913.495 1118.005 ;
        RECT 2913.785 1117.835 2913.955 1118.005 ;
        RECT 5.665 1112.395 5.835 1112.565 ;
        RECT 6.125 1112.395 6.295 1112.565 ;
        RECT 6.585 1112.395 6.755 1112.565 ;
        RECT 8.885 1112.395 9.055 1112.565 ;
        RECT 9.345 1112.395 9.515 1112.565 ;
        RECT 9.805 1112.395 9.975 1112.565 ;
        RECT 2910.105 1112.395 2910.275 1112.565 ;
        RECT 2912.865 1112.395 2913.035 1112.565 ;
        RECT 2913.325 1112.395 2913.495 1112.565 ;
        RECT 2913.785 1112.395 2913.955 1112.565 ;
        RECT 5.665 1106.955 5.835 1107.125 ;
        RECT 6.125 1106.955 6.295 1107.125 ;
        RECT 6.585 1106.955 6.755 1107.125 ;
        RECT 2910.105 1106.955 2910.275 1107.125 ;
        RECT 2912.865 1106.955 2913.035 1107.125 ;
        RECT 2913.325 1106.955 2913.495 1107.125 ;
        RECT 2913.785 1106.955 2913.955 1107.125 ;
        RECT 5.665 1101.515 5.835 1101.685 ;
        RECT 6.125 1101.515 6.295 1101.685 ;
        RECT 6.585 1101.515 6.755 1101.685 ;
        RECT 2910.105 1101.515 2910.275 1101.685 ;
        RECT 2912.865 1101.515 2913.035 1101.685 ;
        RECT 2913.325 1101.515 2913.495 1101.685 ;
        RECT 2913.785 1101.515 2913.955 1101.685 ;
        RECT 5.665 1096.075 5.835 1096.245 ;
        RECT 6.125 1096.075 6.295 1096.245 ;
        RECT 6.585 1096.075 6.755 1096.245 ;
        RECT 2910.105 1096.075 2910.275 1096.245 ;
        RECT 2912.865 1096.075 2913.035 1096.245 ;
        RECT 2913.325 1096.075 2913.495 1096.245 ;
        RECT 2913.785 1096.075 2913.955 1096.245 ;
        RECT 5.665 1090.635 5.835 1090.805 ;
        RECT 6.125 1090.635 6.295 1090.805 ;
        RECT 6.585 1090.635 6.755 1090.805 ;
        RECT 2910.105 1090.635 2910.275 1090.805 ;
        RECT 2912.865 1090.635 2913.035 1090.805 ;
        RECT 2913.325 1090.635 2913.495 1090.805 ;
        RECT 2913.785 1090.635 2913.955 1090.805 ;
        RECT 5.665 1085.195 5.835 1085.365 ;
        RECT 6.125 1085.195 6.295 1085.365 ;
        RECT 6.585 1085.195 6.755 1085.365 ;
        RECT 2910.105 1085.195 2910.275 1085.365 ;
        RECT 2912.865 1085.195 2913.035 1085.365 ;
        RECT 2913.325 1085.195 2913.495 1085.365 ;
        RECT 2913.785 1085.195 2913.955 1085.365 ;
        RECT 5.665 1079.755 5.835 1079.925 ;
        RECT 6.125 1079.755 6.295 1079.925 ;
        RECT 6.585 1079.755 6.755 1079.925 ;
        RECT 2910.105 1079.755 2910.275 1079.925 ;
        RECT 2912.865 1079.755 2913.035 1079.925 ;
        RECT 2913.325 1079.755 2913.495 1079.925 ;
        RECT 2913.785 1079.755 2913.955 1079.925 ;
        RECT 5.665 1074.315 5.835 1074.485 ;
        RECT 6.125 1074.315 6.295 1074.485 ;
        RECT 6.585 1074.315 6.755 1074.485 ;
        RECT 2910.105 1074.315 2910.275 1074.485 ;
        RECT 2912.865 1074.315 2913.035 1074.485 ;
        RECT 2913.325 1074.315 2913.495 1074.485 ;
        RECT 2913.785 1074.315 2913.955 1074.485 ;
        RECT 5.665 1068.875 5.835 1069.045 ;
        RECT 6.125 1068.875 6.295 1069.045 ;
        RECT 6.585 1068.875 6.755 1069.045 ;
        RECT 2910.105 1068.875 2910.275 1069.045 ;
        RECT 2912.865 1068.875 2913.035 1069.045 ;
        RECT 2913.325 1068.875 2913.495 1069.045 ;
        RECT 2913.785 1068.875 2913.955 1069.045 ;
        RECT 5.665 1063.435 5.835 1063.605 ;
        RECT 6.125 1063.435 6.295 1063.605 ;
        RECT 6.585 1063.435 6.755 1063.605 ;
        RECT 2910.105 1063.435 2910.275 1063.605 ;
        RECT 2912.865 1063.435 2913.035 1063.605 ;
        RECT 2913.325 1063.435 2913.495 1063.605 ;
        RECT 2913.785 1063.435 2913.955 1063.605 ;
        RECT 5.665 1057.995 5.835 1058.165 ;
        RECT 6.125 1057.995 6.295 1058.165 ;
        RECT 6.585 1057.995 6.755 1058.165 ;
        RECT 2910.105 1057.995 2910.275 1058.165 ;
        RECT 2912.865 1057.995 2913.035 1058.165 ;
        RECT 2913.325 1057.995 2913.495 1058.165 ;
        RECT 2913.785 1057.995 2913.955 1058.165 ;
        RECT 5.665 1052.555 5.835 1052.725 ;
        RECT 6.125 1052.555 6.295 1052.725 ;
        RECT 6.585 1052.555 6.755 1052.725 ;
        RECT 2910.105 1052.555 2910.275 1052.725 ;
        RECT 2912.865 1052.555 2913.035 1052.725 ;
        RECT 2913.325 1052.555 2913.495 1052.725 ;
        RECT 2913.785 1052.555 2913.955 1052.725 ;
        RECT 5.665 1047.115 5.835 1047.285 ;
        RECT 6.125 1047.115 6.295 1047.285 ;
        RECT 6.585 1047.115 6.755 1047.285 ;
        RECT 2910.105 1047.115 2910.275 1047.285 ;
        RECT 2912.865 1047.115 2913.035 1047.285 ;
        RECT 2913.325 1047.115 2913.495 1047.285 ;
        RECT 2913.785 1047.115 2913.955 1047.285 ;
        RECT 5.665 1041.675 5.835 1041.845 ;
        RECT 6.125 1041.675 6.295 1041.845 ;
        RECT 6.585 1041.675 6.755 1041.845 ;
        RECT 2910.105 1041.675 2910.275 1041.845 ;
        RECT 2912.865 1041.675 2913.035 1041.845 ;
        RECT 2913.325 1041.675 2913.495 1041.845 ;
        RECT 2913.785 1041.675 2913.955 1041.845 ;
        RECT 5.665 1036.235 5.835 1036.405 ;
        RECT 6.125 1036.235 6.295 1036.405 ;
        RECT 6.585 1036.235 6.755 1036.405 ;
        RECT 8.885 1036.235 9.055 1036.405 ;
        RECT 9.345 1036.235 9.515 1036.405 ;
        RECT 9.805 1036.235 9.975 1036.405 ;
        RECT 2910.105 1036.235 2910.275 1036.405 ;
        RECT 2912.865 1036.235 2913.035 1036.405 ;
        RECT 2913.325 1036.235 2913.495 1036.405 ;
        RECT 2913.785 1036.235 2913.955 1036.405 ;
        RECT 5.665 1030.795 5.835 1030.965 ;
        RECT 6.125 1030.795 6.295 1030.965 ;
        RECT 6.585 1030.795 6.755 1030.965 ;
        RECT 2910.105 1030.795 2910.275 1030.965 ;
        RECT 2912.865 1030.795 2913.035 1030.965 ;
        RECT 2913.325 1030.795 2913.495 1030.965 ;
        RECT 2913.785 1030.795 2913.955 1030.965 ;
        RECT 5.665 1025.355 5.835 1025.525 ;
        RECT 6.125 1025.355 6.295 1025.525 ;
        RECT 6.585 1025.355 6.755 1025.525 ;
        RECT 2910.105 1025.355 2910.275 1025.525 ;
        RECT 2912.865 1025.355 2913.035 1025.525 ;
        RECT 2913.325 1025.355 2913.495 1025.525 ;
        RECT 2913.785 1025.355 2913.955 1025.525 ;
        RECT 5.665 1019.915 5.835 1020.085 ;
        RECT 6.125 1019.915 6.295 1020.085 ;
        RECT 6.585 1019.915 6.755 1020.085 ;
        RECT 2910.105 1019.915 2910.275 1020.085 ;
        RECT 2912.865 1019.915 2913.035 1020.085 ;
        RECT 2913.325 1019.915 2913.495 1020.085 ;
        RECT 2913.785 1019.915 2913.955 1020.085 ;
        RECT 5.665 1014.475 5.835 1014.645 ;
        RECT 6.125 1014.475 6.295 1014.645 ;
        RECT 6.585 1014.475 6.755 1014.645 ;
        RECT 2910.105 1014.475 2910.275 1014.645 ;
        RECT 2912.865 1014.475 2913.035 1014.645 ;
        RECT 2913.325 1014.475 2913.495 1014.645 ;
        RECT 2913.785 1014.475 2913.955 1014.645 ;
        RECT 5.665 1009.035 5.835 1009.205 ;
        RECT 6.125 1009.035 6.295 1009.205 ;
        RECT 6.585 1009.035 6.755 1009.205 ;
        RECT 2909.185 1009.035 2909.355 1009.205 ;
        RECT 2909.645 1009.035 2909.815 1009.205 ;
        RECT 2910.105 1009.035 2910.275 1009.205 ;
        RECT 2912.865 1009.035 2913.035 1009.205 ;
        RECT 2913.325 1009.035 2913.495 1009.205 ;
        RECT 2913.785 1009.035 2913.955 1009.205 ;
        RECT 5.665 1003.595 5.835 1003.765 ;
        RECT 6.125 1003.595 6.295 1003.765 ;
        RECT 6.585 1003.595 6.755 1003.765 ;
        RECT 2910.105 1003.595 2910.275 1003.765 ;
        RECT 2912.865 1003.595 2913.035 1003.765 ;
        RECT 2913.325 1003.595 2913.495 1003.765 ;
        RECT 2913.785 1003.595 2913.955 1003.765 ;
        RECT 5.665 998.155 5.835 998.325 ;
        RECT 6.125 998.155 6.295 998.325 ;
        RECT 6.585 998.155 6.755 998.325 ;
        RECT 2909.185 998.155 2909.355 998.325 ;
        RECT 2909.645 998.155 2909.815 998.325 ;
        RECT 2910.105 998.155 2910.275 998.325 ;
        RECT 2912.865 998.155 2913.035 998.325 ;
        RECT 2913.325 998.155 2913.495 998.325 ;
        RECT 2913.785 998.155 2913.955 998.325 ;
        RECT 5.665 992.715 5.835 992.885 ;
        RECT 6.125 992.715 6.295 992.885 ;
        RECT 6.585 992.715 6.755 992.885 ;
        RECT 2910.105 992.715 2910.275 992.885 ;
        RECT 2912.865 992.715 2913.035 992.885 ;
        RECT 2913.325 992.715 2913.495 992.885 ;
        RECT 2913.785 992.715 2913.955 992.885 ;
        RECT 5.665 987.275 5.835 987.445 ;
        RECT 6.125 987.275 6.295 987.445 ;
        RECT 6.585 987.275 6.755 987.445 ;
        RECT 2910.105 987.275 2910.275 987.445 ;
        RECT 2912.865 987.275 2913.035 987.445 ;
        RECT 2913.325 987.275 2913.495 987.445 ;
        RECT 2913.785 987.275 2913.955 987.445 ;
        RECT 5.665 981.835 5.835 982.005 ;
        RECT 6.125 981.835 6.295 982.005 ;
        RECT 6.585 981.835 6.755 982.005 ;
        RECT 2910.105 981.835 2910.275 982.005 ;
        RECT 2912.865 981.835 2913.035 982.005 ;
        RECT 2913.325 981.835 2913.495 982.005 ;
        RECT 2913.785 981.835 2913.955 982.005 ;
        RECT 5.665 976.395 5.835 976.565 ;
        RECT 6.125 976.395 6.295 976.565 ;
        RECT 6.585 976.395 6.755 976.565 ;
        RECT 2910.105 976.395 2910.275 976.565 ;
        RECT 2912.865 976.395 2913.035 976.565 ;
        RECT 2913.325 976.395 2913.495 976.565 ;
        RECT 2913.785 976.395 2913.955 976.565 ;
        RECT 5.665 970.955 5.835 971.125 ;
        RECT 6.125 970.955 6.295 971.125 ;
        RECT 6.585 970.955 6.755 971.125 ;
        RECT 2910.105 970.955 2910.275 971.125 ;
        RECT 2912.865 970.955 2913.035 971.125 ;
        RECT 2913.325 970.955 2913.495 971.125 ;
        RECT 2913.785 970.955 2913.955 971.125 ;
        RECT 5.665 965.515 5.835 965.685 ;
        RECT 6.125 965.515 6.295 965.685 ;
        RECT 6.585 965.515 6.755 965.685 ;
        RECT 2910.105 965.515 2910.275 965.685 ;
        RECT 2912.865 965.515 2913.035 965.685 ;
        RECT 2913.325 965.515 2913.495 965.685 ;
        RECT 2913.785 965.515 2913.955 965.685 ;
        RECT 5.665 960.075 5.835 960.245 ;
        RECT 6.125 960.075 6.295 960.245 ;
        RECT 6.585 960.075 6.755 960.245 ;
        RECT 2910.105 960.075 2910.275 960.245 ;
        RECT 2912.865 960.075 2913.035 960.245 ;
        RECT 2913.325 960.075 2913.495 960.245 ;
        RECT 2913.785 960.075 2913.955 960.245 ;
        RECT 5.665 954.635 5.835 954.805 ;
        RECT 6.125 954.635 6.295 954.805 ;
        RECT 6.585 954.635 6.755 954.805 ;
        RECT 2910.105 954.635 2910.275 954.805 ;
        RECT 2912.865 954.635 2913.035 954.805 ;
        RECT 2913.325 954.635 2913.495 954.805 ;
        RECT 2913.785 954.635 2913.955 954.805 ;
        RECT 5.665 949.195 5.835 949.365 ;
        RECT 6.125 949.195 6.295 949.365 ;
        RECT 6.585 949.195 6.755 949.365 ;
        RECT 2910.105 949.195 2910.275 949.365 ;
        RECT 2912.865 949.195 2913.035 949.365 ;
        RECT 2913.325 949.195 2913.495 949.365 ;
        RECT 2913.785 949.195 2913.955 949.365 ;
        RECT 5.665 943.755 5.835 943.925 ;
        RECT 6.125 943.755 6.295 943.925 ;
        RECT 6.585 943.755 6.755 943.925 ;
        RECT 2910.105 943.755 2910.275 943.925 ;
        RECT 2912.865 943.755 2913.035 943.925 ;
        RECT 2913.325 943.755 2913.495 943.925 ;
        RECT 2913.785 943.755 2913.955 943.925 ;
        RECT 5.665 938.315 5.835 938.485 ;
        RECT 6.125 938.315 6.295 938.485 ;
        RECT 6.585 938.315 6.755 938.485 ;
        RECT 2910.105 938.315 2910.275 938.485 ;
        RECT 2912.865 938.315 2913.035 938.485 ;
        RECT 2913.325 938.315 2913.495 938.485 ;
        RECT 2913.785 938.315 2913.955 938.485 ;
        RECT 5.665 932.875 5.835 933.045 ;
        RECT 6.125 932.875 6.295 933.045 ;
        RECT 6.585 932.875 6.755 933.045 ;
        RECT 2910.105 932.875 2910.275 933.045 ;
        RECT 2912.865 932.875 2913.035 933.045 ;
        RECT 2913.325 932.875 2913.495 933.045 ;
        RECT 2913.785 932.875 2913.955 933.045 ;
        RECT 5.665 927.435 5.835 927.605 ;
        RECT 6.125 927.435 6.295 927.605 ;
        RECT 6.585 927.435 6.755 927.605 ;
        RECT 2910.105 927.435 2910.275 927.605 ;
        RECT 2912.865 927.435 2913.035 927.605 ;
        RECT 2913.325 927.435 2913.495 927.605 ;
        RECT 2913.785 927.435 2913.955 927.605 ;
        RECT 5.665 921.995 5.835 922.165 ;
        RECT 6.125 921.995 6.295 922.165 ;
        RECT 6.585 921.995 6.755 922.165 ;
        RECT 2910.105 921.995 2910.275 922.165 ;
        RECT 2912.865 921.995 2913.035 922.165 ;
        RECT 2913.325 921.995 2913.495 922.165 ;
        RECT 2913.785 921.995 2913.955 922.165 ;
        RECT 5.665 916.555 5.835 916.725 ;
        RECT 6.125 916.555 6.295 916.725 ;
        RECT 6.585 916.555 6.755 916.725 ;
        RECT 2910.105 916.555 2910.275 916.725 ;
        RECT 2912.865 916.555 2913.035 916.725 ;
        RECT 2913.325 916.555 2913.495 916.725 ;
        RECT 2913.785 916.555 2913.955 916.725 ;
        RECT 5.665 911.115 5.835 911.285 ;
        RECT 6.125 911.115 6.295 911.285 ;
        RECT 6.585 911.115 6.755 911.285 ;
        RECT 2910.105 911.115 2910.275 911.285 ;
        RECT 2912.865 911.115 2913.035 911.285 ;
        RECT 2913.325 911.115 2913.495 911.285 ;
        RECT 2913.785 911.115 2913.955 911.285 ;
        RECT 5.665 905.675 5.835 905.845 ;
        RECT 6.125 905.675 6.295 905.845 ;
        RECT 6.585 905.675 6.755 905.845 ;
        RECT 2910.105 905.675 2910.275 905.845 ;
        RECT 2912.865 905.675 2913.035 905.845 ;
        RECT 2913.325 905.675 2913.495 905.845 ;
        RECT 2913.785 905.675 2913.955 905.845 ;
        RECT 5.665 900.235 5.835 900.405 ;
        RECT 6.125 900.235 6.295 900.405 ;
        RECT 6.585 900.235 6.755 900.405 ;
        RECT 2910.105 900.235 2910.275 900.405 ;
        RECT 2912.865 900.235 2913.035 900.405 ;
        RECT 2913.325 900.235 2913.495 900.405 ;
        RECT 2913.785 900.235 2913.955 900.405 ;
        RECT 5.665 894.795 5.835 894.965 ;
        RECT 6.125 894.795 6.295 894.965 ;
        RECT 6.585 894.795 6.755 894.965 ;
        RECT 2910.105 894.795 2910.275 894.965 ;
        RECT 2912.865 894.795 2913.035 894.965 ;
        RECT 2913.325 894.795 2913.495 894.965 ;
        RECT 2913.785 894.795 2913.955 894.965 ;
        RECT 5.665 889.355 5.835 889.525 ;
        RECT 6.125 889.355 6.295 889.525 ;
        RECT 6.585 889.355 6.755 889.525 ;
        RECT 2910.105 889.355 2910.275 889.525 ;
        RECT 2912.865 889.355 2913.035 889.525 ;
        RECT 2913.325 889.355 2913.495 889.525 ;
        RECT 2913.785 889.355 2913.955 889.525 ;
        RECT 5.665 883.915 5.835 884.085 ;
        RECT 6.125 883.915 6.295 884.085 ;
        RECT 6.585 883.915 6.755 884.085 ;
        RECT 2910.105 883.915 2910.275 884.085 ;
        RECT 2912.865 883.915 2913.035 884.085 ;
        RECT 2913.325 883.915 2913.495 884.085 ;
        RECT 2913.785 883.915 2913.955 884.085 ;
        RECT 5.665 878.475 5.835 878.645 ;
        RECT 6.125 878.475 6.295 878.645 ;
        RECT 6.585 878.475 6.755 878.645 ;
        RECT 2910.105 878.475 2910.275 878.645 ;
        RECT 2912.865 878.475 2913.035 878.645 ;
        RECT 2913.325 878.475 2913.495 878.645 ;
        RECT 2913.785 878.475 2913.955 878.645 ;
        RECT 5.665 873.035 5.835 873.205 ;
        RECT 6.125 873.035 6.295 873.205 ;
        RECT 6.585 873.035 6.755 873.205 ;
        RECT 2910.105 873.035 2910.275 873.205 ;
        RECT 2912.865 873.035 2913.035 873.205 ;
        RECT 2913.325 873.035 2913.495 873.205 ;
        RECT 2913.785 873.035 2913.955 873.205 ;
        RECT 5.665 867.595 5.835 867.765 ;
        RECT 6.125 867.595 6.295 867.765 ;
        RECT 6.585 867.595 6.755 867.765 ;
        RECT 2910.105 867.595 2910.275 867.765 ;
        RECT 2912.865 867.595 2913.035 867.765 ;
        RECT 2913.325 867.595 2913.495 867.765 ;
        RECT 2913.785 867.595 2913.955 867.765 ;
        RECT 5.665 862.155 5.835 862.325 ;
        RECT 6.125 862.155 6.295 862.325 ;
        RECT 6.585 862.155 6.755 862.325 ;
        RECT 2910.105 862.155 2910.275 862.325 ;
        RECT 2912.865 862.155 2913.035 862.325 ;
        RECT 2913.325 862.155 2913.495 862.325 ;
        RECT 2913.785 862.155 2913.955 862.325 ;
        RECT 5.665 856.715 5.835 856.885 ;
        RECT 6.125 856.715 6.295 856.885 ;
        RECT 6.585 856.715 6.755 856.885 ;
        RECT 2910.105 856.715 2910.275 856.885 ;
        RECT 2912.865 856.715 2913.035 856.885 ;
        RECT 2913.325 856.715 2913.495 856.885 ;
        RECT 2913.785 856.715 2913.955 856.885 ;
        RECT 5.665 851.275 5.835 851.445 ;
        RECT 6.125 851.275 6.295 851.445 ;
        RECT 6.585 851.275 6.755 851.445 ;
        RECT 2910.105 851.275 2910.275 851.445 ;
        RECT 2912.865 851.275 2913.035 851.445 ;
        RECT 2913.325 851.275 2913.495 851.445 ;
        RECT 2913.785 851.275 2913.955 851.445 ;
        RECT 5.665 845.835 5.835 846.005 ;
        RECT 6.125 845.835 6.295 846.005 ;
        RECT 6.585 845.835 6.755 846.005 ;
        RECT 2910.105 845.835 2910.275 846.005 ;
        RECT 2912.865 845.835 2913.035 846.005 ;
        RECT 2913.325 845.835 2913.495 846.005 ;
        RECT 2913.785 845.835 2913.955 846.005 ;
        RECT 5.665 840.395 5.835 840.565 ;
        RECT 6.125 840.395 6.295 840.565 ;
        RECT 6.585 840.395 6.755 840.565 ;
        RECT 2910.105 840.395 2910.275 840.565 ;
        RECT 2912.865 840.395 2913.035 840.565 ;
        RECT 2913.325 840.395 2913.495 840.565 ;
        RECT 2913.785 840.395 2913.955 840.565 ;
        RECT 5.665 834.955 5.835 835.125 ;
        RECT 6.125 834.955 6.295 835.125 ;
        RECT 6.585 834.955 6.755 835.125 ;
        RECT 2910.105 834.955 2910.275 835.125 ;
        RECT 2912.865 834.955 2913.035 835.125 ;
        RECT 2913.325 834.955 2913.495 835.125 ;
        RECT 2913.785 834.955 2913.955 835.125 ;
        RECT 5.665 829.515 5.835 829.685 ;
        RECT 6.125 829.515 6.295 829.685 ;
        RECT 6.585 829.515 6.755 829.685 ;
        RECT 2910.105 829.515 2910.275 829.685 ;
        RECT 2912.865 829.515 2913.035 829.685 ;
        RECT 2913.325 829.515 2913.495 829.685 ;
        RECT 2913.785 829.515 2913.955 829.685 ;
        RECT 5.665 824.075 5.835 824.245 ;
        RECT 6.125 824.075 6.295 824.245 ;
        RECT 6.585 824.075 6.755 824.245 ;
        RECT 2910.105 824.075 2910.275 824.245 ;
        RECT 2912.865 824.075 2913.035 824.245 ;
        RECT 2913.325 824.075 2913.495 824.245 ;
        RECT 2913.785 824.075 2913.955 824.245 ;
        RECT 5.665 818.635 5.835 818.805 ;
        RECT 6.125 818.635 6.295 818.805 ;
        RECT 6.585 818.635 6.755 818.805 ;
        RECT 2910.105 818.635 2910.275 818.805 ;
        RECT 2912.865 818.635 2913.035 818.805 ;
        RECT 2913.325 818.635 2913.495 818.805 ;
        RECT 2913.785 818.635 2913.955 818.805 ;
        RECT 5.665 813.195 5.835 813.365 ;
        RECT 6.125 813.195 6.295 813.365 ;
        RECT 6.585 813.195 6.755 813.365 ;
        RECT 2909.185 813.195 2909.355 813.365 ;
        RECT 2909.645 813.195 2909.815 813.365 ;
        RECT 2910.105 813.195 2910.275 813.365 ;
        RECT 2912.865 813.195 2913.035 813.365 ;
        RECT 2913.325 813.195 2913.495 813.365 ;
        RECT 2913.785 813.195 2913.955 813.365 ;
        RECT 5.665 807.755 5.835 807.925 ;
        RECT 6.125 807.755 6.295 807.925 ;
        RECT 6.585 807.755 6.755 807.925 ;
        RECT 2910.105 807.755 2910.275 807.925 ;
        RECT 2912.865 807.755 2913.035 807.925 ;
        RECT 2913.325 807.755 2913.495 807.925 ;
        RECT 2913.785 807.755 2913.955 807.925 ;
        RECT 5.665 802.315 5.835 802.485 ;
        RECT 6.125 802.315 6.295 802.485 ;
        RECT 6.585 802.315 6.755 802.485 ;
        RECT 2910.105 802.315 2910.275 802.485 ;
        RECT 2912.865 802.315 2913.035 802.485 ;
        RECT 2913.325 802.315 2913.495 802.485 ;
        RECT 2913.785 802.315 2913.955 802.485 ;
        RECT 5.665 796.875 5.835 797.045 ;
        RECT 6.125 796.875 6.295 797.045 ;
        RECT 6.585 796.875 6.755 797.045 ;
        RECT 2910.105 796.875 2910.275 797.045 ;
        RECT 2912.865 796.875 2913.035 797.045 ;
        RECT 2913.325 796.875 2913.495 797.045 ;
        RECT 2913.785 796.875 2913.955 797.045 ;
        RECT 5.665 791.435 5.835 791.605 ;
        RECT 6.125 791.435 6.295 791.605 ;
        RECT 6.585 791.435 6.755 791.605 ;
        RECT 2910.105 791.435 2910.275 791.605 ;
        RECT 2912.865 791.435 2913.035 791.605 ;
        RECT 2913.325 791.435 2913.495 791.605 ;
        RECT 2913.785 791.435 2913.955 791.605 ;
        RECT 5.665 785.995 5.835 786.165 ;
        RECT 6.125 785.995 6.295 786.165 ;
        RECT 6.585 785.995 6.755 786.165 ;
        RECT 2910.105 785.995 2910.275 786.165 ;
        RECT 2912.865 785.995 2913.035 786.165 ;
        RECT 2913.325 785.995 2913.495 786.165 ;
        RECT 2913.785 785.995 2913.955 786.165 ;
        RECT 5.665 780.555 5.835 780.725 ;
        RECT 6.125 780.555 6.295 780.725 ;
        RECT 6.585 780.555 6.755 780.725 ;
        RECT 2910.105 780.555 2910.275 780.725 ;
        RECT 2912.865 780.555 2913.035 780.725 ;
        RECT 2913.325 780.555 2913.495 780.725 ;
        RECT 2913.785 780.555 2913.955 780.725 ;
        RECT 5.665 775.115 5.835 775.285 ;
        RECT 6.125 775.115 6.295 775.285 ;
        RECT 6.585 775.115 6.755 775.285 ;
        RECT 2910.105 775.115 2910.275 775.285 ;
        RECT 2912.865 775.115 2913.035 775.285 ;
        RECT 2913.325 775.115 2913.495 775.285 ;
        RECT 2913.785 775.115 2913.955 775.285 ;
        RECT 5.665 769.675 5.835 769.845 ;
        RECT 6.125 769.675 6.295 769.845 ;
        RECT 6.585 769.675 6.755 769.845 ;
        RECT 2910.105 769.675 2910.275 769.845 ;
        RECT 2912.865 769.675 2913.035 769.845 ;
        RECT 2913.325 769.675 2913.495 769.845 ;
        RECT 2913.785 769.675 2913.955 769.845 ;
        RECT 5.665 764.235 5.835 764.405 ;
        RECT 6.125 764.235 6.295 764.405 ;
        RECT 6.585 764.235 6.755 764.405 ;
        RECT 2910.105 764.235 2910.275 764.405 ;
        RECT 2912.865 764.235 2913.035 764.405 ;
        RECT 2913.325 764.235 2913.495 764.405 ;
        RECT 2913.785 764.235 2913.955 764.405 ;
        RECT 5.665 758.795 5.835 758.965 ;
        RECT 6.125 758.795 6.295 758.965 ;
        RECT 6.585 758.795 6.755 758.965 ;
        RECT 2910.105 758.795 2910.275 758.965 ;
        RECT 2912.865 758.795 2913.035 758.965 ;
        RECT 2913.325 758.795 2913.495 758.965 ;
        RECT 2913.785 758.795 2913.955 758.965 ;
        RECT 5.665 753.355 5.835 753.525 ;
        RECT 6.125 753.355 6.295 753.525 ;
        RECT 6.585 753.355 6.755 753.525 ;
        RECT 2910.105 753.355 2910.275 753.525 ;
        RECT 2912.865 753.355 2913.035 753.525 ;
        RECT 2913.325 753.355 2913.495 753.525 ;
        RECT 2913.785 753.355 2913.955 753.525 ;
        RECT 5.665 747.915 5.835 748.085 ;
        RECT 6.125 747.915 6.295 748.085 ;
        RECT 6.585 747.915 6.755 748.085 ;
        RECT 2910.105 747.915 2910.275 748.085 ;
        RECT 2912.865 747.915 2913.035 748.085 ;
        RECT 2913.325 747.915 2913.495 748.085 ;
        RECT 2913.785 747.915 2913.955 748.085 ;
        RECT 5.665 742.475 5.835 742.645 ;
        RECT 6.125 742.475 6.295 742.645 ;
        RECT 6.585 742.475 6.755 742.645 ;
        RECT 2910.105 742.475 2910.275 742.645 ;
        RECT 2912.865 742.475 2913.035 742.645 ;
        RECT 2913.325 742.475 2913.495 742.645 ;
        RECT 2913.785 742.475 2913.955 742.645 ;
        RECT 5.665 737.035 5.835 737.205 ;
        RECT 6.125 737.035 6.295 737.205 ;
        RECT 6.585 737.035 6.755 737.205 ;
        RECT 2909.185 737.035 2909.355 737.205 ;
        RECT 2909.645 737.035 2909.815 737.205 ;
        RECT 2910.105 737.035 2910.275 737.205 ;
        RECT 2912.865 737.035 2913.035 737.205 ;
        RECT 2913.325 737.035 2913.495 737.205 ;
        RECT 2913.785 737.035 2913.955 737.205 ;
        RECT 5.665 731.595 5.835 731.765 ;
        RECT 6.125 731.595 6.295 731.765 ;
        RECT 6.585 731.595 6.755 731.765 ;
        RECT 2910.105 731.595 2910.275 731.765 ;
        RECT 2912.865 731.595 2913.035 731.765 ;
        RECT 2913.325 731.595 2913.495 731.765 ;
        RECT 2913.785 731.595 2913.955 731.765 ;
        RECT 5.665 726.155 5.835 726.325 ;
        RECT 6.125 726.155 6.295 726.325 ;
        RECT 6.585 726.155 6.755 726.325 ;
        RECT 2910.105 726.155 2910.275 726.325 ;
        RECT 2912.865 726.155 2913.035 726.325 ;
        RECT 2913.325 726.155 2913.495 726.325 ;
        RECT 2913.785 726.155 2913.955 726.325 ;
        RECT 5.665 720.715 5.835 720.885 ;
        RECT 6.125 720.715 6.295 720.885 ;
        RECT 6.585 720.715 6.755 720.885 ;
        RECT 8.885 720.715 9.055 720.885 ;
        RECT 9.345 720.715 9.515 720.885 ;
        RECT 9.805 720.715 9.975 720.885 ;
        RECT 2910.105 720.715 2910.275 720.885 ;
        RECT 2912.865 720.715 2913.035 720.885 ;
        RECT 2913.325 720.715 2913.495 720.885 ;
        RECT 2913.785 720.715 2913.955 720.885 ;
        RECT 5.665 715.275 5.835 715.445 ;
        RECT 6.125 715.275 6.295 715.445 ;
        RECT 6.585 715.275 6.755 715.445 ;
        RECT 2910.105 715.275 2910.275 715.445 ;
        RECT 2912.865 715.275 2913.035 715.445 ;
        RECT 2913.325 715.275 2913.495 715.445 ;
        RECT 2913.785 715.275 2913.955 715.445 ;
        RECT 5.665 709.835 5.835 710.005 ;
        RECT 6.125 709.835 6.295 710.005 ;
        RECT 6.585 709.835 6.755 710.005 ;
        RECT 2910.105 709.835 2910.275 710.005 ;
        RECT 2912.865 709.835 2913.035 710.005 ;
        RECT 2913.325 709.835 2913.495 710.005 ;
        RECT 2913.785 709.835 2913.955 710.005 ;
        RECT 5.665 704.395 5.835 704.565 ;
        RECT 6.125 704.395 6.295 704.565 ;
        RECT 6.585 704.395 6.755 704.565 ;
        RECT 2910.105 704.395 2910.275 704.565 ;
        RECT 2912.865 704.395 2913.035 704.565 ;
        RECT 2913.325 704.395 2913.495 704.565 ;
        RECT 2913.785 704.395 2913.955 704.565 ;
        RECT 5.665 698.955 5.835 699.125 ;
        RECT 6.125 698.955 6.295 699.125 ;
        RECT 6.585 698.955 6.755 699.125 ;
        RECT 2910.105 698.955 2910.275 699.125 ;
        RECT 2912.865 698.955 2913.035 699.125 ;
        RECT 2913.325 698.955 2913.495 699.125 ;
        RECT 2913.785 698.955 2913.955 699.125 ;
        RECT 5.665 693.515 5.835 693.685 ;
        RECT 6.125 693.515 6.295 693.685 ;
        RECT 6.585 693.515 6.755 693.685 ;
        RECT 2910.105 693.515 2910.275 693.685 ;
        RECT 2912.865 693.515 2913.035 693.685 ;
        RECT 2913.325 693.515 2913.495 693.685 ;
        RECT 2913.785 693.515 2913.955 693.685 ;
        RECT 5.665 688.075 5.835 688.245 ;
        RECT 6.125 688.075 6.295 688.245 ;
        RECT 6.585 688.075 6.755 688.245 ;
        RECT 2910.105 688.075 2910.275 688.245 ;
        RECT 2912.865 688.075 2913.035 688.245 ;
        RECT 2913.325 688.075 2913.495 688.245 ;
        RECT 2913.785 688.075 2913.955 688.245 ;
        RECT 5.665 682.635 5.835 682.805 ;
        RECT 6.125 682.635 6.295 682.805 ;
        RECT 6.585 682.635 6.755 682.805 ;
        RECT 2910.105 682.635 2910.275 682.805 ;
        RECT 2912.865 682.635 2913.035 682.805 ;
        RECT 2913.325 682.635 2913.495 682.805 ;
        RECT 2913.785 682.635 2913.955 682.805 ;
        RECT 5.665 677.195 5.835 677.365 ;
        RECT 6.125 677.195 6.295 677.365 ;
        RECT 6.585 677.195 6.755 677.365 ;
        RECT 2910.105 677.195 2910.275 677.365 ;
        RECT 2912.865 677.195 2913.035 677.365 ;
        RECT 2913.325 677.195 2913.495 677.365 ;
        RECT 2913.785 677.195 2913.955 677.365 ;
        RECT 5.665 671.755 5.835 671.925 ;
        RECT 6.125 671.755 6.295 671.925 ;
        RECT 6.585 671.755 6.755 671.925 ;
        RECT 2910.105 671.755 2910.275 671.925 ;
        RECT 2912.865 671.755 2913.035 671.925 ;
        RECT 2913.325 671.755 2913.495 671.925 ;
        RECT 2913.785 671.755 2913.955 671.925 ;
        RECT 5.665 666.315 5.835 666.485 ;
        RECT 6.125 666.315 6.295 666.485 ;
        RECT 6.585 666.315 6.755 666.485 ;
        RECT 2910.105 666.315 2910.275 666.485 ;
        RECT 2912.865 666.315 2913.035 666.485 ;
        RECT 2913.325 666.315 2913.495 666.485 ;
        RECT 2913.785 666.315 2913.955 666.485 ;
        RECT 5.665 660.875 5.835 661.045 ;
        RECT 6.125 660.875 6.295 661.045 ;
        RECT 6.585 660.875 6.755 661.045 ;
        RECT 2910.105 660.875 2910.275 661.045 ;
        RECT 2912.865 660.875 2913.035 661.045 ;
        RECT 2913.325 660.875 2913.495 661.045 ;
        RECT 2913.785 660.875 2913.955 661.045 ;
        RECT 5.665 655.435 5.835 655.605 ;
        RECT 6.125 655.435 6.295 655.605 ;
        RECT 6.585 655.435 6.755 655.605 ;
        RECT 2910.105 655.435 2910.275 655.605 ;
        RECT 2912.865 655.435 2913.035 655.605 ;
        RECT 2913.325 655.435 2913.495 655.605 ;
        RECT 2913.785 655.435 2913.955 655.605 ;
        RECT 5.665 649.995 5.835 650.165 ;
        RECT 6.125 649.995 6.295 650.165 ;
        RECT 6.585 649.995 6.755 650.165 ;
        RECT 2910.105 649.995 2910.275 650.165 ;
        RECT 2912.865 649.995 2913.035 650.165 ;
        RECT 2913.325 649.995 2913.495 650.165 ;
        RECT 2913.785 649.995 2913.955 650.165 ;
        RECT 5.665 644.555 5.835 644.725 ;
        RECT 6.125 644.555 6.295 644.725 ;
        RECT 6.585 644.555 6.755 644.725 ;
        RECT 2910.105 644.555 2910.275 644.725 ;
        RECT 2912.865 644.555 2913.035 644.725 ;
        RECT 2913.325 644.555 2913.495 644.725 ;
        RECT 2913.785 644.555 2913.955 644.725 ;
        RECT 5.665 639.115 5.835 639.285 ;
        RECT 6.125 639.115 6.295 639.285 ;
        RECT 6.585 639.115 6.755 639.285 ;
        RECT 2910.105 639.115 2910.275 639.285 ;
        RECT 2912.865 639.115 2913.035 639.285 ;
        RECT 2913.325 639.115 2913.495 639.285 ;
        RECT 2913.785 639.115 2913.955 639.285 ;
        RECT 5.665 633.675 5.835 633.845 ;
        RECT 6.125 633.675 6.295 633.845 ;
        RECT 6.585 633.675 6.755 633.845 ;
        RECT 2910.105 633.675 2910.275 633.845 ;
        RECT 2912.865 633.675 2913.035 633.845 ;
        RECT 2913.325 633.675 2913.495 633.845 ;
        RECT 2913.785 633.675 2913.955 633.845 ;
        RECT 5.665 628.235 5.835 628.405 ;
        RECT 6.125 628.235 6.295 628.405 ;
        RECT 6.585 628.235 6.755 628.405 ;
        RECT 8.885 628.235 9.055 628.405 ;
        RECT 9.345 628.235 9.515 628.405 ;
        RECT 9.805 628.235 9.975 628.405 ;
        RECT 2910.105 628.235 2910.275 628.405 ;
        RECT 2912.865 628.235 2913.035 628.405 ;
        RECT 2913.325 628.235 2913.495 628.405 ;
        RECT 2913.785 628.235 2913.955 628.405 ;
        RECT 5.665 622.795 5.835 622.965 ;
        RECT 6.125 622.795 6.295 622.965 ;
        RECT 6.585 622.795 6.755 622.965 ;
        RECT 2910.105 622.795 2910.275 622.965 ;
        RECT 2912.865 622.795 2913.035 622.965 ;
        RECT 2913.325 622.795 2913.495 622.965 ;
        RECT 2913.785 622.795 2913.955 622.965 ;
        RECT 5.665 617.355 5.835 617.525 ;
        RECT 6.125 617.355 6.295 617.525 ;
        RECT 6.585 617.355 6.755 617.525 ;
        RECT 2910.105 617.355 2910.275 617.525 ;
        RECT 2912.865 617.355 2913.035 617.525 ;
        RECT 2913.325 617.355 2913.495 617.525 ;
        RECT 2913.785 617.355 2913.955 617.525 ;
        RECT 5.665 611.915 5.835 612.085 ;
        RECT 6.125 611.915 6.295 612.085 ;
        RECT 6.585 611.915 6.755 612.085 ;
        RECT 2910.105 611.915 2910.275 612.085 ;
        RECT 2912.865 611.915 2913.035 612.085 ;
        RECT 2913.325 611.915 2913.495 612.085 ;
        RECT 2913.785 611.915 2913.955 612.085 ;
        RECT 5.665 606.475 5.835 606.645 ;
        RECT 6.125 606.475 6.295 606.645 ;
        RECT 6.585 606.475 6.755 606.645 ;
        RECT 2910.105 606.475 2910.275 606.645 ;
        RECT 2912.865 606.475 2913.035 606.645 ;
        RECT 2913.325 606.475 2913.495 606.645 ;
        RECT 2913.785 606.475 2913.955 606.645 ;
        RECT 5.665 601.035 5.835 601.205 ;
        RECT 6.125 601.035 6.295 601.205 ;
        RECT 6.585 601.035 6.755 601.205 ;
        RECT 8.885 601.035 9.055 601.205 ;
        RECT 9.345 601.035 9.515 601.205 ;
        RECT 9.805 601.035 9.975 601.205 ;
        RECT 2910.105 601.035 2910.275 601.205 ;
        RECT 2912.865 601.035 2913.035 601.205 ;
        RECT 2913.325 601.035 2913.495 601.205 ;
        RECT 2913.785 601.035 2913.955 601.205 ;
        RECT 5.665 595.595 5.835 595.765 ;
        RECT 6.125 595.595 6.295 595.765 ;
        RECT 6.585 595.595 6.755 595.765 ;
        RECT 2910.105 595.595 2910.275 595.765 ;
        RECT 2912.865 595.595 2913.035 595.765 ;
        RECT 2913.325 595.595 2913.495 595.765 ;
        RECT 2913.785 595.595 2913.955 595.765 ;
        RECT 5.665 590.155 5.835 590.325 ;
        RECT 6.125 590.155 6.295 590.325 ;
        RECT 6.585 590.155 6.755 590.325 ;
        RECT 2910.105 590.155 2910.275 590.325 ;
        RECT 2912.865 590.155 2913.035 590.325 ;
        RECT 2913.325 590.155 2913.495 590.325 ;
        RECT 2913.785 590.155 2913.955 590.325 ;
        RECT 5.665 584.715 5.835 584.885 ;
        RECT 6.125 584.715 6.295 584.885 ;
        RECT 6.585 584.715 6.755 584.885 ;
        RECT 2910.105 584.715 2910.275 584.885 ;
        RECT 2912.865 584.715 2913.035 584.885 ;
        RECT 2913.325 584.715 2913.495 584.885 ;
        RECT 2913.785 584.715 2913.955 584.885 ;
        RECT 5.665 579.275 5.835 579.445 ;
        RECT 6.125 579.275 6.295 579.445 ;
        RECT 6.585 579.275 6.755 579.445 ;
        RECT 2910.105 579.275 2910.275 579.445 ;
        RECT 2912.865 579.275 2913.035 579.445 ;
        RECT 2913.325 579.275 2913.495 579.445 ;
        RECT 2913.785 579.275 2913.955 579.445 ;
        RECT 5.665 573.835 5.835 574.005 ;
        RECT 6.125 573.835 6.295 574.005 ;
        RECT 6.585 573.835 6.755 574.005 ;
        RECT 2910.105 573.835 2910.275 574.005 ;
        RECT 2912.865 573.835 2913.035 574.005 ;
        RECT 2913.325 573.835 2913.495 574.005 ;
        RECT 2913.785 573.835 2913.955 574.005 ;
        RECT 5.665 568.395 5.835 568.565 ;
        RECT 6.125 568.395 6.295 568.565 ;
        RECT 6.585 568.395 6.755 568.565 ;
        RECT 2910.105 568.395 2910.275 568.565 ;
        RECT 2912.865 568.395 2913.035 568.565 ;
        RECT 2913.325 568.395 2913.495 568.565 ;
        RECT 2913.785 568.395 2913.955 568.565 ;
        RECT 5.665 562.955 5.835 563.125 ;
        RECT 6.125 562.955 6.295 563.125 ;
        RECT 6.585 562.955 6.755 563.125 ;
        RECT 2910.105 562.955 2910.275 563.125 ;
        RECT 2912.865 562.955 2913.035 563.125 ;
        RECT 2913.325 562.955 2913.495 563.125 ;
        RECT 2913.785 562.955 2913.955 563.125 ;
        RECT 5.665 557.515 5.835 557.685 ;
        RECT 6.125 557.515 6.295 557.685 ;
        RECT 6.585 557.515 6.755 557.685 ;
        RECT 2910.105 557.515 2910.275 557.685 ;
        RECT 2912.865 557.515 2913.035 557.685 ;
        RECT 2913.325 557.515 2913.495 557.685 ;
        RECT 2913.785 557.515 2913.955 557.685 ;
        RECT 5.665 552.075 5.835 552.245 ;
        RECT 6.125 552.075 6.295 552.245 ;
        RECT 6.585 552.075 6.755 552.245 ;
        RECT 2910.105 552.075 2910.275 552.245 ;
        RECT 2912.865 552.075 2913.035 552.245 ;
        RECT 2913.325 552.075 2913.495 552.245 ;
        RECT 2913.785 552.075 2913.955 552.245 ;
        RECT 5.665 546.635 5.835 546.805 ;
        RECT 6.125 546.635 6.295 546.805 ;
        RECT 6.585 546.635 6.755 546.805 ;
        RECT 2910.105 546.635 2910.275 546.805 ;
        RECT 2912.865 546.635 2913.035 546.805 ;
        RECT 2913.325 546.635 2913.495 546.805 ;
        RECT 2913.785 546.635 2913.955 546.805 ;
        RECT 5.665 541.195 5.835 541.365 ;
        RECT 6.125 541.195 6.295 541.365 ;
        RECT 6.585 541.195 6.755 541.365 ;
        RECT 2910.105 541.195 2910.275 541.365 ;
        RECT 2912.865 541.195 2913.035 541.365 ;
        RECT 2913.325 541.195 2913.495 541.365 ;
        RECT 2913.785 541.195 2913.955 541.365 ;
        RECT 5.665 535.755 5.835 535.925 ;
        RECT 6.125 535.755 6.295 535.925 ;
        RECT 6.585 535.755 6.755 535.925 ;
        RECT 2910.105 535.755 2910.275 535.925 ;
        RECT 2912.865 535.755 2913.035 535.925 ;
        RECT 2913.325 535.755 2913.495 535.925 ;
        RECT 2913.785 535.755 2913.955 535.925 ;
        RECT 5.665 530.315 5.835 530.485 ;
        RECT 6.125 530.315 6.295 530.485 ;
        RECT 6.585 530.315 6.755 530.485 ;
        RECT 2910.105 530.315 2910.275 530.485 ;
        RECT 2912.865 530.315 2913.035 530.485 ;
        RECT 2913.325 530.315 2913.495 530.485 ;
        RECT 2913.785 530.315 2913.955 530.485 ;
        RECT 5.665 524.875 5.835 525.045 ;
        RECT 6.125 524.875 6.295 525.045 ;
        RECT 6.585 524.875 6.755 525.045 ;
        RECT 2910.105 524.875 2910.275 525.045 ;
        RECT 2912.865 524.875 2913.035 525.045 ;
        RECT 2913.325 524.875 2913.495 525.045 ;
        RECT 2913.785 524.875 2913.955 525.045 ;
        RECT 5.665 519.435 5.835 519.605 ;
        RECT 6.125 519.435 6.295 519.605 ;
        RECT 6.585 519.435 6.755 519.605 ;
        RECT 2910.105 519.435 2910.275 519.605 ;
        RECT 2912.865 519.435 2913.035 519.605 ;
        RECT 2913.325 519.435 2913.495 519.605 ;
        RECT 2913.785 519.435 2913.955 519.605 ;
        RECT 5.665 513.995 5.835 514.165 ;
        RECT 6.125 513.995 6.295 514.165 ;
        RECT 6.585 513.995 6.755 514.165 ;
        RECT 2910.105 513.995 2910.275 514.165 ;
        RECT 2912.865 513.995 2913.035 514.165 ;
        RECT 2913.325 513.995 2913.495 514.165 ;
        RECT 2913.785 513.995 2913.955 514.165 ;
        RECT 5.665 508.555 5.835 508.725 ;
        RECT 6.125 508.555 6.295 508.725 ;
        RECT 6.585 508.555 6.755 508.725 ;
        RECT 2910.105 508.555 2910.275 508.725 ;
        RECT 2912.865 508.555 2913.035 508.725 ;
        RECT 2913.325 508.555 2913.495 508.725 ;
        RECT 2913.785 508.555 2913.955 508.725 ;
        RECT 5.665 503.115 5.835 503.285 ;
        RECT 6.125 503.115 6.295 503.285 ;
        RECT 6.585 503.115 6.755 503.285 ;
        RECT 2910.105 503.115 2910.275 503.285 ;
        RECT 2912.865 503.115 2913.035 503.285 ;
        RECT 2913.325 503.115 2913.495 503.285 ;
        RECT 2913.785 503.115 2913.955 503.285 ;
        RECT 5.665 497.675 5.835 497.845 ;
        RECT 6.125 497.675 6.295 497.845 ;
        RECT 6.585 497.675 6.755 497.845 ;
        RECT 2910.105 497.675 2910.275 497.845 ;
        RECT 2912.865 497.675 2913.035 497.845 ;
        RECT 2913.325 497.675 2913.495 497.845 ;
        RECT 2913.785 497.675 2913.955 497.845 ;
        RECT 5.665 492.235 5.835 492.405 ;
        RECT 6.125 492.235 6.295 492.405 ;
        RECT 6.585 492.235 6.755 492.405 ;
        RECT 2910.105 492.235 2910.275 492.405 ;
        RECT 2912.865 492.235 2913.035 492.405 ;
        RECT 2913.325 492.235 2913.495 492.405 ;
        RECT 2913.785 492.235 2913.955 492.405 ;
        RECT 5.665 486.795 5.835 486.965 ;
        RECT 6.125 486.795 6.295 486.965 ;
        RECT 6.585 486.795 6.755 486.965 ;
        RECT 2910.105 486.795 2910.275 486.965 ;
        RECT 2912.865 486.795 2913.035 486.965 ;
        RECT 2913.325 486.795 2913.495 486.965 ;
        RECT 2913.785 486.795 2913.955 486.965 ;
        RECT 5.665 481.355 5.835 481.525 ;
        RECT 6.125 481.355 6.295 481.525 ;
        RECT 6.585 481.355 6.755 481.525 ;
        RECT 2910.105 481.355 2910.275 481.525 ;
        RECT 2912.865 481.355 2913.035 481.525 ;
        RECT 2913.325 481.355 2913.495 481.525 ;
        RECT 2913.785 481.355 2913.955 481.525 ;
        RECT 5.665 475.915 5.835 476.085 ;
        RECT 6.125 475.915 6.295 476.085 ;
        RECT 6.585 475.915 6.755 476.085 ;
        RECT 2910.105 475.915 2910.275 476.085 ;
        RECT 2912.865 475.915 2913.035 476.085 ;
        RECT 2913.325 475.915 2913.495 476.085 ;
        RECT 2913.785 475.915 2913.955 476.085 ;
        RECT 5.665 470.475 5.835 470.645 ;
        RECT 6.125 470.475 6.295 470.645 ;
        RECT 6.585 470.475 6.755 470.645 ;
        RECT 2909.185 470.475 2909.355 470.645 ;
        RECT 2909.645 470.475 2909.815 470.645 ;
        RECT 2910.105 470.475 2910.275 470.645 ;
        RECT 2912.865 470.475 2913.035 470.645 ;
        RECT 2913.325 470.475 2913.495 470.645 ;
        RECT 2913.785 470.475 2913.955 470.645 ;
        RECT 5.665 465.035 5.835 465.205 ;
        RECT 6.125 465.035 6.295 465.205 ;
        RECT 6.585 465.035 6.755 465.205 ;
        RECT 2910.105 465.035 2910.275 465.205 ;
        RECT 2912.865 465.035 2913.035 465.205 ;
        RECT 2913.325 465.035 2913.495 465.205 ;
        RECT 2913.785 465.035 2913.955 465.205 ;
        RECT 5.665 459.595 5.835 459.765 ;
        RECT 6.125 459.595 6.295 459.765 ;
        RECT 6.585 459.595 6.755 459.765 ;
        RECT 2910.105 459.595 2910.275 459.765 ;
        RECT 2912.865 459.595 2913.035 459.765 ;
        RECT 2913.325 459.595 2913.495 459.765 ;
        RECT 2913.785 459.595 2913.955 459.765 ;
        RECT 5.665 454.155 5.835 454.325 ;
        RECT 6.125 454.155 6.295 454.325 ;
        RECT 6.585 454.155 6.755 454.325 ;
        RECT 2910.105 454.155 2910.275 454.325 ;
        RECT 2912.865 454.155 2913.035 454.325 ;
        RECT 2913.325 454.155 2913.495 454.325 ;
        RECT 2913.785 454.155 2913.955 454.325 ;
        RECT 5.665 448.715 5.835 448.885 ;
        RECT 6.125 448.715 6.295 448.885 ;
        RECT 6.585 448.715 6.755 448.885 ;
        RECT 2910.105 448.715 2910.275 448.885 ;
        RECT 2910.565 448.715 2910.735 448.885 ;
        RECT 2911.025 448.715 2911.195 448.885 ;
        RECT 2911.485 448.715 2911.655 448.885 ;
        RECT 2912.865 448.715 2913.035 448.885 ;
        RECT 2913.325 448.715 2913.495 448.885 ;
        RECT 2913.785 448.715 2913.955 448.885 ;
        RECT 5.665 443.275 5.835 443.445 ;
        RECT 6.125 443.275 6.295 443.445 ;
        RECT 6.585 443.275 6.755 443.445 ;
        RECT 8.885 443.275 9.055 443.445 ;
        RECT 9.345 443.275 9.515 443.445 ;
        RECT 9.805 443.275 9.975 443.445 ;
        RECT 2910.105 443.275 2910.275 443.445 ;
        RECT 2912.865 443.275 2913.035 443.445 ;
        RECT 2913.325 443.275 2913.495 443.445 ;
        RECT 2913.785 443.275 2913.955 443.445 ;
        RECT 5.665 437.835 5.835 438.005 ;
        RECT 6.125 437.835 6.295 438.005 ;
        RECT 6.585 437.835 6.755 438.005 ;
        RECT 8.885 437.835 9.055 438.005 ;
        RECT 9.345 437.835 9.515 438.005 ;
        RECT 9.805 437.835 9.975 438.005 ;
        RECT 2910.105 437.835 2910.275 438.005 ;
        RECT 2912.865 437.835 2913.035 438.005 ;
        RECT 2913.325 437.835 2913.495 438.005 ;
        RECT 2913.785 437.835 2913.955 438.005 ;
        RECT 5.665 432.395 5.835 432.565 ;
        RECT 6.125 432.395 6.295 432.565 ;
        RECT 6.585 432.395 6.755 432.565 ;
        RECT 2910.105 432.395 2910.275 432.565 ;
        RECT 2912.865 432.395 2913.035 432.565 ;
        RECT 2913.325 432.395 2913.495 432.565 ;
        RECT 2913.785 432.395 2913.955 432.565 ;
        RECT 5.665 426.955 5.835 427.125 ;
        RECT 6.125 426.955 6.295 427.125 ;
        RECT 6.585 426.955 6.755 427.125 ;
        RECT 2910.105 426.955 2910.275 427.125 ;
        RECT 2912.865 426.955 2913.035 427.125 ;
        RECT 2913.325 426.955 2913.495 427.125 ;
        RECT 2913.785 426.955 2913.955 427.125 ;
        RECT 5.665 421.515 5.835 421.685 ;
        RECT 6.125 421.515 6.295 421.685 ;
        RECT 6.585 421.515 6.755 421.685 ;
        RECT 2910.105 421.515 2910.275 421.685 ;
        RECT 2912.865 421.515 2913.035 421.685 ;
        RECT 2913.325 421.515 2913.495 421.685 ;
        RECT 2913.785 421.515 2913.955 421.685 ;
        RECT 5.665 416.075 5.835 416.245 ;
        RECT 6.125 416.075 6.295 416.245 ;
        RECT 6.585 416.075 6.755 416.245 ;
        RECT 2910.105 416.075 2910.275 416.245 ;
        RECT 2912.865 416.075 2913.035 416.245 ;
        RECT 2913.325 416.075 2913.495 416.245 ;
        RECT 2913.785 416.075 2913.955 416.245 ;
        RECT 5.665 410.635 5.835 410.805 ;
        RECT 6.125 410.635 6.295 410.805 ;
        RECT 6.585 410.635 6.755 410.805 ;
        RECT 2910.105 410.635 2910.275 410.805 ;
        RECT 2912.865 410.635 2913.035 410.805 ;
        RECT 2913.325 410.635 2913.495 410.805 ;
        RECT 2913.785 410.635 2913.955 410.805 ;
        RECT 5.665 405.195 5.835 405.365 ;
        RECT 6.125 405.195 6.295 405.365 ;
        RECT 6.585 405.195 6.755 405.365 ;
        RECT 2910.105 405.195 2910.275 405.365 ;
        RECT 2912.865 405.195 2913.035 405.365 ;
        RECT 2913.325 405.195 2913.495 405.365 ;
        RECT 2913.785 405.195 2913.955 405.365 ;
        RECT 5.665 399.755 5.835 399.925 ;
        RECT 6.125 399.755 6.295 399.925 ;
        RECT 6.585 399.755 6.755 399.925 ;
        RECT 8.885 399.755 9.055 399.925 ;
        RECT 9.345 399.755 9.515 399.925 ;
        RECT 9.805 399.755 9.975 399.925 ;
        RECT 2910.105 399.755 2910.275 399.925 ;
        RECT 2912.865 399.755 2913.035 399.925 ;
        RECT 2913.325 399.755 2913.495 399.925 ;
        RECT 2913.785 399.755 2913.955 399.925 ;
        RECT 5.665 394.315 5.835 394.485 ;
        RECT 6.125 394.315 6.295 394.485 ;
        RECT 6.585 394.315 6.755 394.485 ;
        RECT 8.885 394.315 9.055 394.485 ;
        RECT 9.345 394.315 9.515 394.485 ;
        RECT 9.805 394.315 9.975 394.485 ;
        RECT 2910.105 394.315 2910.275 394.485 ;
        RECT 2912.865 394.315 2913.035 394.485 ;
        RECT 2913.325 394.315 2913.495 394.485 ;
        RECT 2913.785 394.315 2913.955 394.485 ;
        RECT 5.665 388.875 5.835 389.045 ;
        RECT 6.125 388.875 6.295 389.045 ;
        RECT 6.585 388.875 6.755 389.045 ;
        RECT 2910.105 388.875 2910.275 389.045 ;
        RECT 2912.865 388.875 2913.035 389.045 ;
        RECT 2913.325 388.875 2913.495 389.045 ;
        RECT 2913.785 388.875 2913.955 389.045 ;
        RECT 5.665 383.435 5.835 383.605 ;
        RECT 6.125 383.435 6.295 383.605 ;
        RECT 6.585 383.435 6.755 383.605 ;
        RECT 2910.105 383.435 2910.275 383.605 ;
        RECT 2912.865 383.435 2913.035 383.605 ;
        RECT 2913.325 383.435 2913.495 383.605 ;
        RECT 2913.785 383.435 2913.955 383.605 ;
        RECT 5.665 377.995 5.835 378.165 ;
        RECT 6.125 377.995 6.295 378.165 ;
        RECT 6.585 377.995 6.755 378.165 ;
        RECT 2910.105 377.995 2910.275 378.165 ;
        RECT 2912.865 377.995 2913.035 378.165 ;
        RECT 2913.325 377.995 2913.495 378.165 ;
        RECT 2913.785 377.995 2913.955 378.165 ;
        RECT 5.665 372.555 5.835 372.725 ;
        RECT 6.125 372.555 6.295 372.725 ;
        RECT 6.585 372.555 6.755 372.725 ;
        RECT 2910.105 372.555 2910.275 372.725 ;
        RECT 2912.865 372.555 2913.035 372.725 ;
        RECT 2913.325 372.555 2913.495 372.725 ;
        RECT 2913.785 372.555 2913.955 372.725 ;
        RECT 5.665 367.115 5.835 367.285 ;
        RECT 6.125 367.115 6.295 367.285 ;
        RECT 6.585 367.115 6.755 367.285 ;
        RECT 2910.105 367.115 2910.275 367.285 ;
        RECT 2912.865 367.115 2913.035 367.285 ;
        RECT 2913.325 367.115 2913.495 367.285 ;
        RECT 2913.785 367.115 2913.955 367.285 ;
        RECT 5.665 361.675 5.835 361.845 ;
        RECT 6.125 361.675 6.295 361.845 ;
        RECT 6.585 361.675 6.755 361.845 ;
        RECT 2910.105 361.675 2910.275 361.845 ;
        RECT 2912.865 361.675 2913.035 361.845 ;
        RECT 2913.325 361.675 2913.495 361.845 ;
        RECT 2913.785 361.675 2913.955 361.845 ;
        RECT 5.665 356.235 5.835 356.405 ;
        RECT 6.125 356.235 6.295 356.405 ;
        RECT 6.585 356.235 6.755 356.405 ;
        RECT 2910.105 356.235 2910.275 356.405 ;
        RECT 2912.865 356.235 2913.035 356.405 ;
        RECT 2913.325 356.235 2913.495 356.405 ;
        RECT 2913.785 356.235 2913.955 356.405 ;
        RECT 5.665 350.795 5.835 350.965 ;
        RECT 6.125 350.795 6.295 350.965 ;
        RECT 6.585 350.795 6.755 350.965 ;
        RECT 2910.105 350.795 2910.275 350.965 ;
        RECT 2912.865 350.795 2913.035 350.965 ;
        RECT 2913.325 350.795 2913.495 350.965 ;
        RECT 2913.785 350.795 2913.955 350.965 ;
        RECT 5.665 345.355 5.835 345.525 ;
        RECT 6.125 345.355 6.295 345.525 ;
        RECT 6.585 345.355 6.755 345.525 ;
        RECT 2910.105 345.355 2910.275 345.525 ;
        RECT 2912.865 345.355 2913.035 345.525 ;
        RECT 2913.325 345.355 2913.495 345.525 ;
        RECT 2913.785 345.355 2913.955 345.525 ;
        RECT 5.665 339.915 5.835 340.085 ;
        RECT 6.125 339.915 6.295 340.085 ;
        RECT 6.585 339.915 6.755 340.085 ;
        RECT 2910.105 339.915 2910.275 340.085 ;
        RECT 2912.865 339.915 2913.035 340.085 ;
        RECT 2913.325 339.915 2913.495 340.085 ;
        RECT 2913.785 339.915 2913.955 340.085 ;
        RECT 5.665 334.475 5.835 334.645 ;
        RECT 6.125 334.475 6.295 334.645 ;
        RECT 6.585 334.475 6.755 334.645 ;
        RECT 2910.105 334.475 2910.275 334.645 ;
        RECT 2912.865 334.475 2913.035 334.645 ;
        RECT 2913.325 334.475 2913.495 334.645 ;
        RECT 2913.785 334.475 2913.955 334.645 ;
        RECT 5.665 329.035 5.835 329.205 ;
        RECT 6.125 329.035 6.295 329.205 ;
        RECT 6.585 329.035 6.755 329.205 ;
        RECT 2910.105 329.035 2910.275 329.205 ;
        RECT 2912.865 329.035 2913.035 329.205 ;
        RECT 2913.325 329.035 2913.495 329.205 ;
        RECT 2913.785 329.035 2913.955 329.205 ;
        RECT 5.665 323.595 5.835 323.765 ;
        RECT 6.125 323.595 6.295 323.765 ;
        RECT 6.585 323.595 6.755 323.765 ;
        RECT 2910.105 323.595 2910.275 323.765 ;
        RECT 2912.865 323.595 2913.035 323.765 ;
        RECT 2913.325 323.595 2913.495 323.765 ;
        RECT 2913.785 323.595 2913.955 323.765 ;
        RECT 5.665 318.155 5.835 318.325 ;
        RECT 6.125 318.155 6.295 318.325 ;
        RECT 6.585 318.155 6.755 318.325 ;
        RECT 2910.105 318.155 2910.275 318.325 ;
        RECT 2912.865 318.155 2913.035 318.325 ;
        RECT 2913.325 318.155 2913.495 318.325 ;
        RECT 2913.785 318.155 2913.955 318.325 ;
        RECT 5.665 312.715 5.835 312.885 ;
        RECT 6.125 312.715 6.295 312.885 ;
        RECT 6.585 312.715 6.755 312.885 ;
        RECT 8.885 312.715 9.055 312.885 ;
        RECT 9.345 312.715 9.515 312.885 ;
        RECT 9.805 312.715 9.975 312.885 ;
        RECT 2910.105 312.715 2910.275 312.885 ;
        RECT 2912.865 312.715 2913.035 312.885 ;
        RECT 2913.325 312.715 2913.495 312.885 ;
        RECT 2913.785 312.715 2913.955 312.885 ;
        RECT 5.665 307.275 5.835 307.445 ;
        RECT 6.125 307.275 6.295 307.445 ;
        RECT 6.585 307.275 6.755 307.445 ;
        RECT 2910.105 307.275 2910.275 307.445 ;
        RECT 2912.865 307.275 2913.035 307.445 ;
        RECT 2913.325 307.275 2913.495 307.445 ;
        RECT 2913.785 307.275 2913.955 307.445 ;
        RECT 5.665 301.835 5.835 302.005 ;
        RECT 6.125 301.835 6.295 302.005 ;
        RECT 6.585 301.835 6.755 302.005 ;
        RECT 2910.105 301.835 2910.275 302.005 ;
        RECT 2912.865 301.835 2913.035 302.005 ;
        RECT 2913.325 301.835 2913.495 302.005 ;
        RECT 2913.785 301.835 2913.955 302.005 ;
        RECT 5.665 296.395 5.835 296.565 ;
        RECT 6.125 296.395 6.295 296.565 ;
        RECT 6.585 296.395 6.755 296.565 ;
        RECT 2910.105 296.395 2910.275 296.565 ;
        RECT 2912.865 296.395 2913.035 296.565 ;
        RECT 2913.325 296.395 2913.495 296.565 ;
        RECT 2913.785 296.395 2913.955 296.565 ;
        RECT 5.665 290.955 5.835 291.125 ;
        RECT 6.125 290.955 6.295 291.125 ;
        RECT 6.585 290.955 6.755 291.125 ;
        RECT 2909.185 290.955 2909.355 291.125 ;
        RECT 2909.645 290.955 2909.815 291.125 ;
        RECT 2910.105 290.955 2910.275 291.125 ;
        RECT 2912.865 290.955 2913.035 291.125 ;
        RECT 2913.325 290.955 2913.495 291.125 ;
        RECT 2913.785 290.955 2913.955 291.125 ;
        RECT 5.665 285.515 5.835 285.685 ;
        RECT 6.125 285.515 6.295 285.685 ;
        RECT 6.585 285.515 6.755 285.685 ;
        RECT 2910.105 285.515 2910.275 285.685 ;
        RECT 2912.865 285.515 2913.035 285.685 ;
        RECT 2913.325 285.515 2913.495 285.685 ;
        RECT 2913.785 285.515 2913.955 285.685 ;
        RECT 5.665 280.075 5.835 280.245 ;
        RECT 6.125 280.075 6.295 280.245 ;
        RECT 6.585 280.075 6.755 280.245 ;
        RECT 2910.105 280.075 2910.275 280.245 ;
        RECT 2912.865 280.075 2913.035 280.245 ;
        RECT 2913.325 280.075 2913.495 280.245 ;
        RECT 2913.785 280.075 2913.955 280.245 ;
        RECT 5.665 274.635 5.835 274.805 ;
        RECT 6.125 274.635 6.295 274.805 ;
        RECT 6.585 274.635 6.755 274.805 ;
        RECT 2910.105 274.635 2910.275 274.805 ;
        RECT 2912.865 274.635 2913.035 274.805 ;
        RECT 2913.325 274.635 2913.495 274.805 ;
        RECT 2913.785 274.635 2913.955 274.805 ;
        RECT 5.665 269.195 5.835 269.365 ;
        RECT 6.125 269.195 6.295 269.365 ;
        RECT 6.585 269.195 6.755 269.365 ;
        RECT 2910.105 269.195 2910.275 269.365 ;
        RECT 2912.865 269.195 2913.035 269.365 ;
        RECT 2913.325 269.195 2913.495 269.365 ;
        RECT 2913.785 269.195 2913.955 269.365 ;
        RECT 5.665 263.755 5.835 263.925 ;
        RECT 6.125 263.755 6.295 263.925 ;
        RECT 6.585 263.755 6.755 263.925 ;
        RECT 2910.105 263.755 2910.275 263.925 ;
        RECT 2912.865 263.755 2913.035 263.925 ;
        RECT 2913.325 263.755 2913.495 263.925 ;
        RECT 2913.785 263.755 2913.955 263.925 ;
        RECT 5.665 258.315 5.835 258.485 ;
        RECT 6.125 258.315 6.295 258.485 ;
        RECT 6.585 258.315 6.755 258.485 ;
        RECT 2910.105 258.315 2910.275 258.485 ;
        RECT 2912.865 258.315 2913.035 258.485 ;
        RECT 2913.325 258.315 2913.495 258.485 ;
        RECT 2913.785 258.315 2913.955 258.485 ;
        RECT 5.665 252.875 5.835 253.045 ;
        RECT 6.125 252.875 6.295 253.045 ;
        RECT 6.585 252.875 6.755 253.045 ;
        RECT 2910.105 252.875 2910.275 253.045 ;
        RECT 2912.865 252.875 2913.035 253.045 ;
        RECT 2913.325 252.875 2913.495 253.045 ;
        RECT 2913.785 252.875 2913.955 253.045 ;
        RECT 5.665 247.435 5.835 247.605 ;
        RECT 6.125 247.435 6.295 247.605 ;
        RECT 6.585 247.435 6.755 247.605 ;
        RECT 2910.105 247.435 2910.275 247.605 ;
        RECT 2912.865 247.435 2913.035 247.605 ;
        RECT 2913.325 247.435 2913.495 247.605 ;
        RECT 2913.785 247.435 2913.955 247.605 ;
        RECT 5.665 241.995 5.835 242.165 ;
        RECT 6.125 241.995 6.295 242.165 ;
        RECT 6.585 241.995 6.755 242.165 ;
        RECT 2910.105 241.995 2910.275 242.165 ;
        RECT 2912.865 241.995 2913.035 242.165 ;
        RECT 2913.325 241.995 2913.495 242.165 ;
        RECT 2913.785 241.995 2913.955 242.165 ;
        RECT 5.665 236.555 5.835 236.725 ;
        RECT 6.125 236.555 6.295 236.725 ;
        RECT 6.585 236.555 6.755 236.725 ;
        RECT 2910.105 236.555 2910.275 236.725 ;
        RECT 2912.865 236.555 2913.035 236.725 ;
        RECT 2913.325 236.555 2913.495 236.725 ;
        RECT 2913.785 236.555 2913.955 236.725 ;
        RECT 5.665 231.115 5.835 231.285 ;
        RECT 6.125 231.115 6.295 231.285 ;
        RECT 6.585 231.115 6.755 231.285 ;
        RECT 2910.105 231.115 2910.275 231.285 ;
        RECT 2910.565 231.115 2910.735 231.285 ;
        RECT 2911.025 231.115 2911.195 231.285 ;
        RECT 2911.485 231.115 2911.655 231.285 ;
        RECT 2912.865 231.115 2913.035 231.285 ;
        RECT 2913.325 231.115 2913.495 231.285 ;
        RECT 2913.785 231.115 2913.955 231.285 ;
        RECT 5.665 225.675 5.835 225.845 ;
        RECT 6.125 225.675 6.295 225.845 ;
        RECT 6.585 225.675 6.755 225.845 ;
        RECT 2910.105 225.675 2910.275 225.845 ;
        RECT 2912.865 225.675 2913.035 225.845 ;
        RECT 2913.325 225.675 2913.495 225.845 ;
        RECT 2913.785 225.675 2913.955 225.845 ;
        RECT 5.665 220.235 5.835 220.405 ;
        RECT 6.125 220.235 6.295 220.405 ;
        RECT 6.585 220.235 6.755 220.405 ;
        RECT 2910.105 220.235 2910.275 220.405 ;
        RECT 2912.865 220.235 2913.035 220.405 ;
        RECT 2913.325 220.235 2913.495 220.405 ;
        RECT 2913.785 220.235 2913.955 220.405 ;
        RECT 5.665 214.795 5.835 214.965 ;
        RECT 6.125 214.795 6.295 214.965 ;
        RECT 6.585 214.795 6.755 214.965 ;
        RECT 2910.105 214.795 2910.275 214.965 ;
        RECT 2912.865 214.795 2913.035 214.965 ;
        RECT 2913.325 214.795 2913.495 214.965 ;
        RECT 2913.785 214.795 2913.955 214.965 ;
        RECT 5.665 209.355 5.835 209.525 ;
        RECT 6.125 209.355 6.295 209.525 ;
        RECT 6.585 209.355 6.755 209.525 ;
        RECT 2910.105 209.355 2910.275 209.525 ;
        RECT 2912.865 209.355 2913.035 209.525 ;
        RECT 2913.325 209.355 2913.495 209.525 ;
        RECT 2913.785 209.355 2913.955 209.525 ;
        RECT 5.665 203.915 5.835 204.085 ;
        RECT 6.125 203.915 6.295 204.085 ;
        RECT 6.585 203.915 6.755 204.085 ;
        RECT 2910.105 203.915 2910.275 204.085 ;
        RECT 2912.865 203.915 2913.035 204.085 ;
        RECT 2913.325 203.915 2913.495 204.085 ;
        RECT 2913.785 203.915 2913.955 204.085 ;
        RECT 5.665 198.475 5.835 198.645 ;
        RECT 6.125 198.475 6.295 198.645 ;
        RECT 6.585 198.475 6.755 198.645 ;
        RECT 2910.105 198.475 2910.275 198.645 ;
        RECT 2912.865 198.475 2913.035 198.645 ;
        RECT 2913.325 198.475 2913.495 198.645 ;
        RECT 2913.785 198.475 2913.955 198.645 ;
        RECT 5.665 193.035 5.835 193.205 ;
        RECT 6.125 193.035 6.295 193.205 ;
        RECT 6.585 193.035 6.755 193.205 ;
        RECT 2910.105 193.035 2910.275 193.205 ;
        RECT 2912.865 193.035 2913.035 193.205 ;
        RECT 2913.325 193.035 2913.495 193.205 ;
        RECT 2913.785 193.035 2913.955 193.205 ;
        RECT 5.665 187.595 5.835 187.765 ;
        RECT 6.125 187.595 6.295 187.765 ;
        RECT 6.585 187.595 6.755 187.765 ;
        RECT 2910.105 187.595 2910.275 187.765 ;
        RECT 2912.865 187.595 2913.035 187.765 ;
        RECT 2913.325 187.595 2913.495 187.765 ;
        RECT 2913.785 187.595 2913.955 187.765 ;
        RECT 5.665 182.155 5.835 182.325 ;
        RECT 6.125 182.155 6.295 182.325 ;
        RECT 6.585 182.155 6.755 182.325 ;
        RECT 2910.105 182.155 2910.275 182.325 ;
        RECT 2912.865 182.155 2913.035 182.325 ;
        RECT 2913.325 182.155 2913.495 182.325 ;
        RECT 2913.785 182.155 2913.955 182.325 ;
        RECT 5.665 176.715 5.835 176.885 ;
        RECT 6.125 176.715 6.295 176.885 ;
        RECT 6.585 176.715 6.755 176.885 ;
        RECT 2910.105 176.715 2910.275 176.885 ;
        RECT 2912.865 176.715 2913.035 176.885 ;
        RECT 2913.325 176.715 2913.495 176.885 ;
        RECT 2913.785 176.715 2913.955 176.885 ;
        RECT 5.665 171.275 5.835 171.445 ;
        RECT 6.125 171.275 6.295 171.445 ;
        RECT 6.585 171.275 6.755 171.445 ;
        RECT 2910.105 171.275 2910.275 171.445 ;
        RECT 2912.865 171.275 2913.035 171.445 ;
        RECT 2913.325 171.275 2913.495 171.445 ;
        RECT 2913.785 171.275 2913.955 171.445 ;
        RECT 5.665 165.835 5.835 166.005 ;
        RECT 6.125 165.835 6.295 166.005 ;
        RECT 6.585 165.835 6.755 166.005 ;
        RECT 2910.105 165.835 2910.275 166.005 ;
        RECT 2912.865 165.835 2913.035 166.005 ;
        RECT 2913.325 165.835 2913.495 166.005 ;
        RECT 2913.785 165.835 2913.955 166.005 ;
        RECT 5.665 160.395 5.835 160.565 ;
        RECT 6.125 160.395 6.295 160.565 ;
        RECT 6.585 160.395 6.755 160.565 ;
        RECT 2910.105 160.395 2910.275 160.565 ;
        RECT 2912.865 160.395 2913.035 160.565 ;
        RECT 2913.325 160.395 2913.495 160.565 ;
        RECT 2913.785 160.395 2913.955 160.565 ;
        RECT 5.665 154.955 5.835 155.125 ;
        RECT 6.125 154.955 6.295 155.125 ;
        RECT 6.585 154.955 6.755 155.125 ;
        RECT 2910.105 154.955 2910.275 155.125 ;
        RECT 2912.865 154.955 2913.035 155.125 ;
        RECT 2913.325 154.955 2913.495 155.125 ;
        RECT 2913.785 154.955 2913.955 155.125 ;
        RECT 5.665 149.515 5.835 149.685 ;
        RECT 6.125 149.515 6.295 149.685 ;
        RECT 6.585 149.515 6.755 149.685 ;
        RECT 2910.105 149.515 2910.275 149.685 ;
        RECT 2912.865 149.515 2913.035 149.685 ;
        RECT 2913.325 149.515 2913.495 149.685 ;
        RECT 2913.785 149.515 2913.955 149.685 ;
        RECT 5.665 144.075 5.835 144.245 ;
        RECT 6.125 144.075 6.295 144.245 ;
        RECT 6.585 144.075 6.755 144.245 ;
        RECT 2910.105 144.075 2910.275 144.245 ;
        RECT 2912.865 144.075 2913.035 144.245 ;
        RECT 2913.325 144.075 2913.495 144.245 ;
        RECT 2913.785 144.075 2913.955 144.245 ;
        RECT 5.665 138.635 5.835 138.805 ;
        RECT 6.125 138.635 6.295 138.805 ;
        RECT 6.585 138.635 6.755 138.805 ;
        RECT 2910.105 138.635 2910.275 138.805 ;
        RECT 2912.865 138.635 2913.035 138.805 ;
        RECT 2913.325 138.635 2913.495 138.805 ;
        RECT 2913.785 138.635 2913.955 138.805 ;
        RECT 5.665 133.195 5.835 133.365 ;
        RECT 6.125 133.195 6.295 133.365 ;
        RECT 6.585 133.195 6.755 133.365 ;
        RECT 2910.105 133.195 2910.275 133.365 ;
        RECT 2912.865 133.195 2913.035 133.365 ;
        RECT 2913.325 133.195 2913.495 133.365 ;
        RECT 2913.785 133.195 2913.955 133.365 ;
        RECT 5.665 127.755 5.835 127.925 ;
        RECT 6.125 127.755 6.295 127.925 ;
        RECT 6.585 127.755 6.755 127.925 ;
        RECT 7.045 127.755 7.215 127.925 ;
        RECT 7.505 127.755 7.675 127.925 ;
        RECT 7.965 127.755 8.135 127.925 ;
        RECT 8.425 127.755 8.595 127.925 ;
        RECT 8.885 127.755 9.055 127.925 ;
        RECT 9.345 127.755 9.515 127.925 ;
        RECT 9.805 127.755 9.975 127.925 ;
        RECT 10.265 127.755 10.435 127.925 ;
        RECT 10.725 127.755 10.895 127.925 ;
        RECT 11.185 127.755 11.355 127.925 ;
        RECT 11.645 127.755 11.815 127.925 ;
        RECT 12.105 127.755 12.275 127.925 ;
        RECT 12.565 127.755 12.735 127.925 ;
        RECT 13.025 127.755 13.195 127.925 ;
        RECT 13.485 127.755 13.655 127.925 ;
        RECT 2910.105 127.755 2910.275 127.925 ;
        RECT 2912.865 127.755 2913.035 127.925 ;
        RECT 2913.325 127.755 2913.495 127.925 ;
        RECT 2913.785 127.755 2913.955 127.925 ;
        RECT 5.665 122.315 5.835 122.485 ;
        RECT 6.125 122.315 6.295 122.485 ;
        RECT 6.585 122.315 6.755 122.485 ;
        RECT 2910.105 122.315 2910.275 122.485 ;
        RECT 2912.865 122.315 2913.035 122.485 ;
        RECT 2913.325 122.315 2913.495 122.485 ;
        RECT 2913.785 122.315 2913.955 122.485 ;
        RECT 5.665 116.875 5.835 117.045 ;
        RECT 6.125 116.875 6.295 117.045 ;
        RECT 6.585 116.875 6.755 117.045 ;
        RECT 2910.105 116.875 2910.275 117.045 ;
        RECT 2912.865 116.875 2913.035 117.045 ;
        RECT 2913.325 116.875 2913.495 117.045 ;
        RECT 2913.785 116.875 2913.955 117.045 ;
        RECT 5.665 111.435 5.835 111.605 ;
        RECT 6.125 111.435 6.295 111.605 ;
        RECT 6.585 111.435 6.755 111.605 ;
        RECT 2910.105 111.435 2910.275 111.605 ;
        RECT 2912.865 111.435 2913.035 111.605 ;
        RECT 2913.325 111.435 2913.495 111.605 ;
        RECT 2913.785 111.435 2913.955 111.605 ;
        RECT 5.665 105.995 5.835 106.165 ;
        RECT 6.125 105.995 6.295 106.165 ;
        RECT 6.585 105.995 6.755 106.165 ;
        RECT 8.885 105.995 9.055 106.165 ;
        RECT 9.345 105.995 9.515 106.165 ;
        RECT 9.805 105.995 9.975 106.165 ;
        RECT 2910.105 105.995 2910.275 106.165 ;
        RECT 2912.865 105.995 2913.035 106.165 ;
        RECT 2913.325 105.995 2913.495 106.165 ;
        RECT 2913.785 105.995 2913.955 106.165 ;
        RECT 5.665 100.555 5.835 100.725 ;
        RECT 6.125 100.555 6.295 100.725 ;
        RECT 6.585 100.555 6.755 100.725 ;
        RECT 2910.105 100.555 2910.275 100.725 ;
        RECT 2912.865 100.555 2913.035 100.725 ;
        RECT 2913.325 100.555 2913.495 100.725 ;
        RECT 2913.785 100.555 2913.955 100.725 ;
        RECT 5.665 95.115 5.835 95.285 ;
        RECT 6.125 95.115 6.295 95.285 ;
        RECT 6.585 95.115 6.755 95.285 ;
        RECT 2910.105 95.115 2910.275 95.285 ;
        RECT 2912.865 95.115 2913.035 95.285 ;
        RECT 2913.325 95.115 2913.495 95.285 ;
        RECT 2913.785 95.115 2913.955 95.285 ;
        RECT 5.665 89.675 5.835 89.845 ;
        RECT 6.125 89.675 6.295 89.845 ;
        RECT 6.585 89.675 6.755 89.845 ;
        RECT 2910.105 89.675 2910.275 89.845 ;
        RECT 2912.865 89.675 2913.035 89.845 ;
        RECT 2913.325 89.675 2913.495 89.845 ;
        RECT 2913.785 89.675 2913.955 89.845 ;
        RECT 5.665 84.235 5.835 84.405 ;
        RECT 6.125 84.235 6.295 84.405 ;
        RECT 6.585 84.235 6.755 84.405 ;
        RECT 2910.105 84.235 2910.275 84.405 ;
        RECT 2912.865 84.235 2913.035 84.405 ;
        RECT 2913.325 84.235 2913.495 84.405 ;
        RECT 2913.785 84.235 2913.955 84.405 ;
        RECT 5.665 78.795 5.835 78.965 ;
        RECT 6.125 78.795 6.295 78.965 ;
        RECT 6.585 78.795 6.755 78.965 ;
        RECT 2910.105 78.795 2910.275 78.965 ;
        RECT 2912.865 78.795 2913.035 78.965 ;
        RECT 2913.325 78.795 2913.495 78.965 ;
        RECT 2913.785 78.795 2913.955 78.965 ;
        RECT 5.665 73.355 5.835 73.525 ;
        RECT 6.125 73.355 6.295 73.525 ;
        RECT 6.585 73.355 6.755 73.525 ;
        RECT 2910.105 73.355 2910.275 73.525 ;
        RECT 2912.865 73.355 2913.035 73.525 ;
        RECT 2913.325 73.355 2913.495 73.525 ;
        RECT 2913.785 73.355 2913.955 73.525 ;
        RECT 5.665 67.915 5.835 68.085 ;
        RECT 6.125 67.915 6.295 68.085 ;
        RECT 6.585 67.915 6.755 68.085 ;
        RECT 2910.105 67.915 2910.275 68.085 ;
        RECT 2912.865 67.915 2913.035 68.085 ;
        RECT 2913.325 67.915 2913.495 68.085 ;
        RECT 2913.785 67.915 2913.955 68.085 ;
        RECT 5.665 62.475 5.835 62.645 ;
        RECT 6.125 62.475 6.295 62.645 ;
        RECT 6.585 62.475 6.755 62.645 ;
        RECT 2909.185 62.475 2909.355 62.645 ;
        RECT 2909.645 62.475 2909.815 62.645 ;
        RECT 2910.105 62.475 2910.275 62.645 ;
        RECT 2912.865 62.475 2913.035 62.645 ;
        RECT 2913.325 62.475 2913.495 62.645 ;
        RECT 2913.785 62.475 2913.955 62.645 ;
        RECT 5.665 57.035 5.835 57.205 ;
        RECT 6.125 57.035 6.295 57.205 ;
        RECT 6.585 57.035 6.755 57.205 ;
        RECT 2910.105 57.035 2910.275 57.205 ;
        RECT 2912.865 57.035 2913.035 57.205 ;
        RECT 2913.325 57.035 2913.495 57.205 ;
        RECT 2913.785 57.035 2913.955 57.205 ;
        RECT 5.665 51.595 5.835 51.765 ;
        RECT 6.125 51.595 6.295 51.765 ;
        RECT 6.585 51.595 6.755 51.765 ;
        RECT 2910.105 51.595 2910.275 51.765 ;
        RECT 2912.865 51.595 2913.035 51.765 ;
        RECT 2913.325 51.595 2913.495 51.765 ;
        RECT 2913.785 51.595 2913.955 51.765 ;
        RECT 5.665 46.155 5.835 46.325 ;
        RECT 6.125 46.155 6.295 46.325 ;
        RECT 6.585 46.155 6.755 46.325 ;
        RECT 2910.105 46.155 2910.275 46.325 ;
        RECT 2912.865 46.155 2913.035 46.325 ;
        RECT 2913.325 46.155 2913.495 46.325 ;
        RECT 2913.785 46.155 2913.955 46.325 ;
        RECT 5.665 40.715 5.835 40.885 ;
        RECT 6.125 40.715 6.295 40.885 ;
        RECT 6.585 40.715 6.755 40.885 ;
        RECT 7.045 40.715 7.215 40.885 ;
        RECT 7.505 40.715 7.675 40.885 ;
        RECT 7.965 40.715 8.135 40.885 ;
        RECT 8.425 40.715 8.595 40.885 ;
        RECT 8.885 40.715 9.055 40.885 ;
        RECT 9.345 40.715 9.515 40.885 ;
        RECT 9.805 40.715 9.975 40.885 ;
        RECT 10.265 40.715 10.435 40.885 ;
        RECT 10.725 40.715 10.895 40.885 ;
        RECT 11.185 40.715 11.355 40.885 ;
        RECT 11.645 40.715 11.815 40.885 ;
        RECT 12.105 40.715 12.275 40.885 ;
        RECT 12.565 40.715 12.735 40.885 ;
        RECT 13.025 40.715 13.195 40.885 ;
        RECT 13.485 40.715 13.655 40.885 ;
        RECT 2910.105 40.715 2910.275 40.885 ;
        RECT 2912.865 40.715 2913.035 40.885 ;
        RECT 2913.325 40.715 2913.495 40.885 ;
        RECT 2913.785 40.715 2913.955 40.885 ;
        RECT 5.665 35.275 5.835 35.445 ;
        RECT 6.125 35.275 6.295 35.445 ;
        RECT 6.585 35.275 6.755 35.445 ;
        RECT 2910.105 35.275 2910.275 35.445 ;
        RECT 2912.865 35.275 2913.035 35.445 ;
        RECT 2913.325 35.275 2913.495 35.445 ;
        RECT 2913.785 35.275 2913.955 35.445 ;
        RECT 5.665 29.835 5.835 30.005 ;
        RECT 6.125 29.835 6.295 30.005 ;
        RECT 6.585 29.835 6.755 30.005 ;
        RECT 2910.105 29.835 2910.275 30.005 ;
        RECT 2912.865 29.835 2913.035 30.005 ;
        RECT 2913.325 29.835 2913.495 30.005 ;
        RECT 2913.785 29.835 2913.955 30.005 ;
        RECT 5.665 24.395 5.835 24.565 ;
        RECT 6.125 24.395 6.295 24.565 ;
        RECT 6.585 24.395 6.755 24.565 ;
        RECT 2910.105 24.395 2910.275 24.565 ;
        RECT 2912.865 24.395 2913.035 24.565 ;
        RECT 2913.325 24.395 2913.495 24.565 ;
        RECT 2913.785 24.395 2913.955 24.565 ;
        RECT 5.665 18.955 5.835 19.125 ;
        RECT 6.125 18.955 6.295 19.125 ;
        RECT 6.585 18.955 6.755 19.125 ;
        RECT 7.045 18.955 7.215 19.125 ;
        RECT 7.505 18.955 7.675 19.125 ;
        RECT 7.965 18.955 8.135 19.125 ;
        RECT 8.425 18.955 8.595 19.125 ;
        RECT 8.885 18.955 9.055 19.125 ;
        RECT 9.345 18.955 9.515 19.125 ;
        RECT 9.805 18.955 9.975 19.125 ;
        RECT 10.265 18.955 10.435 19.125 ;
        RECT 10.725 18.955 10.895 19.125 ;
        RECT 11.185 18.955 11.355 19.125 ;
        RECT 11.645 18.955 11.815 19.125 ;
        RECT 12.105 18.955 12.275 19.125 ;
        RECT 12.565 18.955 12.735 19.125 ;
        RECT 13.025 18.955 13.195 19.125 ;
        RECT 13.485 18.955 13.655 19.125 ;
        RECT 2909.185 18.955 2909.355 19.125 ;
        RECT 2909.645 18.955 2909.815 19.125 ;
        RECT 2910.105 18.955 2910.275 19.125 ;
        RECT 2910.565 18.955 2910.735 19.125 ;
        RECT 2911.025 18.955 2911.195 19.125 ;
        RECT 2911.485 18.955 2911.655 19.125 ;
        RECT 2912.865 18.955 2913.035 19.125 ;
        RECT 2913.325 18.955 2913.495 19.125 ;
        RECT 2913.785 18.955 2913.955 19.125 ;
        RECT 5.665 13.515 5.835 13.685 ;
        RECT 6.125 13.515 6.295 13.685 ;
        RECT 6.585 13.515 6.755 13.685 ;
        RECT 7.045 13.515 7.215 13.685 ;
        RECT 7.505 13.515 7.675 13.685 ;
        RECT 7.965 13.515 8.135 13.685 ;
        RECT 8.425 13.515 8.595 13.685 ;
        RECT 8.885 13.515 9.055 13.685 ;
        RECT 9.345 13.515 9.515 13.685 ;
        RECT 9.805 13.515 9.975 13.685 ;
        RECT 10.265 13.515 10.435 13.685 ;
        RECT 10.725 13.515 10.895 13.685 ;
        RECT 11.185 13.515 11.355 13.685 ;
        RECT 11.645 13.515 11.815 13.685 ;
        RECT 12.105 13.515 12.275 13.685 ;
        RECT 12.565 13.515 12.735 13.685 ;
        RECT 13.025 13.515 13.195 13.685 ;
        RECT 13.485 13.515 13.655 13.685 ;
        RECT 13.945 13.515 14.115 13.685 ;
        RECT 14.405 13.515 14.575 13.685 ;
        RECT 14.865 13.515 15.035 13.685 ;
        RECT 15.325 13.515 15.495 13.685 ;
        RECT 16.705 13.515 16.875 13.685 ;
        RECT 17.165 13.515 17.335 13.685 ;
        RECT 17.625 13.515 17.795 13.685 ;
        RECT 18.085 13.515 18.255 13.685 ;
        RECT 19.925 13.515 20.095 13.685 ;
        RECT 34.185 13.515 34.355 13.685 ;
        RECT 47.985 13.515 48.155 13.685 ;
        RECT 48.445 13.515 48.615 13.685 ;
        RECT 58.105 13.515 58.275 13.685 ;
        RECT 58.565 13.515 58.735 13.685 ;
        RECT 59.025 13.515 59.195 13.685 ;
        RECT 59.485 13.515 59.655 13.685 ;
        RECT 59.945 13.515 60.115 13.685 ;
        RECT 60.405 13.515 60.575 13.685 ;
        RECT 60.865 13.515 61.035 13.685 ;
        RECT 61.325 13.515 61.495 13.685 ;
        RECT 61.785 13.515 61.955 13.685 ;
        RECT 62.245 13.515 62.415 13.685 ;
        RECT 62.705 13.515 62.875 13.685 ;
        RECT 63.165 13.515 63.335 13.685 ;
        RECT 63.625 13.515 63.795 13.685 ;
        RECT 64.085 13.515 64.255 13.685 ;
        RECT 64.545 13.515 64.715 13.685 ;
        RECT 65.005 13.515 65.175 13.685 ;
        RECT 65.465 13.515 65.635 13.685 ;
        RECT 76.045 13.515 76.215 13.685 ;
        RECT 76.965 13.515 77.135 13.685 ;
        RECT 77.425 13.515 77.595 13.685 ;
        RECT 77.885 13.515 78.055 13.685 ;
        RECT 78.345 13.515 78.515 13.685 ;
        RECT 78.805 13.515 78.975 13.685 ;
        RECT 79.265 13.515 79.435 13.685 ;
        RECT 79.725 13.515 79.895 13.685 ;
        RECT 80.185 13.515 80.355 13.685 ;
        RECT 80.645 13.515 80.815 13.685 ;
        RECT 81.105 13.515 81.275 13.685 ;
        RECT 82.025 13.515 82.195 13.685 ;
        RECT 82.485 13.515 82.655 13.685 ;
        RECT 82.945 13.515 83.115 13.685 ;
        RECT 83.405 13.515 83.575 13.685 ;
        RECT 83.865 13.515 84.035 13.685 ;
        RECT 84.325 13.515 84.495 13.685 ;
        RECT 84.785 13.515 84.955 13.685 ;
        RECT 85.245 13.515 85.415 13.685 ;
        RECT 85.705 13.515 85.875 13.685 ;
        RECT 86.165 13.515 86.335 13.685 ;
        RECT 86.625 13.515 86.795 13.685 ;
        RECT 87.085 13.515 87.255 13.685 ;
        RECT 87.545 13.515 87.715 13.685 ;
        RECT 88.005 13.515 88.175 13.685 ;
        RECT 88.465 13.515 88.635 13.685 ;
        RECT 88.925 13.515 89.095 13.685 ;
        RECT 89.385 13.515 89.555 13.685 ;
        RECT 89.845 13.515 90.015 13.685 ;
        RECT 90.305 13.515 90.475 13.685 ;
        RECT 90.765 13.515 90.935 13.685 ;
        RECT 91.225 13.515 91.395 13.685 ;
        RECT 101.345 13.515 101.515 13.685 ;
        RECT 101.805 13.515 101.975 13.685 ;
        RECT 102.265 13.515 102.435 13.685 ;
        RECT 102.725 13.515 102.895 13.685 ;
        RECT 104.105 13.515 104.275 13.685 ;
        RECT 104.565 13.515 104.735 13.685 ;
        RECT 105.025 13.515 105.195 13.685 ;
        RECT 105.485 13.515 105.655 13.685 ;
        RECT 105.945 13.515 106.115 13.685 ;
        RECT 106.405 13.515 106.575 13.685 ;
        RECT 106.865 13.515 107.035 13.685 ;
        RECT 107.325 13.515 107.495 13.685 ;
        RECT 107.785 13.515 107.955 13.685 ;
        RECT 108.245 13.515 108.415 13.685 ;
        RECT 108.705 13.515 108.875 13.685 ;
        RECT 109.165 13.515 109.335 13.685 ;
        RECT 109.625 13.515 109.795 13.685 ;
        RECT 110.085 13.515 110.255 13.685 ;
        RECT 110.545 13.515 110.715 13.685 ;
        RECT 111.005 13.515 111.175 13.685 ;
        RECT 111.465 13.515 111.635 13.685 ;
        RECT 119.745 13.515 119.915 13.685 ;
        RECT 120.205 13.515 120.375 13.685 ;
        RECT 120.665 13.515 120.835 13.685 ;
        RECT 121.125 13.515 121.295 13.685 ;
        RECT 132.165 13.515 132.335 13.685 ;
        RECT 134.005 13.515 134.175 13.685 ;
        RECT 134.465 13.515 134.635 13.685 ;
        RECT 134.925 13.515 135.095 13.685 ;
        RECT 135.385 13.515 135.555 13.685 ;
        RECT 135.845 13.515 136.015 13.685 ;
        RECT 136.305 13.515 136.475 13.685 ;
        RECT 136.765 13.515 136.935 13.685 ;
        RECT 137.225 13.515 137.395 13.685 ;
        RECT 137.685 13.515 137.855 13.685 ;
        RECT 138.145 13.515 138.315 13.685 ;
        RECT 138.605 13.515 138.775 13.685 ;
        RECT 139.065 13.515 139.235 13.685 ;
        RECT 139.525 13.515 139.695 13.685 ;
        RECT 139.985 13.515 140.155 13.685 ;
        RECT 140.445 13.515 140.615 13.685 ;
        RECT 142.285 13.515 142.455 13.685 ;
        RECT 142.745 13.515 142.915 13.685 ;
        RECT 143.205 13.515 143.375 13.685 ;
        RECT 143.665 13.515 143.835 13.685 ;
        RECT 144.125 13.515 144.295 13.685 ;
        RECT 144.585 13.515 144.755 13.685 ;
        RECT 145.045 13.515 145.215 13.685 ;
        RECT 145.505 13.515 145.675 13.685 ;
        RECT 145.965 13.515 146.135 13.685 ;
        RECT 146.425 13.515 146.595 13.685 ;
        RECT 146.885 13.515 147.055 13.685 ;
        RECT 147.345 13.515 147.515 13.685 ;
        RECT 147.805 13.515 147.975 13.685 ;
        RECT 148.265 13.515 148.435 13.685 ;
        RECT 152.865 13.515 153.035 13.685 ;
        RECT 153.325 13.515 153.495 13.685 ;
        RECT 153.785 13.515 153.955 13.685 ;
        RECT 154.245 13.515 154.415 13.685 ;
        RECT 154.705 13.515 154.875 13.685 ;
        RECT 155.165 13.515 155.335 13.685 ;
        RECT 155.625 13.515 155.795 13.685 ;
        RECT 156.085 13.515 156.255 13.685 ;
        RECT 156.545 13.515 156.715 13.685 ;
        RECT 157.005 13.515 157.175 13.685 ;
        RECT 157.465 13.515 157.635 13.685 ;
        RECT 157.925 13.515 158.095 13.685 ;
        RECT 158.385 13.515 158.555 13.685 ;
        RECT 158.845 13.515 159.015 13.685 ;
        RECT 159.305 13.515 159.475 13.685 ;
        RECT 159.765 13.515 159.935 13.685 ;
        RECT 160.225 13.515 160.395 13.685 ;
        RECT 160.685 13.515 160.855 13.685 ;
        RECT 161.145 13.515 161.315 13.685 ;
        RECT 161.605 13.515 161.775 13.685 ;
        RECT 162.525 13.515 162.695 13.685 ;
        RECT 162.985 13.515 163.155 13.685 ;
        RECT 163.445 13.515 163.615 13.685 ;
        RECT 163.905 13.515 164.075 13.685 ;
        RECT 164.365 13.515 164.535 13.685 ;
        RECT 164.825 13.515 164.995 13.685 ;
        RECT 165.285 13.515 165.455 13.685 ;
        RECT 165.745 13.515 165.915 13.685 ;
        RECT 166.205 13.515 166.375 13.685 ;
        RECT 166.665 13.515 166.835 13.685 ;
        RECT 167.125 13.515 167.295 13.685 ;
        RECT 167.585 13.515 167.755 13.685 ;
        RECT 168.045 13.515 168.215 13.685 ;
        RECT 168.505 13.515 168.675 13.685 ;
        RECT 168.965 13.515 169.135 13.685 ;
        RECT 169.425 13.515 169.595 13.685 ;
        RECT 169.885 13.515 170.055 13.685 ;
        RECT 170.345 13.515 170.515 13.685 ;
        RECT 170.805 13.515 170.975 13.685 ;
        RECT 176.785 13.515 176.955 13.685 ;
        RECT 181.385 13.515 181.555 13.685 ;
        RECT 181.845 13.515 182.015 13.685 ;
        RECT 182.305 13.515 182.475 13.685 ;
        RECT 182.765 13.515 182.935 13.685 ;
        RECT 183.225 13.515 183.395 13.685 ;
        RECT 183.685 13.515 183.855 13.685 ;
        RECT 184.145 13.515 184.315 13.685 ;
        RECT 184.605 13.515 184.775 13.685 ;
        RECT 185.065 13.515 185.235 13.685 ;
        RECT 185.525 13.515 185.695 13.685 ;
        RECT 185.985 13.515 186.155 13.685 ;
        RECT 186.445 13.515 186.615 13.685 ;
        RECT 186.905 13.515 187.075 13.685 ;
        RECT 187.365 13.515 187.535 13.685 ;
        RECT 188.285 13.515 188.455 13.685 ;
        RECT 191.045 13.515 191.215 13.685 ;
        RECT 194.265 13.515 194.435 13.685 ;
        RECT 194.725 13.515 194.895 13.685 ;
        RECT 195.185 13.515 195.355 13.685 ;
        RECT 195.645 13.515 195.815 13.685 ;
        RECT 196.105 13.515 196.275 13.685 ;
        RECT 196.565 13.515 196.735 13.685 ;
        RECT 197.025 13.515 197.195 13.685 ;
        RECT 197.485 13.515 197.655 13.685 ;
        RECT 197.945 13.515 198.115 13.685 ;
        RECT 198.405 13.515 198.575 13.685 ;
        RECT 198.865 13.515 199.035 13.685 ;
        RECT 199.325 13.515 199.495 13.685 ;
        RECT 199.785 13.515 199.955 13.685 ;
        RECT 200.245 13.515 200.415 13.685 ;
        RECT 200.705 13.515 200.875 13.685 ;
        RECT 201.165 13.515 201.335 13.685 ;
        RECT 201.625 13.515 201.795 13.685 ;
        RECT 202.085 13.515 202.255 13.685 ;
        RECT 205.305 13.515 205.475 13.685 ;
        RECT 205.765 13.515 205.935 13.685 ;
        RECT 206.225 13.515 206.395 13.685 ;
        RECT 206.685 13.515 206.855 13.685 ;
        RECT 207.145 13.515 207.315 13.685 ;
        RECT 207.605 13.515 207.775 13.685 ;
        RECT 208.065 13.515 208.235 13.685 ;
        RECT 208.525 13.515 208.695 13.685 ;
        RECT 208.985 13.515 209.155 13.685 ;
        RECT 209.445 13.515 209.615 13.685 ;
        RECT 209.905 13.515 210.075 13.685 ;
        RECT 210.365 13.515 210.535 13.685 ;
        RECT 210.825 13.515 210.995 13.685 ;
        RECT 211.285 13.515 211.455 13.685 ;
        RECT 211.745 13.515 211.915 13.685 ;
        RECT 212.205 13.515 212.375 13.685 ;
        RECT 212.665 13.515 212.835 13.685 ;
        RECT 213.125 13.515 213.295 13.685 ;
        RECT 213.585 13.515 213.755 13.685 ;
        RECT 214.045 13.515 214.215 13.685 ;
        RECT 214.505 13.515 214.675 13.685 ;
        RECT 214.965 13.515 215.135 13.685 ;
        RECT 215.425 13.515 215.595 13.685 ;
        RECT 216.345 13.515 216.515 13.685 ;
        RECT 218.185 13.515 218.355 13.685 ;
        RECT 218.645 13.515 218.815 13.685 ;
        RECT 219.105 13.515 219.275 13.685 ;
        RECT 219.565 13.515 219.735 13.685 ;
        RECT 220.025 13.515 220.195 13.685 ;
        RECT 220.485 13.515 220.655 13.685 ;
        RECT 220.945 13.515 221.115 13.685 ;
        RECT 221.405 13.515 221.575 13.685 ;
        RECT 221.865 13.515 222.035 13.685 ;
        RECT 222.325 13.515 222.495 13.685 ;
        RECT 222.785 13.515 222.955 13.685 ;
        RECT 223.245 13.515 223.415 13.685 ;
        RECT 223.705 13.515 223.875 13.685 ;
        RECT 224.165 13.515 224.335 13.685 ;
        RECT 225.545 13.515 225.715 13.685 ;
        RECT 226.005 13.515 226.175 13.685 ;
        RECT 226.465 13.515 226.635 13.685 ;
        RECT 226.925 13.515 227.095 13.685 ;
        RECT 227.385 13.515 227.555 13.685 ;
        RECT 227.845 13.515 228.015 13.685 ;
        RECT 228.305 13.515 228.475 13.685 ;
        RECT 228.765 13.515 228.935 13.685 ;
        RECT 229.225 13.515 229.395 13.685 ;
        RECT 229.685 13.515 229.855 13.685 ;
        RECT 230.145 13.515 230.315 13.685 ;
        RECT 230.605 13.515 230.775 13.685 ;
        RECT 231.065 13.515 231.235 13.685 ;
        RECT 231.525 13.515 231.695 13.685 ;
        RECT 231.985 13.515 232.155 13.685 ;
        RECT 232.445 13.515 232.615 13.685 ;
        RECT 232.905 13.515 233.075 13.685 ;
        RECT 233.365 13.515 233.535 13.685 ;
        RECT 233.825 13.515 233.995 13.685 ;
        RECT 234.285 13.515 234.455 13.685 ;
        RECT 234.745 13.515 234.915 13.685 ;
        RECT 235.205 13.515 235.375 13.685 ;
        RECT 235.665 13.515 235.835 13.685 ;
        RECT 236.125 13.515 236.295 13.685 ;
        RECT 237.045 13.515 237.215 13.685 ;
        RECT 237.505 13.515 237.675 13.685 ;
        RECT 237.965 13.515 238.135 13.685 ;
        RECT 238.425 13.515 238.595 13.685 ;
        RECT 238.885 13.515 239.055 13.685 ;
        RECT 239.345 13.515 239.515 13.685 ;
        RECT 239.805 13.515 239.975 13.685 ;
        RECT 240.265 13.515 240.435 13.685 ;
        RECT 240.725 13.515 240.895 13.685 ;
        RECT 241.185 13.515 241.355 13.685 ;
        RECT 241.645 13.515 241.815 13.685 ;
        RECT 242.105 13.515 242.275 13.685 ;
        RECT 242.565 13.515 242.735 13.685 ;
        RECT 243.025 13.515 243.195 13.685 ;
        RECT 243.485 13.515 243.655 13.685 ;
        RECT 243.945 13.515 244.115 13.685 ;
        RECT 244.405 13.515 244.575 13.685 ;
        RECT 248.085 13.515 248.255 13.685 ;
        RECT 259.125 13.515 259.295 13.685 ;
        RECT 259.585 13.515 259.755 13.685 ;
        RECT 260.045 13.515 260.215 13.685 ;
        RECT 260.505 13.515 260.675 13.685 ;
        RECT 260.965 13.515 261.135 13.685 ;
        RECT 261.425 13.515 261.595 13.685 ;
        RECT 261.885 13.515 262.055 13.685 ;
        RECT 262.345 13.515 262.515 13.685 ;
        RECT 262.805 13.515 262.975 13.685 ;
        RECT 263.265 13.515 263.435 13.685 ;
        RECT 263.725 13.515 263.895 13.685 ;
        RECT 264.185 13.515 264.355 13.685 ;
        RECT 264.645 13.515 264.815 13.685 ;
        RECT 265.105 13.515 265.275 13.685 ;
        RECT 265.565 13.515 265.735 13.685 ;
        RECT 266.025 13.515 266.195 13.685 ;
        RECT 266.485 13.515 266.655 13.685 ;
        RECT 266.945 13.515 267.115 13.685 ;
        RECT 267.405 13.515 267.575 13.685 ;
        RECT 267.865 13.515 268.035 13.685 ;
        RECT 268.325 13.515 268.495 13.685 ;
        RECT 268.785 13.515 268.955 13.685 ;
        RECT 269.245 13.515 269.415 13.685 ;
        RECT 272.465 13.515 272.635 13.685 ;
        RECT 276.605 13.515 276.775 13.685 ;
        RECT 277.525 13.515 277.695 13.685 ;
        RECT 277.985 13.515 278.155 13.685 ;
        RECT 278.445 13.515 278.615 13.685 ;
        RECT 283.045 13.515 283.215 13.685 ;
        RECT 283.505 13.515 283.675 13.685 ;
        RECT 283.965 13.515 284.135 13.685 ;
        RECT 284.425 13.515 284.595 13.685 ;
        RECT 289.025 13.515 289.195 13.685 ;
        RECT 289.485 13.515 289.655 13.685 ;
        RECT 289.945 13.515 290.115 13.685 ;
        RECT 290.865 13.515 291.035 13.685 ;
        RECT 292.705 13.515 292.875 13.685 ;
        RECT 293.165 13.515 293.335 13.685 ;
        RECT 293.625 13.515 293.795 13.685 ;
        RECT 294.085 13.515 294.255 13.685 ;
        RECT 294.545 13.515 294.715 13.685 ;
        RECT 295.005 13.515 295.175 13.685 ;
        RECT 295.465 13.515 295.635 13.685 ;
        RECT 295.925 13.515 296.095 13.685 ;
        RECT 296.385 13.515 296.555 13.685 ;
        RECT 296.845 13.515 297.015 13.685 ;
        RECT 297.305 13.515 297.475 13.685 ;
        RECT 297.765 13.515 297.935 13.685 ;
        RECT 298.225 13.515 298.395 13.685 ;
        RECT 298.685 13.515 298.855 13.685 ;
        RECT 300.525 13.515 300.695 13.685 ;
        RECT 304.665 13.515 304.835 13.685 ;
        RECT 305.125 13.515 305.295 13.685 ;
        RECT 305.585 13.515 305.755 13.685 ;
        RECT 306.045 13.515 306.215 13.685 ;
        RECT 306.505 13.515 306.675 13.685 ;
        RECT 306.965 13.515 307.135 13.685 ;
        RECT 307.885 13.515 308.055 13.685 ;
        RECT 308.345 13.515 308.515 13.685 ;
        RECT 308.805 13.515 308.975 13.685 ;
        RECT 309.265 13.515 309.435 13.685 ;
        RECT 309.725 13.515 309.895 13.685 ;
        RECT 310.185 13.515 310.355 13.685 ;
        RECT 310.645 13.515 310.815 13.685 ;
        RECT 311.105 13.515 311.275 13.685 ;
        RECT 314.325 13.515 314.495 13.685 ;
        RECT 314.785 13.515 314.955 13.685 ;
        RECT 315.245 13.515 315.415 13.685 ;
        RECT 317.545 13.515 317.715 13.685 ;
        RECT 318.005 13.515 318.175 13.685 ;
        RECT 318.465 13.515 318.635 13.685 ;
        RECT 318.925 13.515 319.095 13.685 ;
        RECT 319.385 13.515 319.555 13.685 ;
        RECT 319.845 13.515 320.015 13.685 ;
        RECT 320.305 13.515 320.475 13.685 ;
        RECT 320.765 13.515 320.935 13.685 ;
        RECT 321.225 13.515 321.395 13.685 ;
        RECT 321.685 13.515 321.855 13.685 ;
        RECT 322.145 13.515 322.315 13.685 ;
        RECT 322.605 13.515 322.775 13.685 ;
        RECT 323.065 13.515 323.235 13.685 ;
        RECT 323.525 13.515 323.695 13.685 ;
        RECT 323.985 13.515 324.155 13.685 ;
        RECT 324.445 13.515 324.615 13.685 ;
        RECT 324.905 13.515 325.075 13.685 ;
        RECT 325.365 13.515 325.535 13.685 ;
        RECT 325.825 13.515 325.995 13.685 ;
        RECT 328.585 13.515 328.755 13.685 ;
        RECT 329.045 13.515 329.215 13.685 ;
        RECT 329.505 13.515 329.675 13.685 ;
        RECT 329.965 13.515 330.135 13.685 ;
        RECT 330.425 13.515 330.595 13.685 ;
        RECT 330.885 13.515 331.055 13.685 ;
        RECT 331.345 13.515 331.515 13.685 ;
        RECT 331.805 13.515 331.975 13.685 ;
        RECT 332.265 13.515 332.435 13.685 ;
        RECT 332.725 13.515 332.895 13.685 ;
        RECT 333.185 13.515 333.355 13.685 ;
        RECT 333.645 13.515 333.815 13.685 ;
        RECT 334.105 13.515 334.275 13.685 ;
        RECT 334.565 13.515 334.735 13.685 ;
        RECT 335.025 13.515 335.195 13.685 ;
        RECT 335.485 13.515 335.655 13.685 ;
        RECT 335.945 13.515 336.115 13.685 ;
        RECT 336.405 13.515 336.575 13.685 ;
        RECT 336.865 13.515 337.035 13.685 ;
        RECT 337.325 13.515 337.495 13.685 ;
        RECT 339.165 13.515 339.335 13.685 ;
        RECT 339.625 13.515 339.795 13.685 ;
        RECT 340.085 13.515 340.255 13.685 ;
        RECT 340.545 13.515 340.715 13.685 ;
        RECT 347.905 13.515 348.075 13.685 ;
        RECT 348.365 13.515 348.535 13.685 ;
        RECT 348.825 13.515 348.995 13.685 ;
        RECT 349.285 13.515 349.455 13.685 ;
        RECT 349.745 13.515 349.915 13.685 ;
        RECT 350.205 13.515 350.375 13.685 ;
        RECT 350.665 13.515 350.835 13.685 ;
        RECT 351.125 13.515 351.295 13.685 ;
        RECT 351.585 13.515 351.755 13.685 ;
        RECT 352.045 13.515 352.215 13.685 ;
        RECT 352.505 13.515 352.675 13.685 ;
        RECT 352.965 13.515 353.135 13.685 ;
        RECT 353.425 13.515 353.595 13.685 ;
        RECT 353.885 13.515 354.055 13.685 ;
        RECT 354.345 13.515 354.515 13.685 ;
        RECT 354.805 13.515 354.975 13.685 ;
        RECT 355.265 13.515 355.435 13.685 ;
        RECT 355.725 13.515 355.895 13.685 ;
        RECT 356.185 13.515 356.355 13.685 ;
        RECT 356.645 13.515 356.815 13.685 ;
        RECT 357.105 13.515 357.275 13.685 ;
        RECT 357.565 13.515 357.735 13.685 ;
        RECT 358.025 13.515 358.195 13.685 ;
        RECT 358.485 13.515 358.655 13.685 ;
        RECT 359.865 13.515 360.035 13.685 ;
        RECT 360.325 13.515 360.495 13.685 ;
        RECT 360.785 13.515 360.955 13.685 ;
        RECT 361.245 13.515 361.415 13.685 ;
        RECT 361.705 13.515 361.875 13.685 ;
        RECT 362.165 13.515 362.335 13.685 ;
        RECT 362.625 13.515 362.795 13.685 ;
        RECT 363.085 13.515 363.255 13.685 ;
        RECT 363.545 13.515 363.715 13.685 ;
        RECT 364.005 13.515 364.175 13.685 ;
        RECT 364.465 13.515 364.635 13.685 ;
        RECT 364.925 13.515 365.095 13.685 ;
        RECT 365.385 13.515 365.555 13.685 ;
        RECT 365.845 13.515 366.015 13.685 ;
        RECT 366.305 13.515 366.475 13.685 ;
        RECT 366.765 13.515 366.935 13.685 ;
        RECT 368.145 13.515 368.315 13.685 ;
        RECT 368.605 13.515 368.775 13.685 ;
        RECT 369.065 13.515 369.235 13.685 ;
        RECT 369.525 13.515 369.695 13.685 ;
        RECT 369.985 13.515 370.155 13.685 ;
        RECT 370.445 13.515 370.615 13.685 ;
        RECT 370.905 13.515 371.075 13.685 ;
        RECT 371.365 13.515 371.535 13.685 ;
        RECT 371.825 13.515 371.995 13.685 ;
        RECT 372.285 13.515 372.455 13.685 ;
        RECT 372.745 13.515 372.915 13.685 ;
        RECT 373.205 13.515 373.375 13.685 ;
        RECT 373.665 13.515 373.835 13.685 ;
        RECT 374.125 13.515 374.295 13.685 ;
        RECT 374.585 13.515 374.755 13.685 ;
        RECT 375.045 13.515 375.215 13.685 ;
        RECT 376.425 13.515 376.595 13.685 ;
        RECT 384.705 13.515 384.875 13.685 ;
        RECT 385.165 13.515 385.335 13.685 ;
        RECT 385.625 13.515 385.795 13.685 ;
        RECT 386.085 13.515 386.255 13.685 ;
        RECT 386.545 13.515 386.715 13.685 ;
        RECT 387.005 13.515 387.175 13.685 ;
        RECT 387.465 13.515 387.635 13.685 ;
        RECT 387.925 13.515 388.095 13.685 ;
        RECT 388.385 13.515 388.555 13.685 ;
        RECT 388.845 13.515 389.015 13.685 ;
        RECT 389.305 13.515 389.475 13.685 ;
        RECT 389.765 13.515 389.935 13.685 ;
        RECT 390.225 13.515 390.395 13.685 ;
        RECT 390.685 13.515 390.855 13.685 ;
        RECT 391.145 13.515 391.315 13.685 ;
        RECT 391.605 13.515 391.775 13.685 ;
        RECT 392.065 13.515 392.235 13.685 ;
        RECT 392.525 13.515 392.695 13.685 ;
        RECT 392.985 13.515 393.155 13.685 ;
        RECT 393.445 13.515 393.615 13.685 ;
        RECT 393.905 13.515 394.075 13.685 ;
        RECT 394.365 13.515 394.535 13.685 ;
        RECT 394.825 13.515 394.995 13.685 ;
        RECT 395.285 13.515 395.455 13.685 ;
        RECT 395.745 13.515 395.915 13.685 ;
        RECT 396.205 13.515 396.375 13.685 ;
        RECT 396.665 13.515 396.835 13.685 ;
        RECT 397.125 13.515 397.295 13.685 ;
        RECT 397.585 13.515 397.755 13.685 ;
        RECT 398.045 13.515 398.215 13.685 ;
        RECT 398.505 13.515 398.675 13.685 ;
        RECT 398.965 13.515 399.135 13.685 ;
        RECT 399.425 13.515 399.595 13.685 ;
        RECT 399.885 13.515 400.055 13.685 ;
        RECT 400.345 13.515 400.515 13.685 ;
        RECT 400.805 13.515 400.975 13.685 ;
        RECT 401.265 13.515 401.435 13.685 ;
        RECT 401.725 13.515 401.895 13.685 ;
        RECT 402.185 13.515 402.355 13.685 ;
        RECT 402.645 13.515 402.815 13.685 ;
        RECT 403.105 13.515 403.275 13.685 ;
        RECT 403.565 13.515 403.735 13.685 ;
        RECT 404.025 13.515 404.195 13.685 ;
        RECT 404.945 13.515 405.115 13.685 ;
        RECT 412.765 13.515 412.935 13.685 ;
        RECT 413.685 13.515 413.855 13.685 ;
        RECT 414.145 13.515 414.315 13.685 ;
        RECT 414.605 13.515 414.775 13.685 ;
        RECT 415.065 13.515 415.235 13.685 ;
        RECT 415.525 13.515 415.695 13.685 ;
        RECT 415.985 13.515 416.155 13.685 ;
        RECT 416.445 13.515 416.615 13.685 ;
        RECT 416.905 13.515 417.075 13.685 ;
        RECT 417.365 13.515 417.535 13.685 ;
        RECT 417.825 13.515 417.995 13.685 ;
        RECT 418.285 13.515 418.455 13.685 ;
        RECT 418.745 13.515 418.915 13.685 ;
        RECT 419.205 13.515 419.375 13.685 ;
        RECT 419.665 13.515 419.835 13.685 ;
        RECT 420.125 13.515 420.295 13.685 ;
        RECT 420.585 13.515 420.755 13.685 ;
        RECT 425.645 13.515 425.815 13.685 ;
        RECT 426.105 13.515 426.275 13.685 ;
        RECT 426.565 13.515 426.735 13.685 ;
        RECT 427.025 13.515 427.195 13.685 ;
        RECT 427.485 13.515 427.655 13.685 ;
        RECT 427.945 13.515 428.115 13.685 ;
        RECT 428.405 13.515 428.575 13.685 ;
        RECT 428.865 13.515 429.035 13.685 ;
        RECT 429.325 13.515 429.495 13.685 ;
        RECT 429.785 13.515 429.955 13.685 ;
        RECT 430.245 13.515 430.415 13.685 ;
        RECT 430.705 13.515 430.875 13.685 ;
        RECT 431.165 13.515 431.335 13.685 ;
        RECT 431.625 13.515 431.795 13.685 ;
        RECT 432.085 13.515 432.255 13.685 ;
        RECT 432.545 13.515 432.715 13.685 ;
        RECT 433.005 13.515 433.175 13.685 ;
        RECT 433.465 13.515 433.635 13.685 ;
        RECT 433.925 13.515 434.095 13.685 ;
        RECT 440.825 13.515 440.995 13.685 ;
        RECT 445.425 13.515 445.595 13.685 ;
        RECT 445.885 13.515 446.055 13.685 ;
        RECT 446.345 13.515 446.515 13.685 ;
        RECT 446.805 13.515 446.975 13.685 ;
        RECT 447.265 13.515 447.435 13.685 ;
        RECT 447.725 13.515 447.895 13.685 ;
        RECT 448.185 13.515 448.355 13.685 ;
        RECT 448.645 13.515 448.815 13.685 ;
        RECT 449.105 13.515 449.275 13.685 ;
        RECT 449.565 13.515 449.735 13.685 ;
        RECT 450.025 13.515 450.195 13.685 ;
        RECT 450.485 13.515 450.655 13.685 ;
        RECT 450.945 13.515 451.115 13.685 ;
        RECT 451.405 13.515 451.575 13.685 ;
        RECT 451.865 13.515 452.035 13.685 ;
        RECT 452.325 13.515 452.495 13.685 ;
        RECT 452.785 13.515 452.955 13.685 ;
        RECT 453.245 13.515 453.415 13.685 ;
        RECT 453.705 13.515 453.875 13.685 ;
        RECT 454.165 13.515 454.335 13.685 ;
        RECT 454.625 13.515 454.795 13.685 ;
        RECT 455.085 13.515 455.255 13.685 ;
        RECT 455.545 13.515 455.715 13.685 ;
        RECT 456.005 13.515 456.175 13.685 ;
        RECT 456.465 13.515 456.635 13.685 ;
        RECT 456.925 13.515 457.095 13.685 ;
        RECT 457.845 13.515 458.015 13.685 ;
        RECT 458.305 13.515 458.475 13.685 ;
        RECT 458.765 13.515 458.935 13.685 ;
        RECT 459.225 13.515 459.395 13.685 ;
        RECT 459.685 13.515 459.855 13.685 ;
        RECT 460.145 13.515 460.315 13.685 ;
        RECT 460.605 13.515 460.775 13.685 ;
        RECT 461.065 13.515 461.235 13.685 ;
        RECT 461.525 13.515 461.695 13.685 ;
        RECT 461.985 13.515 462.155 13.685 ;
        RECT 462.445 13.515 462.615 13.685 ;
        RECT 462.905 13.515 463.075 13.685 ;
        RECT 463.365 13.515 463.535 13.685 ;
        RECT 463.825 13.515 463.995 13.685 ;
        RECT 464.285 13.515 464.455 13.685 ;
        RECT 464.745 13.515 464.915 13.685 ;
        RECT 465.205 13.515 465.375 13.685 ;
        RECT 465.665 13.515 465.835 13.685 ;
        RECT 466.125 13.515 466.295 13.685 ;
        RECT 467.045 13.515 467.215 13.685 ;
        RECT 467.505 13.515 467.675 13.685 ;
        RECT 467.965 13.515 468.135 13.685 ;
        RECT 468.425 13.515 468.595 13.685 ;
        RECT 468.885 13.515 469.055 13.685 ;
        RECT 476.245 13.515 476.415 13.685 ;
        RECT 480.845 13.515 481.015 13.685 ;
        RECT 481.305 13.515 481.475 13.685 ;
        RECT 481.765 13.515 481.935 13.685 ;
        RECT 482.225 13.515 482.395 13.685 ;
        RECT 490.505 13.515 490.675 13.685 ;
        RECT 494.645 13.515 494.815 13.685 ;
        RECT 495.105 13.515 495.275 13.685 ;
        RECT 495.565 13.515 495.735 13.685 ;
        RECT 496.945 13.515 497.115 13.685 ;
        RECT 504.765 13.515 504.935 13.685 ;
        RECT 519.025 13.515 519.195 13.685 ;
        RECT 525.005 13.515 525.175 13.685 ;
        RECT 527.765 13.515 527.935 13.685 ;
        RECT 528.225 13.515 528.395 13.685 ;
        RECT 528.685 13.515 528.855 13.685 ;
        RECT 529.145 13.515 529.315 13.685 ;
        RECT 529.605 13.515 529.775 13.685 ;
        RECT 530.065 13.515 530.235 13.685 ;
        RECT 530.525 13.515 530.695 13.685 ;
        RECT 530.985 13.515 531.155 13.685 ;
        RECT 531.445 13.515 531.615 13.685 ;
        RECT 531.905 13.515 532.075 13.685 ;
        RECT 532.365 13.515 532.535 13.685 ;
        RECT 532.825 13.515 532.995 13.685 ;
        RECT 533.285 13.515 533.455 13.685 ;
        RECT 533.745 13.515 533.915 13.685 ;
        RECT 536.045 13.515 536.215 13.685 ;
        RECT 536.505 13.515 536.675 13.685 ;
        RECT 536.965 13.515 537.135 13.685 ;
        RECT 538.805 13.515 538.975 13.685 ;
        RECT 539.265 13.515 539.435 13.685 ;
        RECT 539.725 13.515 539.895 13.685 ;
        RECT 540.185 13.515 540.355 13.685 ;
        RECT 547.545 13.515 547.715 13.685 ;
        RECT 553.065 13.515 553.235 13.685 ;
        RECT 561.805 13.515 561.975 13.685 ;
        RECT 564.105 13.515 564.275 13.685 ;
        RECT 564.565 13.515 564.735 13.685 ;
        RECT 565.025 13.515 565.195 13.685 ;
        RECT 565.485 13.515 565.655 13.685 ;
        RECT 571.005 13.515 571.175 13.685 ;
        RECT 571.465 13.515 571.635 13.685 ;
        RECT 571.925 13.515 572.095 13.685 ;
        RECT 572.385 13.515 572.555 13.685 ;
        RECT 572.845 13.515 573.015 13.685 ;
        RECT 573.305 13.515 573.475 13.685 ;
        RECT 573.765 13.515 573.935 13.685 ;
        RECT 574.225 13.515 574.395 13.685 ;
        RECT 574.685 13.515 574.855 13.685 ;
        RECT 575.145 13.515 575.315 13.685 ;
        RECT 575.605 13.515 575.775 13.685 ;
        RECT 576.065 13.515 576.235 13.685 ;
        RECT 576.525 13.515 576.695 13.685 ;
        RECT 576.985 13.515 577.155 13.685 ;
        RECT 577.445 13.515 577.615 13.685 ;
        RECT 577.905 13.515 578.075 13.685 ;
        RECT 578.365 13.515 578.535 13.685 ;
        RECT 578.825 13.515 578.995 13.685 ;
        RECT 579.285 13.515 579.455 13.685 ;
        RECT 579.745 13.515 579.915 13.685 ;
        RECT 580.205 13.515 580.375 13.685 ;
        RECT 581.125 13.515 581.295 13.685 ;
        RECT 590.325 13.515 590.495 13.685 ;
        RECT 604.585 13.515 604.755 13.685 ;
        RECT 609.185 13.515 609.355 13.685 ;
        RECT 618.845 13.515 619.015 13.685 ;
        RECT 633.105 13.515 633.275 13.685 ;
        RECT 637.245 13.515 637.415 13.685 ;
        RECT 647.365 13.515 647.535 13.685 ;
        RECT 661.625 13.515 661.795 13.685 ;
        RECT 665.305 13.515 665.475 13.685 ;
        RECT 675.885 13.515 676.055 13.685 ;
        RECT 690.145 13.515 690.315 13.685 ;
        RECT 693.365 13.515 693.535 13.685 ;
        RECT 704.405 13.515 704.575 13.685 ;
        RECT 718.665 13.515 718.835 13.685 ;
        RECT 721.425 13.515 721.595 13.685 ;
        RECT 732.925 13.515 733.095 13.685 ;
        RECT 747.185 13.515 747.355 13.685 ;
        RECT 749.485 13.515 749.655 13.685 ;
        RECT 761.445 13.515 761.615 13.685 ;
        RECT 775.705 13.515 775.875 13.685 ;
        RECT 777.545 13.515 777.715 13.685 ;
        RECT 789.965 13.515 790.135 13.685 ;
        RECT 804.225 13.515 804.395 13.685 ;
        RECT 805.605 13.515 805.775 13.685 ;
        RECT 818.485 13.515 818.655 13.685 ;
        RECT 832.745 13.515 832.915 13.685 ;
        RECT 833.665 13.515 833.835 13.685 ;
        RECT 847.005 13.515 847.175 13.685 ;
        RECT 861.265 13.515 861.435 13.685 ;
        RECT 861.725 13.515 861.895 13.685 ;
        RECT 875.525 13.515 875.695 13.685 ;
        RECT 889.785 13.515 889.955 13.685 ;
        RECT 904.045 13.515 904.215 13.685 ;
        RECT 917.845 13.515 918.015 13.685 ;
        RECT 918.305 13.515 918.475 13.685 ;
        RECT 932.565 13.515 932.735 13.685 ;
        RECT 945.905 13.515 946.075 13.685 ;
        RECT 946.825 13.515 946.995 13.685 ;
        RECT 961.085 13.515 961.255 13.685 ;
        RECT 973.965 13.515 974.135 13.685 ;
        RECT 975.345 13.515 975.515 13.685 ;
        RECT 989.605 13.515 989.775 13.685 ;
        RECT 1002.025 13.515 1002.195 13.685 ;
        RECT 1003.865 13.515 1004.035 13.685 ;
        RECT 1018.125 13.515 1018.295 13.685 ;
        RECT 1030.085 13.515 1030.255 13.685 ;
        RECT 1032.385 13.515 1032.555 13.685 ;
        RECT 1046.645 13.515 1046.815 13.685 ;
        RECT 1058.145 13.515 1058.315 13.685 ;
        RECT 1060.905 13.515 1061.075 13.685 ;
        RECT 1075.165 13.515 1075.335 13.685 ;
        RECT 1086.205 13.515 1086.375 13.685 ;
        RECT 1089.425 13.515 1089.595 13.685 ;
        RECT 1103.685 13.515 1103.855 13.685 ;
        RECT 1114.265 13.515 1114.435 13.685 ;
        RECT 1117.945 13.515 1118.115 13.685 ;
        RECT 1132.205 13.515 1132.375 13.685 ;
        RECT 1142.325 13.515 1142.495 13.685 ;
        RECT 1146.465 13.515 1146.635 13.685 ;
        RECT 1160.725 13.515 1160.895 13.685 ;
        RECT 1170.385 13.515 1170.555 13.685 ;
        RECT 1174.985 13.515 1175.155 13.685 ;
        RECT 1189.245 13.515 1189.415 13.685 ;
        RECT 1198.445 13.515 1198.615 13.685 ;
        RECT 1203.505 13.515 1203.675 13.685 ;
        RECT 1217.765 13.515 1217.935 13.685 ;
        RECT 1226.505 13.515 1226.675 13.685 ;
        RECT 1232.025 13.515 1232.195 13.685 ;
        RECT 1246.285 13.515 1246.455 13.685 ;
        RECT 1254.565 13.515 1254.735 13.685 ;
        RECT 1260.545 13.515 1260.715 13.685 ;
        RECT 1274.805 13.515 1274.975 13.685 ;
        RECT 1282.625 13.515 1282.795 13.685 ;
        RECT 1289.065 13.515 1289.235 13.685 ;
        RECT 1303.325 13.515 1303.495 13.685 ;
        RECT 1310.685 13.515 1310.855 13.685 ;
        RECT 1317.585 13.515 1317.755 13.685 ;
        RECT 1331.845 13.515 1332.015 13.685 ;
        RECT 1338.745 13.515 1338.915 13.685 ;
        RECT 1346.105 13.515 1346.275 13.685 ;
        RECT 1360.365 13.515 1360.535 13.685 ;
        RECT 1366.805 13.515 1366.975 13.685 ;
        RECT 1374.625 13.515 1374.795 13.685 ;
        RECT 1382.445 13.515 1382.615 13.685 ;
        RECT 1382.905 13.515 1383.075 13.685 ;
        RECT 1383.365 13.515 1383.535 13.685 ;
        RECT 1388.885 13.515 1389.055 13.685 ;
        RECT 1394.865 13.515 1395.035 13.685 ;
        RECT 1400.845 13.515 1401.015 13.685 ;
        RECT 1401.305 13.515 1401.475 13.685 ;
        RECT 1401.765 13.515 1401.935 13.685 ;
        RECT 1403.145 13.515 1403.315 13.685 ;
        RECT 1417.405 13.515 1417.575 13.685 ;
        RECT 1422.925 13.515 1423.095 13.685 ;
        RECT 1431.665 13.515 1431.835 13.685 ;
        RECT 1445.925 13.515 1446.095 13.685 ;
        RECT 1450.985 13.515 1451.155 13.685 ;
        RECT 1460.185 13.515 1460.355 13.685 ;
        RECT 1474.445 13.515 1474.615 13.685 ;
        RECT 1479.045 13.515 1479.215 13.685 ;
        RECT 1488.705 13.515 1488.875 13.685 ;
        RECT 1502.965 13.515 1503.135 13.685 ;
        RECT 1503.885 13.515 1504.055 13.685 ;
        RECT 1504.345 13.515 1504.515 13.685 ;
        RECT 1504.805 13.515 1504.975 13.685 ;
        RECT 1507.105 13.515 1507.275 13.685 ;
        RECT 1517.225 13.515 1517.395 13.685 ;
        RECT 1525.965 13.515 1526.135 13.685 ;
        RECT 1526.425 13.515 1526.595 13.685 ;
        RECT 1526.885 13.515 1527.055 13.685 ;
        RECT 1531.485 13.515 1531.655 13.685 ;
        RECT 1535.165 13.515 1535.335 13.685 ;
        RECT 1535.625 13.515 1535.795 13.685 ;
        RECT 1536.085 13.515 1536.255 13.685 ;
        RECT 1536.545 13.515 1536.715 13.685 ;
        RECT 1539.305 13.515 1539.475 13.685 ;
        RECT 1539.765 13.515 1539.935 13.685 ;
        RECT 1540.225 13.515 1540.395 13.685 ;
        RECT 1542.525 13.515 1542.695 13.685 ;
        RECT 1542.985 13.515 1543.155 13.685 ;
        RECT 1543.445 13.515 1543.615 13.685 ;
        RECT 1545.745 13.515 1545.915 13.685 ;
        RECT 1559.085 13.515 1559.255 13.685 ;
        RECT 1559.545 13.515 1559.715 13.685 ;
        RECT 1560.005 13.515 1560.175 13.685 ;
        RECT 1563.225 13.515 1563.395 13.685 ;
        RECT 1574.265 13.515 1574.435 13.685 ;
        RECT 1575.645 13.515 1575.815 13.685 ;
        RECT 1576.105 13.515 1576.275 13.685 ;
        RECT 1576.565 13.515 1576.735 13.685 ;
        RECT 1588.525 13.515 1588.695 13.685 ;
        RECT 1588.985 13.515 1589.155 13.685 ;
        RECT 1589.445 13.515 1589.615 13.685 ;
        RECT 1591.285 13.515 1591.455 13.685 ;
        RECT 1602.785 13.515 1602.955 13.685 ;
        RECT 1617.045 13.515 1617.215 13.685 ;
        RECT 1619.345 13.515 1619.515 13.685 ;
        RECT 1625.785 13.515 1625.955 13.685 ;
        RECT 1626.245 13.515 1626.415 13.685 ;
        RECT 1626.705 13.515 1626.875 13.685 ;
        RECT 1631.305 13.515 1631.475 13.685 ;
        RECT 1645.565 13.515 1645.735 13.685 ;
        RECT 1647.405 13.515 1647.575 13.685 ;
        RECT 1648.785 13.515 1648.955 13.685 ;
        RECT 1649.245 13.515 1649.415 13.685 ;
        RECT 1649.705 13.515 1649.875 13.685 ;
        RECT 1659.825 13.515 1659.995 13.685 ;
        RECT 1674.085 13.515 1674.255 13.685 ;
        RECT 1675.465 13.515 1675.635 13.685 ;
        RECT 1688.345 13.515 1688.515 13.685 ;
        RECT 1702.605 13.515 1702.775 13.685 ;
        RECT 1703.525 13.515 1703.695 13.685 ;
        RECT 1716.865 13.515 1717.035 13.685 ;
        RECT 1731.125 13.515 1731.295 13.685 ;
        RECT 1731.585 13.515 1731.755 13.685 ;
        RECT 1745.385 13.515 1745.555 13.685 ;
        RECT 1759.645 13.515 1759.815 13.685 ;
        RECT 1760.105 13.515 1760.275 13.685 ;
        RECT 1760.565 13.515 1760.735 13.685 ;
        RECT 1761.025 13.515 1761.195 13.685 ;
        RECT 1773.905 13.515 1774.075 13.685 ;
        RECT 1774.365 13.515 1774.535 13.685 ;
        RECT 1774.825 13.515 1774.995 13.685 ;
        RECT 1787.705 13.515 1787.875 13.685 ;
        RECT 1788.165 13.515 1788.335 13.685 ;
        RECT 1802.425 13.515 1802.595 13.685 ;
        RECT 1815.765 13.515 1815.935 13.685 ;
        RECT 1816.685 13.515 1816.855 13.685 ;
        RECT 1830.025 13.515 1830.195 13.685 ;
        RECT 1830.485 13.515 1830.655 13.685 ;
        RECT 1830.945 13.515 1831.115 13.685 ;
        RECT 1843.825 13.515 1843.995 13.685 ;
        RECT 1845.205 13.515 1845.375 13.685 ;
        RECT 1859.465 13.515 1859.635 13.685 ;
        RECT 1871.885 13.515 1872.055 13.685 ;
        RECT 1873.725 13.515 1873.895 13.685 ;
        RECT 1887.985 13.515 1888.155 13.685 ;
        RECT 1899.945 13.515 1900.115 13.685 ;
        RECT 1902.245 13.515 1902.415 13.685 ;
        RECT 1913.285 13.515 1913.455 13.685 ;
        RECT 1913.745 13.515 1913.915 13.685 ;
        RECT 1914.205 13.515 1914.375 13.685 ;
        RECT 1916.505 13.515 1916.675 13.685 ;
        RECT 1925.705 13.515 1925.875 13.685 ;
        RECT 1926.165 13.515 1926.335 13.685 ;
        RECT 1926.625 13.515 1926.795 13.685 ;
        RECT 1928.005 13.515 1928.175 13.685 ;
        RECT 1930.765 13.515 1930.935 13.685 ;
        RECT 1931.685 13.515 1931.855 13.685 ;
        RECT 1932.145 13.515 1932.315 13.685 ;
        RECT 1932.605 13.515 1932.775 13.685 ;
        RECT 1945.025 13.515 1945.195 13.685 ;
        RECT 1947.785 13.515 1947.955 13.685 ;
        RECT 1948.245 13.515 1948.415 13.685 ;
        RECT 1948.705 13.515 1948.875 13.685 ;
        RECT 1956.065 13.515 1956.235 13.685 ;
        RECT 1959.285 13.515 1959.455 13.685 ;
        RECT 1973.085 13.515 1973.255 13.685 ;
        RECT 1973.545 13.515 1973.715 13.685 ;
        RECT 1974.005 13.515 1974.175 13.685 ;
        RECT 1982.745 13.515 1982.915 13.685 ;
        RECT 1983.205 13.515 1983.375 13.685 ;
        RECT 1983.665 13.515 1983.835 13.685 ;
        RECT 1984.125 13.515 1984.295 13.685 ;
        RECT 1987.805 13.515 1987.975 13.685 ;
        RECT 1991.945 13.515 1992.115 13.685 ;
        RECT 1992.405 13.515 1992.575 13.685 ;
        RECT 1992.865 13.515 1993.035 13.685 ;
        RECT 1995.165 13.515 1995.335 13.685 ;
        RECT 1995.625 13.515 1995.795 13.685 ;
        RECT 1996.085 13.515 1996.255 13.685 ;
        RECT 1999.765 13.515 1999.935 13.685 ;
        RECT 2000.225 13.515 2000.395 13.685 ;
        RECT 2000.685 13.515 2000.855 13.685 ;
        RECT 2002.065 13.515 2002.235 13.685 ;
        RECT 2012.185 13.515 2012.355 13.685 ;
        RECT 2016.325 13.515 2016.495 13.685 ;
        RECT 2018.165 13.515 2018.335 13.685 ;
        RECT 2018.625 13.515 2018.795 13.685 ;
        RECT 2019.085 13.515 2019.255 13.685 ;
        RECT 2024.605 13.515 2024.775 13.685 ;
        RECT 2025.065 13.515 2025.235 13.685 ;
        RECT 2025.525 13.515 2025.695 13.685 ;
        RECT 2030.585 13.515 2030.755 13.685 ;
        RECT 2037.485 13.515 2037.655 13.685 ;
        RECT 2037.945 13.515 2038.115 13.685 ;
        RECT 2038.405 13.515 2038.575 13.685 ;
        RECT 2040.245 13.515 2040.415 13.685 ;
        RECT 2044.845 13.515 2045.015 13.685 ;
        RECT 2059.105 13.515 2059.275 13.685 ;
        RECT 2059.565 13.515 2059.735 13.685 ;
        RECT 2060.025 13.515 2060.195 13.685 ;
        RECT 2060.485 13.515 2060.655 13.685 ;
        RECT 2060.945 13.515 2061.115 13.685 ;
        RECT 2061.405 13.515 2061.575 13.685 ;
        RECT 2068.305 13.515 2068.475 13.685 ;
        RECT 2073.365 13.515 2073.535 13.685 ;
        RECT 2073.825 13.515 2073.995 13.685 ;
        RECT 2074.285 13.515 2074.455 13.685 ;
        RECT 2074.745 13.515 2074.915 13.685 ;
        RECT 2087.625 13.515 2087.795 13.685 ;
        RECT 2089.925 13.515 2090.095 13.685 ;
        RECT 2090.385 13.515 2090.555 13.685 ;
        RECT 2090.845 13.515 2091.015 13.685 ;
        RECT 2096.365 13.515 2096.535 13.685 ;
        RECT 2101.885 13.515 2102.055 13.685 ;
        RECT 2105.105 13.515 2105.275 13.685 ;
        RECT 2105.565 13.515 2105.735 13.685 ;
        RECT 2106.025 13.515 2106.195 13.685 ;
        RECT 2116.145 13.515 2116.315 13.685 ;
        RECT 2124.425 13.515 2124.595 13.685 ;
        RECT 2124.885 13.515 2125.055 13.685 ;
        RECT 2125.345 13.515 2125.515 13.685 ;
        RECT 2125.805 13.515 2125.975 13.685 ;
        RECT 2130.405 13.515 2130.575 13.685 ;
        RECT 2135.465 13.515 2135.635 13.685 ;
        RECT 2135.925 13.515 2136.095 13.685 ;
        RECT 2136.385 13.515 2136.555 13.685 ;
        RECT 2136.845 13.515 2137.015 13.685 ;
        RECT 2137.305 13.515 2137.475 13.685 ;
        RECT 2137.765 13.515 2137.935 13.685 ;
        RECT 2140.985 13.515 2141.155 13.685 ;
        RECT 2141.445 13.515 2141.615 13.685 ;
        RECT 2141.905 13.515 2142.075 13.685 ;
        RECT 2144.665 13.515 2144.835 13.685 ;
        RECT 2152.485 13.515 2152.655 13.685 ;
        RECT 2158.925 13.515 2159.095 13.685 ;
        RECT 2173.185 13.515 2173.355 13.685 ;
        RECT 2174.105 13.515 2174.275 13.685 ;
        RECT 2174.565 13.515 2174.735 13.685 ;
        RECT 2175.025 13.515 2175.195 13.685 ;
        RECT 2179.165 13.515 2179.335 13.685 ;
        RECT 2179.625 13.515 2179.795 13.685 ;
        RECT 2180.085 13.515 2180.255 13.685 ;
        RECT 2180.545 13.515 2180.715 13.685 ;
        RECT 2187.445 13.515 2187.615 13.685 ;
        RECT 2189.745 13.515 2189.915 13.685 ;
        RECT 2190.205 13.515 2190.375 13.685 ;
        RECT 2190.665 13.515 2190.835 13.685 ;
        RECT 2192.045 13.515 2192.215 13.685 ;
        RECT 2192.505 13.515 2192.675 13.685 ;
        RECT 2192.965 13.515 2193.135 13.685 ;
        RECT 2201.705 13.515 2201.875 13.685 ;
        RECT 2208.605 13.515 2208.775 13.685 ;
        RECT 2215.965 13.515 2216.135 13.685 ;
        RECT 2230.225 13.515 2230.395 13.685 ;
        RECT 2233.905 13.515 2234.075 13.685 ;
        RECT 2234.365 13.515 2234.535 13.685 ;
        RECT 2234.825 13.515 2234.995 13.685 ;
        RECT 2236.665 13.515 2236.835 13.685 ;
        RECT 2238.505 13.515 2238.675 13.685 ;
        RECT 2238.965 13.515 2239.135 13.685 ;
        RECT 2239.425 13.515 2239.595 13.685 ;
        RECT 2240.805 13.515 2240.975 13.685 ;
        RECT 2241.265 13.515 2241.435 13.685 ;
        RECT 2241.725 13.515 2241.895 13.685 ;
        RECT 2244.485 13.515 2244.655 13.685 ;
        RECT 2258.745 13.515 2258.915 13.685 ;
        RECT 2264.725 13.515 2264.895 13.685 ;
        RECT 2271.625 13.515 2271.795 13.685 ;
        RECT 2272.085 13.515 2272.255 13.685 ;
        RECT 2272.545 13.515 2272.715 13.685 ;
        RECT 2273.005 13.515 2273.175 13.685 ;
        RECT 2276.685 13.515 2276.855 13.685 ;
        RECT 2277.145 13.515 2277.315 13.685 ;
        RECT 2277.605 13.515 2277.775 13.685 ;
        RECT 2287.265 13.515 2287.435 13.685 ;
        RECT 2292.785 13.515 2292.955 13.685 ;
        RECT 2296.465 13.515 2296.635 13.685 ;
        RECT 2296.925 13.515 2297.095 13.685 ;
        RECT 2297.385 13.515 2297.555 13.685 ;
        RECT 2301.525 13.515 2301.695 13.685 ;
        RECT 2315.785 13.515 2315.955 13.685 ;
        RECT 2320.845 13.515 2321.015 13.685 ;
        RECT 2321.305 13.515 2321.475 13.685 ;
        RECT 2321.765 13.515 2321.935 13.685 ;
        RECT 2322.225 13.515 2322.395 13.685 ;
        RECT 2330.045 13.515 2330.215 13.685 ;
        RECT 2344.305 13.515 2344.475 13.685 ;
        RECT 2348.905 13.515 2349.075 13.685 ;
        RECT 2358.565 13.515 2358.735 13.685 ;
        RECT 2372.825 13.515 2372.995 13.685 ;
        RECT 2376.965 13.515 2377.135 13.685 ;
        RECT 2387.085 13.515 2387.255 13.685 ;
        RECT 2401.345 13.515 2401.515 13.685 ;
        RECT 2405.025 13.515 2405.195 13.685 ;
        RECT 2415.605 13.515 2415.775 13.685 ;
        RECT 2427.565 13.515 2427.735 13.685 ;
        RECT 2428.025 13.515 2428.195 13.685 ;
        RECT 2428.485 13.515 2428.655 13.685 ;
        RECT 2429.865 13.515 2430.035 13.685 ;
        RECT 2433.085 13.515 2433.255 13.685 ;
        RECT 2439.525 13.515 2439.695 13.685 ;
        RECT 2439.985 13.515 2440.155 13.685 ;
        RECT 2440.445 13.515 2440.615 13.685 ;
        RECT 2444.125 13.515 2444.295 13.685 ;
        RECT 2458.385 13.515 2458.555 13.685 ;
        RECT 2461.145 13.515 2461.315 13.685 ;
        RECT 2472.645 13.515 2472.815 13.685 ;
        RECT 2486.905 13.515 2487.075 13.685 ;
        RECT 2489.205 13.515 2489.375 13.685 ;
        RECT 2490.125 13.515 2490.295 13.685 ;
        RECT 2490.585 13.515 2490.755 13.685 ;
        RECT 2491.045 13.515 2491.215 13.685 ;
        RECT 2496.105 13.515 2496.275 13.685 ;
        RECT 2496.565 13.515 2496.735 13.685 ;
        RECT 2497.025 13.515 2497.195 13.685 ;
        RECT 2497.485 13.515 2497.655 13.685 ;
        RECT 2497.945 13.515 2498.115 13.685 ;
        RECT 2498.405 13.515 2498.575 13.685 ;
        RECT 2500.245 13.515 2500.415 13.685 ;
        RECT 2500.705 13.515 2500.875 13.685 ;
        RECT 2501.165 13.515 2501.335 13.685 ;
        RECT 2501.625 13.515 2501.795 13.685 ;
        RECT 2502.085 13.515 2502.255 13.685 ;
        RECT 2502.545 13.515 2502.715 13.685 ;
        RECT 2509.445 13.515 2509.615 13.685 ;
        RECT 2509.905 13.515 2510.075 13.685 ;
        RECT 2510.365 13.515 2510.535 13.685 ;
        RECT 2515.425 13.515 2515.595 13.685 ;
        RECT 2517.265 13.515 2517.435 13.685 ;
        RECT 2525.085 13.515 2525.255 13.685 ;
        RECT 2525.545 13.515 2525.715 13.685 ;
        RECT 2526.005 13.515 2526.175 13.685 ;
        RECT 2529.685 13.515 2529.855 13.685 ;
        RECT 2530.145 13.515 2530.315 13.685 ;
        RECT 2530.605 13.515 2530.775 13.685 ;
        RECT 2531.065 13.515 2531.235 13.685 ;
        RECT 2533.825 13.515 2533.995 13.685 ;
        RECT 2534.285 13.515 2534.455 13.685 ;
        RECT 2534.745 13.515 2534.915 13.685 ;
        RECT 2543.945 13.515 2544.115 13.685 ;
        RECT 2545.325 13.515 2545.495 13.685 ;
        RECT 2547.625 13.515 2547.795 13.685 ;
        RECT 2548.085 13.515 2548.255 13.685 ;
        RECT 2548.545 13.515 2548.715 13.685 ;
        RECT 2551.305 13.515 2551.475 13.685 ;
        RECT 2551.765 13.515 2551.935 13.685 ;
        RECT 2552.225 13.515 2552.395 13.685 ;
        RECT 2554.065 13.515 2554.235 13.685 ;
        RECT 2554.525 13.515 2554.695 13.685 ;
        RECT 2554.985 13.515 2555.155 13.685 ;
        RECT 2558.205 13.515 2558.375 13.685 ;
        RECT 2569.245 13.515 2569.415 13.685 ;
        RECT 2569.705 13.515 2569.875 13.685 ;
        RECT 2570.165 13.515 2570.335 13.685 ;
        RECT 2572.465 13.515 2572.635 13.685 ;
        RECT 2573.385 13.515 2573.555 13.685 ;
        RECT 2580.745 13.515 2580.915 13.685 ;
        RECT 2581.205 13.515 2581.375 13.685 ;
        RECT 2581.665 13.515 2581.835 13.685 ;
        RECT 2585.805 13.515 2585.975 13.685 ;
        RECT 2586.265 13.515 2586.435 13.685 ;
        RECT 2586.725 13.515 2586.895 13.685 ;
        RECT 2592.705 13.515 2592.875 13.685 ;
        RECT 2593.165 13.515 2593.335 13.685 ;
        RECT 2593.625 13.515 2593.795 13.685 ;
        RECT 2597.765 13.515 2597.935 13.685 ;
        RECT 2598.225 13.515 2598.395 13.685 ;
        RECT 2598.685 13.515 2598.855 13.685 ;
        RECT 2600.985 13.515 2601.155 13.685 ;
        RECT 2601.445 13.515 2601.615 13.685 ;
        RECT 2609.265 13.515 2609.435 13.685 ;
        RECT 2609.725 13.515 2609.895 13.685 ;
        RECT 2610.185 13.515 2610.355 13.685 ;
        RECT 2615.245 13.515 2615.415 13.685 ;
        RECT 2629.505 13.515 2629.675 13.685 ;
        RECT 2643.765 13.515 2643.935 13.685 ;
        RECT 2655.265 13.515 2655.435 13.685 ;
        RECT 2655.725 13.515 2655.895 13.685 ;
        RECT 2656.185 13.515 2656.355 13.685 ;
        RECT 2657.565 13.515 2657.735 13.685 ;
        RECT 2658.025 13.515 2658.195 13.685 ;
        RECT 2672.285 13.515 2672.455 13.685 ;
        RECT 2685.625 13.515 2685.795 13.685 ;
        RECT 2686.085 13.515 2686.255 13.685 ;
        RECT 2686.545 13.515 2686.715 13.685 ;
        RECT 2687.005 13.515 2687.175 13.685 ;
        RECT 2688.385 13.515 2688.555 13.685 ;
        RECT 2688.845 13.515 2689.015 13.685 ;
        RECT 2689.305 13.515 2689.475 13.685 ;
        RECT 2700.805 13.515 2700.975 13.685 ;
        RECT 2713.685 13.515 2713.855 13.685 ;
        RECT 2715.065 13.515 2715.235 13.685 ;
        RECT 2725.645 13.515 2725.815 13.685 ;
        RECT 2726.105 13.515 2726.275 13.685 ;
        RECT 2726.565 13.515 2726.735 13.685 ;
        RECT 2727.025 13.515 2727.195 13.685 ;
        RECT 2727.485 13.515 2727.655 13.685 ;
        RECT 2727.945 13.515 2728.115 13.685 ;
        RECT 2729.325 13.515 2729.495 13.685 ;
        RECT 2730.245 13.515 2730.415 13.685 ;
        RECT 2730.705 13.515 2730.875 13.685 ;
        RECT 2731.165 13.515 2731.335 13.685 ;
        RECT 2741.745 13.515 2741.915 13.685 ;
        RECT 2743.585 13.515 2743.755 13.685 ;
        RECT 2757.845 13.515 2758.015 13.685 ;
        RECT 2769.805 13.515 2769.975 13.685 ;
        RECT 2772.105 13.515 2772.275 13.685 ;
        RECT 2786.365 13.515 2786.535 13.685 ;
        RECT 2797.865 13.515 2798.035 13.685 ;
        RECT 2800.625 13.515 2800.795 13.685 ;
        RECT 2814.885 13.515 2815.055 13.685 ;
        RECT 2825.925 13.515 2826.095 13.685 ;
        RECT 2829.145 13.515 2829.315 13.685 ;
        RECT 2843.405 13.515 2843.575 13.685 ;
        RECT 2853.985 13.515 2854.155 13.685 ;
        RECT 2855.365 13.515 2855.535 13.685 ;
        RECT 2855.825 13.515 2855.995 13.685 ;
        RECT 2856.285 13.515 2856.455 13.685 ;
        RECT 2857.665 13.515 2857.835 13.685 ;
        RECT 2871.925 13.515 2872.095 13.685 ;
        RECT 2882.045 13.515 2882.215 13.685 ;
        RECT 2886.185 13.515 2886.355 13.685 ;
        RECT 2900.445 13.515 2900.615 13.685 ;
        RECT 2907.345 13.515 2907.515 13.685 ;
        RECT 2907.805 13.515 2907.975 13.685 ;
        RECT 2908.265 13.515 2908.435 13.685 ;
        RECT 2908.725 13.515 2908.895 13.685 ;
        RECT 2909.185 13.515 2909.355 13.685 ;
        RECT 2909.645 13.515 2909.815 13.685 ;
        RECT 2910.105 13.515 2910.275 13.685 ;
        RECT 2910.565 13.515 2910.735 13.685 ;
        RECT 2911.025 13.515 2911.195 13.685 ;
        RECT 2911.485 13.515 2911.655 13.685 ;
        RECT 2912.865 13.515 2913.035 13.685 ;
        RECT 2913.325 13.515 2913.495 13.685 ;
        RECT 2913.785 13.515 2913.955 13.685 ;
      LAYER met1 ;
        RECT 5.520 3506.300 2914.100 3506.320 ;
        RECT 5.520 3505.840 13.700 3506.300 ;
        RECT 2906.300 3505.840 2914.100 3506.300 ;
        RECT 5.520 3500.400 13.700 3500.880 ;
        RECT 2906.300 3500.400 2914.100 3500.880 ;
        RECT 5.520 3494.960 13.700 3495.440 ;
        RECT 2906.300 3494.960 2914.100 3495.440 ;
        RECT 5.520 3489.520 13.700 3490.000 ;
        RECT 2906.300 3489.520 2914.100 3490.000 ;
        RECT 5.520 3484.080 13.700 3484.560 ;
        RECT 2906.300 3484.080 2914.100 3484.560 ;
        RECT 5.520 3478.640 13.700 3479.120 ;
        RECT 2906.300 3478.640 2914.100 3479.120 ;
        RECT 5.520 3473.200 13.700 3473.680 ;
        RECT 2906.300 3473.200 2914.100 3473.680 ;
        RECT 5.520 3467.760 13.700 3468.240 ;
        RECT 2906.300 3467.760 2914.100 3468.240 ;
        RECT 5.520 3462.320 13.700 3462.800 ;
        RECT 2906.300 3462.320 2914.100 3462.800 ;
        RECT 5.520 3456.880 13.700 3457.360 ;
        RECT 2906.300 3456.880 2914.100 3457.360 ;
        RECT 5.520 3451.440 13.700 3451.920 ;
        RECT 2906.300 3451.440 2914.100 3451.920 ;
        RECT 5.520 3446.000 13.700 3446.480 ;
        RECT 2906.300 3446.000 2914.100 3446.480 ;
        RECT 5.520 3440.560 13.700 3441.040 ;
        RECT 2906.300 3440.560 2914.100 3441.040 ;
        RECT 5.520 3435.120 13.700 3435.600 ;
        RECT 2906.300 3435.120 2914.100 3435.600 ;
        RECT 5.520 3429.680 13.700 3430.160 ;
        RECT 2906.300 3429.680 2914.100 3430.160 ;
        RECT 5.520 3424.240 13.700 3424.720 ;
        RECT 2906.300 3424.240 2914.100 3424.720 ;
        RECT 5.520 3418.800 13.700 3419.280 ;
        RECT 2906.300 3418.800 2914.100 3419.280 ;
        RECT 5.520 3413.360 13.700 3413.840 ;
        RECT 2906.300 3413.360 2914.100 3413.840 ;
        RECT 5.520 3407.920 13.700 3408.400 ;
        RECT 2906.300 3407.920 2914.100 3408.400 ;
        RECT 5.520 3402.480 13.700 3402.960 ;
        RECT 2906.300 3402.480 2914.100 3402.960 ;
        RECT 5.520 3397.040 13.700 3397.520 ;
        RECT 2906.300 3397.040 2914.100 3397.520 ;
        RECT 5.520 3391.600 13.700 3392.080 ;
        RECT 2906.300 3391.600 2914.100 3392.080 ;
        RECT 5.520 3386.160 13.700 3386.640 ;
        RECT 2906.300 3386.160 2914.100 3386.640 ;
        RECT 5.520 3380.720 13.700 3381.200 ;
        RECT 2906.300 3380.720 2914.100 3381.200 ;
        RECT 5.520 3375.280 13.700 3375.760 ;
        RECT 2906.300 3375.280 2914.100 3375.760 ;
        RECT 5.520 3369.840 13.700 3370.320 ;
        RECT 2906.300 3369.840 2914.100 3370.320 ;
        RECT 5.520 3364.400 13.700 3364.880 ;
        RECT 2906.300 3364.400 2914.100 3364.880 ;
        RECT 5.520 3358.960 13.700 3359.440 ;
        RECT 2906.300 3358.960 2914.100 3359.440 ;
        RECT 5.520 3353.520 13.700 3354.000 ;
        RECT 2906.300 3353.520 2914.100 3354.000 ;
        RECT 5.520 3348.080 13.700 3348.560 ;
        RECT 2906.300 3348.080 2914.100 3348.560 ;
        RECT 5.520 3342.640 13.700 3343.120 ;
        RECT 2906.300 3342.640 2914.100 3343.120 ;
        RECT 5.520 3337.200 13.700 3337.680 ;
        RECT 2906.300 3337.200 2914.100 3337.680 ;
        RECT 5.520 3331.760 13.700 3332.240 ;
        RECT 2906.300 3331.760 2914.100 3332.240 ;
        RECT 5.520 3326.320 13.700 3326.800 ;
        RECT 2906.300 3326.320 2914.100 3326.800 ;
        RECT 5.520 3320.880 13.700 3321.360 ;
        RECT 2906.300 3320.880 2914.100 3321.360 ;
        RECT 5.520 3315.440 13.700 3315.920 ;
        RECT 2906.300 3315.440 2914.100 3315.920 ;
        RECT 5.520 3310.000 13.700 3310.480 ;
        RECT 2906.300 3310.000 2914.100 3310.480 ;
        RECT 5.520 3304.560 13.700 3305.040 ;
        RECT 2906.300 3304.560 2914.100 3305.040 ;
        RECT 5.520 3299.120 13.700 3299.600 ;
        RECT 2906.300 3299.120 2914.100 3299.600 ;
        RECT 5.520 3293.680 13.700 3294.160 ;
        RECT 2906.300 3293.680 2914.100 3294.160 ;
        RECT 5.520 3288.240 13.700 3288.720 ;
        RECT 2906.300 3288.240 2914.100 3288.720 ;
        RECT 5.520 3282.800 13.700 3283.280 ;
        RECT 2906.300 3282.800 2914.100 3283.280 ;
        RECT 5.520 3277.360 13.700 3277.840 ;
        RECT 2906.300 3277.360 2914.100 3277.840 ;
        RECT 5.520 3271.920 13.700 3272.400 ;
        RECT 2906.300 3271.920 2914.100 3272.400 ;
        RECT 5.520 3266.480 13.700 3266.960 ;
        RECT 2906.300 3266.480 2914.100 3266.960 ;
        RECT 5.520 3261.040 13.700 3261.520 ;
        RECT 2906.300 3261.040 2914.100 3261.520 ;
        RECT 5.520 3255.600 13.700 3256.080 ;
        RECT 2906.300 3255.600 2914.100 3256.080 ;
        RECT 5.520 3250.160 13.700 3250.640 ;
        RECT 2906.300 3250.160 2914.100 3250.640 ;
        RECT 5.520 3244.720 13.700 3245.200 ;
        RECT 2906.300 3244.720 2914.100 3245.200 ;
        RECT 5.520 3239.280 13.700 3239.760 ;
        RECT 2906.300 3239.280 2914.100 3239.760 ;
        RECT 5.520 3233.840 13.700 3234.320 ;
        RECT 2906.300 3233.840 2914.100 3234.320 ;
        RECT 5.520 3228.400 13.700 3228.880 ;
        RECT 2906.300 3228.400 2914.100 3228.880 ;
        RECT 5.520 3222.960 13.700 3223.440 ;
        RECT 2906.300 3222.960 2914.100 3223.440 ;
        RECT 5.520 3217.520 13.700 3218.000 ;
        RECT 2906.300 3217.520 2914.100 3218.000 ;
        RECT 5.520 3212.080 13.700 3212.560 ;
        RECT 2906.300 3212.080 2914.100 3212.560 ;
        RECT 5.520 3206.640 13.700 3207.120 ;
        RECT 2906.300 3206.640 2914.100 3207.120 ;
        RECT 5.520 3201.200 13.700 3201.680 ;
        RECT 2906.300 3201.200 2914.100 3201.680 ;
        RECT 5.520 3195.760 13.700 3196.240 ;
        RECT 2906.300 3195.760 2914.100 3196.240 ;
        RECT 5.520 3190.320 13.700 3190.800 ;
        RECT 2906.300 3190.320 2914.100 3190.800 ;
        RECT 5.520 3184.880 13.700 3185.360 ;
        RECT 2906.300 3184.880 2914.100 3185.360 ;
        RECT 5.520 3179.440 13.700 3179.920 ;
        RECT 2906.300 3179.440 2914.100 3179.920 ;
        RECT 5.520 3174.000 13.700 3174.480 ;
        RECT 2906.300 3174.000 2914.100 3174.480 ;
        RECT 5.520 3168.560 13.700 3169.040 ;
        RECT 2906.300 3168.560 2914.100 3169.040 ;
        RECT 5.520 3163.120 13.700 3163.600 ;
        RECT 2906.300 3163.120 2914.100 3163.600 ;
        RECT 5.520 3157.680 13.700 3158.160 ;
        RECT 2906.300 3157.680 2914.100 3158.160 ;
        RECT 5.520 3152.240 13.700 3152.720 ;
        RECT 2906.300 3152.240 2914.100 3152.720 ;
        RECT 5.520 3146.800 13.700 3147.280 ;
        RECT 2906.300 3146.800 2914.100 3147.280 ;
        RECT 5.520 3141.360 13.700 3141.840 ;
        RECT 2906.300 3141.360 2914.100 3141.840 ;
        RECT 5.520 3135.920 13.700 3136.400 ;
        RECT 2906.300 3135.920 2914.100 3136.400 ;
        RECT 5.520 3130.480 13.700 3130.960 ;
        RECT 2906.300 3130.480 2914.100 3130.960 ;
        RECT 5.520 3125.040 13.700 3125.520 ;
        RECT 2906.300 3125.040 2914.100 3125.520 ;
        RECT 5.520 3119.600 13.700 3120.080 ;
        RECT 2906.300 3119.600 2914.100 3120.080 ;
        RECT 5.520 3114.160 13.700 3114.640 ;
        RECT 2906.300 3114.160 2914.100 3114.640 ;
        RECT 5.520 3108.720 13.700 3109.200 ;
        RECT 2906.300 3108.720 2914.100 3109.200 ;
        RECT 5.520 3103.280 13.700 3103.760 ;
        RECT 2906.300 3103.280 2914.100 3103.760 ;
        RECT 5.520 3097.840 13.700 3098.320 ;
        RECT 2906.300 3097.840 2914.100 3098.320 ;
        RECT 5.520 3092.400 13.700 3092.880 ;
        RECT 2906.300 3092.400 2914.100 3092.880 ;
        RECT 5.520 3086.960 13.700 3087.440 ;
        RECT 2906.300 3086.960 2914.100 3087.440 ;
        RECT 5.520 3081.520 13.700 3082.000 ;
        RECT 2906.300 3081.520 2914.100 3082.000 ;
        RECT 5.520 3076.080 13.700 3076.560 ;
        RECT 2906.300 3076.080 2914.100 3076.560 ;
        RECT 5.520 3070.640 13.700 3071.120 ;
        RECT 2906.300 3070.640 2914.100 3071.120 ;
        RECT 5.520 3065.200 13.700 3065.680 ;
        RECT 2906.300 3065.200 2914.100 3065.680 ;
        RECT 5.520 3059.760 13.700 3060.240 ;
        RECT 2906.300 3059.760 2914.100 3060.240 ;
        RECT 5.520 3054.320 13.700 3054.800 ;
        RECT 2906.300 3054.320 2914.100 3054.800 ;
        RECT 5.520 3048.880 13.700 3049.360 ;
        RECT 2906.300 3048.880 2914.100 3049.360 ;
        RECT 5.520 3043.440 13.700 3043.920 ;
        RECT 2906.300 3043.440 2914.100 3043.920 ;
        RECT 5.520 3038.000 13.700 3038.480 ;
        RECT 2906.300 3038.000 2914.100 3038.480 ;
        RECT 5.520 3032.560 13.700 3033.040 ;
        RECT 2906.300 3032.560 2914.100 3033.040 ;
        RECT 5.520 3027.120 13.700 3027.600 ;
        RECT 2906.300 3027.120 2914.100 3027.600 ;
        RECT 5.520 3021.680 13.700 3022.160 ;
        RECT 2906.300 3021.680 2914.100 3022.160 ;
        RECT 5.520 3016.240 13.700 3016.720 ;
        RECT 2906.300 3016.240 2914.100 3016.720 ;
        RECT 5.520 3010.800 13.700 3011.280 ;
        RECT 2906.300 3010.800 2914.100 3011.280 ;
        RECT 5.520 3005.360 13.700 3005.840 ;
        RECT 2906.300 3005.360 2914.100 3005.840 ;
        RECT 5.520 2999.920 13.700 3000.400 ;
        RECT 2906.300 2999.920 2914.100 3000.400 ;
        RECT 5.520 2994.480 13.700 2994.960 ;
        RECT 2906.300 2994.480 2914.100 2994.960 ;
        RECT 5.520 2989.040 13.700 2989.520 ;
        RECT 2906.300 2989.040 2914.100 2989.520 ;
        RECT 5.520 2983.600 13.700 2984.080 ;
        RECT 2906.300 2983.600 2914.100 2984.080 ;
        RECT 5.520 2978.160 13.700 2978.640 ;
        RECT 2906.300 2978.160 2914.100 2978.640 ;
        RECT 5.520 2972.720 13.700 2973.200 ;
        RECT 2906.300 2972.720 2914.100 2973.200 ;
        RECT 5.520 2967.280 13.700 2967.760 ;
        RECT 2906.300 2967.280 2914.100 2967.760 ;
        RECT 5.520 2961.840 13.700 2962.320 ;
        RECT 2906.300 2961.840 2914.100 2962.320 ;
        RECT 5.520 2956.400 13.700 2956.880 ;
        RECT 2906.300 2956.400 2914.100 2956.880 ;
        RECT 5.520 2950.960 13.700 2951.440 ;
        RECT 2906.300 2950.960 2914.100 2951.440 ;
        RECT 5.520 2945.520 13.700 2946.000 ;
        RECT 2906.300 2945.520 2914.100 2946.000 ;
        RECT 5.520 2940.080 13.700 2940.560 ;
        RECT 2906.300 2940.080 2914.100 2940.560 ;
        RECT 5.520 2934.640 13.700 2935.120 ;
        RECT 2906.300 2934.640 2914.100 2935.120 ;
        RECT 5.520 2929.200 13.700 2929.680 ;
        RECT 2906.300 2929.200 2914.100 2929.680 ;
        RECT 5.520 2923.760 13.700 2924.240 ;
        RECT 2906.300 2923.760 2914.100 2924.240 ;
        RECT 5.520 2918.320 13.700 2918.800 ;
        RECT 2906.300 2918.320 2914.100 2918.800 ;
        RECT 5.520 2912.880 13.700 2913.360 ;
        RECT 2906.300 2912.880 2914.100 2913.360 ;
        RECT 5.520 2907.440 13.700 2907.920 ;
        RECT 2906.300 2907.440 2914.100 2907.920 ;
        RECT 5.520 2902.000 13.700 2902.480 ;
        RECT 2906.300 2902.000 2914.100 2902.480 ;
        RECT 5.520 2896.560 13.700 2897.040 ;
        RECT 2906.300 2896.560 2914.100 2897.040 ;
        RECT 5.520 2891.120 13.700 2891.600 ;
        RECT 2906.300 2891.120 2914.100 2891.600 ;
        RECT 5.520 2885.680 13.700 2886.160 ;
        RECT 2906.300 2885.680 2914.100 2886.160 ;
        RECT 5.520 2880.240 13.700 2880.720 ;
        RECT 2906.300 2880.240 2914.100 2880.720 ;
        RECT 5.520 2874.800 13.700 2875.280 ;
        RECT 2906.300 2874.800 2914.100 2875.280 ;
        RECT 5.520 2869.360 13.700 2869.840 ;
        RECT 2906.300 2869.360 2914.100 2869.840 ;
        RECT 5.520 2863.920 13.700 2864.400 ;
        RECT 2906.300 2863.920 2914.100 2864.400 ;
        RECT 5.520 2858.480 13.700 2858.960 ;
        RECT 2906.300 2858.480 2914.100 2858.960 ;
        RECT 5.520 2853.040 13.700 2853.520 ;
        RECT 2906.300 2853.040 2914.100 2853.520 ;
        RECT 5.520 2847.600 13.700 2848.080 ;
        RECT 2906.300 2847.600 2914.100 2848.080 ;
        RECT 5.520 2842.160 13.700 2842.640 ;
        RECT 2906.300 2842.160 2914.100 2842.640 ;
        RECT 5.520 2836.720 13.700 2837.200 ;
        RECT 2906.300 2836.720 2914.100 2837.200 ;
        RECT 5.520 2831.280 13.700 2831.760 ;
        RECT 2906.300 2831.280 2914.100 2831.760 ;
        RECT 5.520 2825.840 13.700 2826.320 ;
        RECT 2906.300 2825.840 2914.100 2826.320 ;
        RECT 5.520 2820.400 13.700 2820.880 ;
        RECT 2906.300 2820.400 2914.100 2820.880 ;
        RECT 5.520 2814.960 13.700 2815.440 ;
        RECT 2906.300 2814.960 2914.100 2815.440 ;
        RECT 5.520 2809.520 13.700 2810.000 ;
        RECT 2906.300 2809.520 2914.100 2810.000 ;
        RECT 5.520 2804.080 13.700 2804.560 ;
        RECT 2906.300 2804.080 2914.100 2804.560 ;
        RECT 5.520 2798.640 13.700 2799.120 ;
        RECT 2906.300 2798.640 2914.100 2799.120 ;
        RECT 5.520 2793.200 13.700 2793.680 ;
        RECT 2906.300 2793.200 2914.100 2793.680 ;
        RECT 5.520 2787.760 13.700 2788.240 ;
        RECT 2906.300 2787.760 2914.100 2788.240 ;
        RECT 5.520 2782.320 13.700 2782.800 ;
        RECT 2906.300 2782.320 2914.100 2782.800 ;
        RECT 5.520 2776.880 13.700 2777.360 ;
        RECT 2906.300 2776.880 2914.100 2777.360 ;
        RECT 5.520 2771.440 13.700 2771.920 ;
        RECT 2906.300 2771.440 2914.100 2771.920 ;
        RECT 5.520 2766.000 13.700 2766.480 ;
        RECT 2906.300 2766.000 2914.100 2766.480 ;
        RECT 5.520 2760.560 13.700 2761.040 ;
        RECT 2906.300 2760.560 2914.100 2761.040 ;
        RECT 5.520 2755.120 13.700 2755.600 ;
        RECT 2906.300 2755.120 2914.100 2755.600 ;
        RECT 5.520 2749.680 13.700 2750.160 ;
        RECT 2906.300 2749.680 2914.100 2750.160 ;
        RECT 5.520 2744.240 13.700 2744.720 ;
        RECT 2906.300 2744.240 2914.100 2744.720 ;
        RECT 5.520 2738.800 13.700 2739.280 ;
        RECT 2906.300 2738.800 2914.100 2739.280 ;
        RECT 5.520 2733.360 13.700 2733.840 ;
        RECT 2906.300 2733.360 2914.100 2733.840 ;
        RECT 5.520 2727.920 13.700 2728.400 ;
        RECT 2906.300 2727.920 2914.100 2728.400 ;
        RECT 5.520 2722.480 13.700 2722.960 ;
        RECT 2906.300 2722.480 2914.100 2722.960 ;
        RECT 5.520 2717.040 13.700 2717.520 ;
        RECT 2906.300 2717.040 2914.100 2717.520 ;
        RECT 5.520 2711.600 13.700 2712.080 ;
        RECT 2906.300 2711.600 2914.100 2712.080 ;
        RECT 5.520 2706.160 13.700 2706.640 ;
        RECT 2906.300 2706.160 2914.100 2706.640 ;
        RECT 5.520 2700.720 13.700 2701.200 ;
        RECT 2906.300 2700.720 2914.100 2701.200 ;
        RECT 5.520 2695.280 13.700 2695.760 ;
        RECT 2906.300 2695.280 2914.100 2695.760 ;
        RECT 5.520 2689.840 13.700 2690.320 ;
        RECT 2906.300 2689.840 2914.100 2690.320 ;
        RECT 5.520 2684.400 13.700 2684.880 ;
        RECT 2906.300 2684.400 2914.100 2684.880 ;
        RECT 5.520 2678.960 13.700 2679.440 ;
        RECT 2906.300 2678.960 2914.100 2679.440 ;
        RECT 5.520 2673.520 13.700 2674.000 ;
        RECT 2906.300 2673.520 2914.100 2674.000 ;
        RECT 5.520 2668.080 13.700 2668.560 ;
        RECT 2906.300 2668.080 2914.100 2668.560 ;
        RECT 5.520 2662.640 13.700 2663.120 ;
        RECT 2906.300 2662.640 2914.100 2663.120 ;
        RECT 5.520 2657.200 13.700 2657.680 ;
        RECT 2906.300 2657.200 2914.100 2657.680 ;
        RECT 5.520 2651.760 13.700 2652.240 ;
        RECT 2906.300 2651.760 2914.100 2652.240 ;
        RECT 5.520 2646.320 13.700 2646.800 ;
        RECT 2906.300 2646.320 2914.100 2646.800 ;
        RECT 5.520 2640.880 13.700 2641.360 ;
        RECT 2906.300 2640.880 2914.100 2641.360 ;
        RECT 5.520 2635.440 13.700 2635.920 ;
        RECT 2906.300 2635.440 2914.100 2635.920 ;
        RECT 5.520 2630.000 13.700 2630.480 ;
        RECT 2906.300 2630.000 2914.100 2630.480 ;
        RECT 5.520 2624.560 13.700 2625.040 ;
        RECT 2906.300 2624.560 2914.100 2625.040 ;
        RECT 5.520 2619.120 13.700 2619.600 ;
        RECT 2906.300 2619.120 2914.100 2619.600 ;
        RECT 5.520 2613.680 13.700 2614.160 ;
        RECT 2906.300 2613.680 2914.100 2614.160 ;
        RECT 5.520 2608.240 13.700 2608.720 ;
        RECT 2906.300 2608.240 2914.100 2608.720 ;
        RECT 5.520 2602.800 13.700 2603.280 ;
        RECT 2906.300 2602.800 2914.100 2603.280 ;
        RECT 5.520 2597.360 13.700 2597.840 ;
        RECT 2906.300 2597.360 2914.100 2597.840 ;
        RECT 5.520 2591.920 13.700 2592.400 ;
        RECT 2906.300 2591.920 2914.100 2592.400 ;
        RECT 5.520 2586.480 13.700 2586.960 ;
        RECT 2906.300 2586.480 2914.100 2586.960 ;
        RECT 5.520 2581.040 13.700 2581.520 ;
        RECT 2906.300 2581.040 2914.100 2581.520 ;
        RECT 5.520 2575.600 13.700 2576.080 ;
        RECT 2906.300 2575.600 2914.100 2576.080 ;
        RECT 5.520 2570.160 13.700 2570.640 ;
        RECT 2906.300 2570.160 2914.100 2570.640 ;
        RECT 5.520 2564.720 13.700 2565.200 ;
        RECT 2906.300 2564.720 2914.100 2565.200 ;
        RECT 5.520 2559.280 13.700 2559.760 ;
        RECT 2906.300 2559.280 2914.100 2559.760 ;
        RECT 5.520 2553.840 13.700 2554.320 ;
        RECT 2906.300 2553.840 2914.100 2554.320 ;
        RECT 5.520 2548.400 13.700 2548.880 ;
        RECT 2906.300 2548.400 2914.100 2548.880 ;
        RECT 5.520 2542.960 13.700 2543.440 ;
        RECT 2906.300 2542.960 2914.100 2543.440 ;
        RECT 5.520 2537.520 13.700 2538.000 ;
        RECT 2906.300 2537.520 2914.100 2538.000 ;
        RECT 5.520 2532.080 13.700 2532.560 ;
        RECT 2906.300 2532.080 2914.100 2532.560 ;
        RECT 5.520 2526.640 13.700 2527.120 ;
        RECT 2906.300 2526.640 2914.100 2527.120 ;
        RECT 5.520 2521.200 13.700 2521.680 ;
        RECT 2906.300 2521.200 2914.100 2521.680 ;
        RECT 5.520 2515.760 13.700 2516.240 ;
        RECT 2906.300 2515.760 2914.100 2516.240 ;
        RECT 5.520 2510.320 13.700 2510.800 ;
        RECT 2906.300 2510.320 2914.100 2510.800 ;
        RECT 5.520 2504.880 13.700 2505.360 ;
        RECT 2906.300 2504.880 2914.100 2505.360 ;
        RECT 5.520 2499.440 13.700 2499.920 ;
        RECT 2906.300 2499.440 2914.100 2499.920 ;
        RECT 5.520 2494.000 13.700 2494.480 ;
        RECT 2906.300 2494.000 2914.100 2494.480 ;
        RECT 5.520 2488.560 13.700 2489.040 ;
        RECT 2906.300 2488.560 2914.100 2489.040 ;
        RECT 5.520 2483.120 13.700 2483.600 ;
        RECT 2906.300 2483.120 2914.100 2483.600 ;
        RECT 5.520 2477.680 13.700 2478.160 ;
        RECT 2906.300 2477.680 2914.100 2478.160 ;
        RECT 5.520 2472.240 13.700 2472.720 ;
        RECT 2906.300 2472.240 2914.100 2472.720 ;
        RECT 5.520 2466.800 13.700 2467.280 ;
        RECT 2906.300 2466.800 2914.100 2467.280 ;
        RECT 5.520 2461.360 13.700 2461.840 ;
        RECT 2906.300 2461.360 2914.100 2461.840 ;
        RECT 5.520 2455.920 13.700 2456.400 ;
        RECT 2906.300 2455.920 2914.100 2456.400 ;
        RECT 5.520 2450.480 13.700 2450.960 ;
        RECT 2906.300 2450.480 2914.100 2450.960 ;
        RECT 5.520 2445.040 13.700 2445.520 ;
        RECT 2906.300 2445.040 2914.100 2445.520 ;
        RECT 5.520 2439.600 13.700 2440.080 ;
        RECT 2906.300 2439.600 2914.100 2440.080 ;
        RECT 5.520 2434.160 13.700 2434.640 ;
        RECT 2906.300 2434.160 2914.100 2434.640 ;
        RECT 5.520 2428.720 13.700 2429.200 ;
        RECT 2906.300 2428.720 2914.100 2429.200 ;
        RECT 5.520 2423.280 13.700 2423.760 ;
        RECT 2906.300 2423.280 2914.100 2423.760 ;
        RECT 5.520 2417.840 13.700 2418.320 ;
        RECT 2906.300 2417.840 2914.100 2418.320 ;
        RECT 5.520 2412.400 13.700 2412.880 ;
        RECT 2906.300 2412.400 2914.100 2412.880 ;
        RECT 5.520 2406.960 13.700 2407.440 ;
        RECT 2906.300 2406.960 2914.100 2407.440 ;
        RECT 5.520 2401.520 13.700 2402.000 ;
        RECT 2906.300 2401.520 2914.100 2402.000 ;
        RECT 5.520 2396.080 13.700 2396.560 ;
        RECT 2906.300 2396.080 2914.100 2396.560 ;
        RECT 5.520 2390.640 13.700 2391.120 ;
        RECT 2906.300 2390.640 2914.100 2391.120 ;
        RECT 5.520 2385.200 13.700 2385.680 ;
        RECT 2906.300 2385.200 2914.100 2385.680 ;
        RECT 5.520 2379.760 13.700 2380.240 ;
        RECT 2906.300 2379.760 2914.100 2380.240 ;
        RECT 5.520 2374.320 13.700 2374.800 ;
        RECT 2906.300 2374.320 2914.100 2374.800 ;
        RECT 5.520 2368.880 13.700 2369.360 ;
        RECT 2906.300 2368.880 2914.100 2369.360 ;
        RECT 5.520 2363.440 13.700 2363.920 ;
        RECT 2906.300 2363.440 2914.100 2363.920 ;
        RECT 5.520 2358.000 13.700 2358.480 ;
        RECT 2906.300 2358.000 2914.100 2358.480 ;
        RECT 5.520 2352.560 13.700 2353.040 ;
        RECT 2906.300 2352.560 2914.100 2353.040 ;
        RECT 5.520 2347.120 13.700 2347.600 ;
        RECT 2906.300 2347.120 2914.100 2347.600 ;
        RECT 5.520 2341.680 13.700 2342.160 ;
        RECT 2906.300 2341.680 2914.100 2342.160 ;
        RECT 5.520 2336.240 13.700 2336.720 ;
        RECT 2906.300 2336.240 2914.100 2336.720 ;
        RECT 5.520 2330.800 13.700 2331.280 ;
        RECT 2906.300 2330.800 2914.100 2331.280 ;
        RECT 5.520 2325.360 13.700 2325.840 ;
        RECT 2906.300 2325.360 2914.100 2325.840 ;
        RECT 5.520 2319.920 13.700 2320.400 ;
        RECT 2906.300 2319.920 2914.100 2320.400 ;
        RECT 5.520 2314.480 13.700 2314.960 ;
        RECT 2906.300 2314.480 2914.100 2314.960 ;
        RECT 5.520 2309.040 13.700 2309.520 ;
        RECT 2906.300 2309.040 2914.100 2309.520 ;
        RECT 5.520 2303.600 13.700 2304.080 ;
        RECT 2906.300 2303.600 2914.100 2304.080 ;
        RECT 5.520 2298.160 13.700 2298.640 ;
        RECT 2906.300 2298.160 2914.100 2298.640 ;
        RECT 5.520 2292.720 13.700 2293.200 ;
        RECT 2906.300 2292.720 2914.100 2293.200 ;
        RECT 5.520 2287.280 13.700 2287.760 ;
        RECT 2906.300 2287.280 2914.100 2287.760 ;
        RECT 5.520 2281.840 13.700 2282.320 ;
        RECT 2906.300 2281.840 2914.100 2282.320 ;
        RECT 5.520 2276.400 13.700 2276.880 ;
        RECT 2906.300 2276.400 2914.100 2276.880 ;
        RECT 5.520 2270.960 13.700 2271.440 ;
        RECT 2906.300 2270.960 2914.100 2271.440 ;
        RECT 5.520 2265.520 13.700 2266.000 ;
        RECT 2906.300 2265.520 2914.100 2266.000 ;
        RECT 5.520 2260.080 13.700 2260.560 ;
        RECT 2906.300 2260.080 2914.100 2260.560 ;
        RECT 5.520 2254.640 13.700 2255.120 ;
        RECT 2906.300 2254.640 2914.100 2255.120 ;
        RECT 5.520 2249.200 13.700 2249.680 ;
        RECT 2906.300 2249.200 2914.100 2249.680 ;
        RECT 5.520 2243.760 13.700 2244.240 ;
        RECT 2906.300 2243.760 2914.100 2244.240 ;
        RECT 5.520 2238.320 13.700 2238.800 ;
        RECT 2906.300 2238.320 2914.100 2238.800 ;
        RECT 5.520 2232.880 13.700 2233.360 ;
        RECT 2906.300 2232.880 2914.100 2233.360 ;
        RECT 5.520 2227.440 13.700 2227.920 ;
        RECT 2906.300 2227.440 2914.100 2227.920 ;
        RECT 5.520 2222.000 13.700 2222.480 ;
        RECT 2906.300 2222.000 2914.100 2222.480 ;
        RECT 5.520 2216.560 13.700 2217.040 ;
        RECT 2906.300 2216.560 2914.100 2217.040 ;
        RECT 5.520 2211.120 13.700 2211.600 ;
        RECT 2906.300 2211.120 2914.100 2211.600 ;
        RECT 5.520 2205.680 13.700 2206.160 ;
        RECT 2906.300 2205.680 2914.100 2206.160 ;
        RECT 5.520 2200.240 13.700 2200.720 ;
        RECT 2906.300 2200.240 2914.100 2200.720 ;
        RECT 5.520 2194.800 13.700 2195.280 ;
        RECT 2906.300 2194.800 2914.100 2195.280 ;
        RECT 5.520 2189.360 13.700 2189.840 ;
        RECT 2906.300 2189.360 2914.100 2189.840 ;
        RECT 5.520 2183.920 13.700 2184.400 ;
        RECT 2906.300 2183.920 2914.100 2184.400 ;
        RECT 5.520 2178.480 13.700 2178.960 ;
        RECT 2906.300 2178.480 2914.100 2178.960 ;
        RECT 5.520 2173.040 13.700 2173.520 ;
        RECT 2906.300 2173.040 2914.100 2173.520 ;
        RECT 5.520 2167.600 13.700 2168.080 ;
        RECT 2906.300 2167.600 2914.100 2168.080 ;
        RECT 5.520 2162.160 13.700 2162.640 ;
        RECT 2906.300 2162.160 2914.100 2162.640 ;
        RECT 5.520 2156.720 13.700 2157.200 ;
        RECT 2906.300 2156.720 2914.100 2157.200 ;
        RECT 5.520 2151.280 13.700 2151.760 ;
        RECT 2906.300 2151.280 2914.100 2151.760 ;
        RECT 5.520 2145.840 13.700 2146.320 ;
        RECT 2906.300 2145.840 2914.100 2146.320 ;
        RECT 5.520 2140.400 13.700 2140.880 ;
        RECT 2906.300 2140.400 2914.100 2140.880 ;
        RECT 5.520 2134.960 13.700 2135.440 ;
        RECT 2906.300 2134.960 2914.100 2135.440 ;
        RECT 5.520 2129.520 13.700 2130.000 ;
        RECT 2906.300 2129.520 2914.100 2130.000 ;
        RECT 5.520 2124.080 13.700 2124.560 ;
        RECT 2906.300 2124.080 2914.100 2124.560 ;
        RECT 5.520 2118.640 13.700 2119.120 ;
        RECT 2906.300 2118.640 2914.100 2119.120 ;
        RECT 5.520 2113.200 13.700 2113.680 ;
        RECT 2906.300 2113.200 2914.100 2113.680 ;
        RECT 5.520 2107.760 13.700 2108.240 ;
        RECT 2906.300 2107.760 2914.100 2108.240 ;
        RECT 5.520 2102.320 13.700 2102.800 ;
        RECT 2906.300 2102.320 2914.100 2102.800 ;
        RECT 5.520 2096.880 13.700 2097.360 ;
        RECT 2906.300 2096.880 2914.100 2097.360 ;
        RECT 5.520 2091.440 13.700 2091.920 ;
        RECT 2906.300 2091.440 2914.100 2091.920 ;
        RECT 5.520 2086.000 13.700 2086.480 ;
        RECT 2906.300 2086.000 2914.100 2086.480 ;
        RECT 5.520 2080.560 13.700 2081.040 ;
        RECT 2906.300 2080.560 2914.100 2081.040 ;
        RECT 5.520 2075.120 13.700 2075.600 ;
        RECT 2906.300 2075.120 2914.100 2075.600 ;
        RECT 5.520 2069.680 13.700 2070.160 ;
        RECT 2906.300 2069.680 2914.100 2070.160 ;
        RECT 5.520 2064.240 13.700 2064.720 ;
        RECT 2906.300 2064.240 2914.100 2064.720 ;
        RECT 5.520 2058.800 13.700 2059.280 ;
        RECT 2906.300 2058.800 2914.100 2059.280 ;
        RECT 5.520 2053.360 13.700 2053.840 ;
        RECT 2906.300 2053.360 2914.100 2053.840 ;
        RECT 5.520 2047.920 13.700 2048.400 ;
        RECT 2906.300 2047.920 2914.100 2048.400 ;
        RECT 5.520 2042.480 13.700 2042.960 ;
        RECT 2906.300 2042.480 2914.100 2042.960 ;
        RECT 5.520 2037.040 13.700 2037.520 ;
        RECT 2906.300 2037.040 2914.100 2037.520 ;
        RECT 5.520 2031.600 13.700 2032.080 ;
        RECT 2906.300 2031.600 2914.100 2032.080 ;
        RECT 5.520 2026.160 13.700 2026.640 ;
        RECT 2906.300 2026.160 2914.100 2026.640 ;
        RECT 5.520 2020.720 13.700 2021.200 ;
        RECT 2906.300 2020.720 2914.100 2021.200 ;
        RECT 5.520 2015.280 13.700 2015.760 ;
        RECT 2906.300 2015.280 2914.100 2015.760 ;
        RECT 5.520 2009.840 13.700 2010.320 ;
        RECT 2906.300 2009.840 2914.100 2010.320 ;
        RECT 5.520 2004.400 13.700 2004.880 ;
        RECT 2906.300 2004.400 2914.100 2004.880 ;
        RECT 5.520 1998.960 13.700 1999.440 ;
        RECT 2906.300 1998.960 2914.100 1999.440 ;
        RECT 5.520 1993.520 13.700 1994.000 ;
        RECT 2906.300 1993.520 2914.100 1994.000 ;
        RECT 5.520 1988.080 13.700 1988.560 ;
        RECT 2906.300 1988.080 2914.100 1988.560 ;
        RECT 5.520 1982.640 13.700 1983.120 ;
        RECT 2906.300 1982.640 2914.100 1983.120 ;
        RECT 5.520 1977.200 13.700 1977.680 ;
        RECT 2906.300 1977.200 2914.100 1977.680 ;
        RECT 5.520 1971.760 13.700 1972.240 ;
        RECT 2906.300 1971.760 2914.100 1972.240 ;
        RECT 5.520 1966.320 13.700 1966.800 ;
        RECT 2906.300 1966.320 2914.100 1966.800 ;
        RECT 5.520 1960.880 13.700 1961.360 ;
        RECT 2906.300 1960.880 2914.100 1961.360 ;
        RECT 5.520 1955.440 13.700 1955.920 ;
        RECT 2906.300 1955.440 2914.100 1955.920 ;
        RECT 5.520 1950.000 13.700 1950.480 ;
        RECT 2906.300 1950.000 2914.100 1950.480 ;
        RECT 5.520 1944.560 13.700 1945.040 ;
        RECT 2906.300 1944.560 2914.100 1945.040 ;
        RECT 5.520 1939.120 13.700 1939.600 ;
        RECT 2906.300 1939.120 2914.100 1939.600 ;
        RECT 5.520 1933.680 13.700 1934.160 ;
        RECT 2906.300 1933.680 2914.100 1934.160 ;
        RECT 5.520 1928.240 13.700 1928.720 ;
        RECT 2906.300 1928.240 2914.100 1928.720 ;
        RECT 5.520 1922.800 13.700 1923.280 ;
        RECT 2906.300 1922.800 2914.100 1923.280 ;
        RECT 5.520 1917.360 13.700 1917.840 ;
        RECT 2906.300 1917.360 2914.100 1917.840 ;
        RECT 5.520 1911.920 13.700 1912.400 ;
        RECT 2906.300 1911.920 2914.100 1912.400 ;
        RECT 5.520 1906.480 13.700 1906.960 ;
        RECT 2906.300 1906.480 2914.100 1906.960 ;
        RECT 5.520 1901.040 13.700 1901.520 ;
        RECT 2906.300 1901.040 2914.100 1901.520 ;
        RECT 5.520 1895.600 13.700 1896.080 ;
        RECT 2906.300 1895.600 2914.100 1896.080 ;
        RECT 5.520 1890.160 13.700 1890.640 ;
        RECT 2906.300 1890.160 2914.100 1890.640 ;
        RECT 5.520 1884.720 13.700 1885.200 ;
        RECT 2906.300 1884.720 2914.100 1885.200 ;
        RECT 5.520 1879.280 13.700 1879.760 ;
        RECT 2906.300 1879.280 2914.100 1879.760 ;
        RECT 5.520 1873.840 13.700 1874.320 ;
        RECT 2906.300 1873.840 2914.100 1874.320 ;
        RECT 5.520 1868.400 13.700 1868.880 ;
        RECT 2906.300 1868.400 2914.100 1868.880 ;
        RECT 5.520 1862.960 13.700 1863.440 ;
        RECT 2906.300 1862.960 2914.100 1863.440 ;
        RECT 5.520 1857.520 13.700 1858.000 ;
        RECT 2906.300 1857.520 2914.100 1858.000 ;
        RECT 5.520 1852.080 13.700 1852.560 ;
        RECT 2906.300 1852.080 2914.100 1852.560 ;
        RECT 5.520 1846.640 13.700 1847.120 ;
        RECT 2906.300 1846.640 2914.100 1847.120 ;
        RECT 5.520 1841.200 13.700 1841.680 ;
        RECT 2906.300 1841.200 2914.100 1841.680 ;
        RECT 5.520 1835.760 13.700 1836.240 ;
        RECT 2906.300 1835.760 2914.100 1836.240 ;
        RECT 5.520 1830.320 13.700 1830.800 ;
        RECT 2906.300 1830.320 2914.100 1830.800 ;
        RECT 5.520 1824.880 13.700 1825.360 ;
        RECT 2906.300 1824.880 2914.100 1825.360 ;
        RECT 5.520 1819.440 13.700 1819.920 ;
        RECT 2906.300 1819.440 2914.100 1819.920 ;
        RECT 5.520 1814.000 13.700 1814.480 ;
        RECT 2906.300 1814.000 2914.100 1814.480 ;
        RECT 5.520 1808.560 13.700 1809.040 ;
        RECT 2906.300 1808.560 2914.100 1809.040 ;
        RECT 5.520 1803.120 13.700 1803.600 ;
        RECT 2906.300 1803.120 2914.100 1803.600 ;
        RECT 5.520 1797.680 13.700 1798.160 ;
        RECT 2906.300 1797.680 2914.100 1798.160 ;
        RECT 5.520 1792.240 13.700 1792.720 ;
        RECT 2906.300 1792.240 2914.100 1792.720 ;
        RECT 5.520 1786.800 13.700 1787.280 ;
        RECT 2906.300 1786.800 2914.100 1787.280 ;
        RECT 5.520 1781.360 13.700 1781.840 ;
        RECT 2906.300 1781.360 2914.100 1781.840 ;
        RECT 5.520 1775.920 13.700 1776.400 ;
        RECT 2906.300 1775.920 2914.100 1776.400 ;
        RECT 5.520 1770.480 13.700 1770.960 ;
        RECT 2906.300 1770.480 2914.100 1770.960 ;
        RECT 5.520 1765.040 13.700 1765.520 ;
        RECT 2906.300 1765.040 2914.100 1765.520 ;
        RECT 5.520 1759.600 13.700 1760.080 ;
        RECT 2906.300 1759.600 2914.100 1760.080 ;
        RECT 5.520 1754.160 13.700 1754.640 ;
        RECT 2906.300 1754.160 2914.100 1754.640 ;
        RECT 5.520 1748.720 13.700 1749.200 ;
        RECT 2906.300 1748.720 2914.100 1749.200 ;
        RECT 5.520 1743.280 13.700 1743.760 ;
        RECT 2906.300 1743.280 2914.100 1743.760 ;
        RECT 5.520 1737.840 13.700 1738.320 ;
        RECT 2906.300 1737.840 2914.100 1738.320 ;
        RECT 5.520 1732.400 13.700 1732.880 ;
        RECT 2906.300 1732.400 2914.100 1732.880 ;
        RECT 5.520 1726.960 13.700 1727.440 ;
        RECT 2906.300 1726.960 2914.100 1727.440 ;
        RECT 5.520 1721.520 13.700 1722.000 ;
        RECT 2906.300 1721.520 2914.100 1722.000 ;
        RECT 5.520 1716.080 13.700 1716.560 ;
        RECT 2906.300 1716.080 2914.100 1716.560 ;
        RECT 5.520 1710.640 13.700 1711.120 ;
        RECT 2906.300 1710.640 2914.100 1711.120 ;
        RECT 5.520 1705.200 13.700 1705.680 ;
        RECT 2906.300 1705.200 2914.100 1705.680 ;
        RECT 5.520 1699.760 13.700 1700.240 ;
        RECT 2906.300 1699.760 2914.100 1700.240 ;
        RECT 5.520 1694.320 13.700 1694.800 ;
        RECT 2906.300 1694.320 2914.100 1694.800 ;
        RECT 5.520 1688.880 13.700 1689.360 ;
        RECT 2906.300 1688.880 2914.100 1689.360 ;
        RECT 5.520 1683.440 13.700 1683.920 ;
        RECT 2906.300 1683.440 2914.100 1683.920 ;
        RECT 5.520 1678.000 13.700 1678.480 ;
        RECT 2906.300 1678.000 2914.100 1678.480 ;
        RECT 5.520 1672.560 13.700 1673.040 ;
        RECT 2906.300 1672.560 2914.100 1673.040 ;
        RECT 5.520 1667.120 13.700 1667.600 ;
        RECT 2906.300 1667.120 2914.100 1667.600 ;
        RECT 5.520 1661.680 13.700 1662.160 ;
        RECT 2906.300 1661.680 2914.100 1662.160 ;
        RECT 5.520 1656.240 13.700 1656.720 ;
        RECT 2906.300 1656.240 2914.100 1656.720 ;
        RECT 5.520 1650.800 13.700 1651.280 ;
        RECT 2906.300 1650.800 2914.100 1651.280 ;
        RECT 5.520 1645.360 13.700 1645.840 ;
        RECT 2906.300 1645.360 2914.100 1645.840 ;
        RECT 5.520 1639.920 13.700 1640.400 ;
        RECT 2906.300 1639.920 2914.100 1640.400 ;
        RECT 5.520 1634.480 13.700 1634.960 ;
        RECT 2906.300 1634.480 2914.100 1634.960 ;
        RECT 5.520 1629.040 13.700 1629.520 ;
        RECT 2906.300 1629.040 2914.100 1629.520 ;
        RECT 5.520 1623.600 13.700 1624.080 ;
        RECT 2906.300 1623.600 2914.100 1624.080 ;
        RECT 5.520 1618.160 13.700 1618.640 ;
        RECT 2906.300 1618.160 2914.100 1618.640 ;
        RECT 5.520 1612.720 13.700 1613.200 ;
        RECT 2906.300 1612.720 2914.100 1613.200 ;
        RECT 5.520 1607.280 13.700 1607.760 ;
        RECT 2906.300 1607.280 2914.100 1607.760 ;
        RECT 5.520 1601.840 13.700 1602.320 ;
        RECT 2906.300 1601.840 2914.100 1602.320 ;
        RECT 5.520 1596.400 13.700 1596.880 ;
        RECT 2906.300 1596.400 2914.100 1596.880 ;
        RECT 5.520 1590.960 13.700 1591.440 ;
        RECT 2906.300 1590.960 2914.100 1591.440 ;
        RECT 5.520 1585.520 13.700 1586.000 ;
        RECT 2906.300 1585.520 2914.100 1586.000 ;
        RECT 5.520 1580.080 13.700 1580.560 ;
        RECT 2906.300 1580.080 2914.100 1580.560 ;
        RECT 5.520 1574.640 13.700 1575.120 ;
        RECT 2906.300 1574.640 2914.100 1575.120 ;
        RECT 5.520 1569.200 13.700 1569.680 ;
        RECT 2906.300 1569.200 2914.100 1569.680 ;
        RECT 5.520 1563.760 13.700 1564.240 ;
        RECT 2906.300 1563.760 2914.100 1564.240 ;
        RECT 5.520 1558.320 13.700 1558.800 ;
        RECT 2906.300 1558.320 2914.100 1558.800 ;
        RECT 5.520 1552.880 13.700 1553.360 ;
        RECT 2906.300 1552.880 2914.100 1553.360 ;
        RECT 5.520 1547.440 13.700 1547.920 ;
        RECT 2906.300 1547.440 2914.100 1547.920 ;
        RECT 5.520 1542.000 13.700 1542.480 ;
        RECT 2906.300 1542.000 2914.100 1542.480 ;
        RECT 5.520 1536.560 13.700 1537.040 ;
        RECT 2906.300 1536.560 2914.100 1537.040 ;
        RECT 5.520 1531.120 13.700 1531.600 ;
        RECT 2906.300 1531.120 2914.100 1531.600 ;
        RECT 5.520 1525.680 13.700 1526.160 ;
        RECT 2906.300 1525.680 2914.100 1526.160 ;
        RECT 5.520 1520.240 13.700 1520.720 ;
        RECT 2906.300 1520.240 2914.100 1520.720 ;
        RECT 5.520 1514.800 13.700 1515.280 ;
        RECT 2906.300 1514.800 2914.100 1515.280 ;
        RECT 5.520 1509.360 13.700 1509.840 ;
        RECT 2906.300 1509.360 2914.100 1509.840 ;
        RECT 5.520 1503.920 13.700 1504.400 ;
        RECT 2906.300 1503.920 2914.100 1504.400 ;
        RECT 5.520 1498.480 13.700 1498.960 ;
        RECT 2906.300 1498.480 2914.100 1498.960 ;
        RECT 5.520 1493.040 13.700 1493.520 ;
        RECT 2906.300 1493.040 2914.100 1493.520 ;
        RECT 5.520 1487.600 13.700 1488.080 ;
        RECT 2906.300 1487.600 2914.100 1488.080 ;
        RECT 5.520 1482.160 13.700 1482.640 ;
        RECT 2906.300 1482.160 2914.100 1482.640 ;
        RECT 5.520 1476.720 13.700 1477.200 ;
        RECT 2906.300 1476.720 2914.100 1477.200 ;
        RECT 5.520 1471.280 13.700 1471.760 ;
        RECT 2906.300 1471.280 2914.100 1471.760 ;
        RECT 5.520 1465.840 13.700 1466.320 ;
        RECT 2906.300 1465.840 2914.100 1466.320 ;
        RECT 5.520 1460.400 13.700 1460.880 ;
        RECT 2906.300 1460.400 2914.100 1460.880 ;
        RECT 5.520 1454.960 13.700 1455.440 ;
        RECT 2906.300 1454.960 2914.100 1455.440 ;
        RECT 5.520 1449.520 13.700 1450.000 ;
        RECT 2906.300 1449.520 2914.100 1450.000 ;
        RECT 5.520 1444.080 13.700 1444.560 ;
        RECT 2906.300 1444.080 2914.100 1444.560 ;
        RECT 5.520 1438.640 13.700 1439.120 ;
        RECT 2906.300 1438.640 2914.100 1439.120 ;
        RECT 5.520 1433.200 13.700 1433.680 ;
        RECT 2906.300 1433.200 2914.100 1433.680 ;
        RECT 5.520 1427.760 13.700 1428.240 ;
        RECT 2906.300 1427.760 2914.100 1428.240 ;
        RECT 5.520 1422.320 13.700 1422.800 ;
        RECT 2906.300 1422.320 2914.100 1422.800 ;
        RECT 5.520 1416.880 13.700 1417.360 ;
        RECT 2906.300 1416.880 2914.100 1417.360 ;
        RECT 5.520 1411.440 13.700 1411.920 ;
        RECT 2906.300 1411.440 2914.100 1411.920 ;
        RECT 5.520 1406.000 13.700 1406.480 ;
        RECT 2906.300 1406.000 2914.100 1406.480 ;
        RECT 5.520 1400.560 13.700 1401.040 ;
        RECT 2906.300 1400.560 2914.100 1401.040 ;
        RECT 5.520 1395.120 13.700 1395.600 ;
        RECT 2906.300 1395.120 2914.100 1395.600 ;
        RECT 5.520 1389.680 13.700 1390.160 ;
        RECT 2906.300 1389.680 2914.100 1390.160 ;
        RECT 5.520 1384.240 13.700 1384.720 ;
        RECT 2906.300 1384.240 2914.100 1384.720 ;
        RECT 5.520 1378.800 13.700 1379.280 ;
        RECT 2906.300 1378.800 2914.100 1379.280 ;
        RECT 5.520 1373.360 13.700 1373.840 ;
        RECT 2906.300 1373.360 2914.100 1373.840 ;
        RECT 5.520 1367.920 13.700 1368.400 ;
        RECT 2906.300 1367.920 2914.100 1368.400 ;
        RECT 5.520 1362.480 13.700 1362.960 ;
        RECT 2906.300 1362.480 2914.100 1362.960 ;
        RECT 5.520 1357.040 13.700 1357.520 ;
        RECT 2906.300 1357.040 2914.100 1357.520 ;
        RECT 5.520 1351.600 13.700 1352.080 ;
        RECT 2906.300 1351.600 2914.100 1352.080 ;
        RECT 5.520 1346.160 13.700 1346.640 ;
        RECT 2906.300 1346.160 2914.100 1346.640 ;
        RECT 5.520 1340.720 13.700 1341.200 ;
        RECT 2906.300 1340.720 2914.100 1341.200 ;
        RECT 5.520 1335.280 13.700 1335.760 ;
        RECT 2906.300 1335.280 2914.100 1335.760 ;
        RECT 5.520 1329.840 13.700 1330.320 ;
        RECT 2906.300 1329.840 2914.100 1330.320 ;
        RECT 5.520 1324.400 13.700 1324.880 ;
        RECT 2906.300 1324.400 2914.100 1324.880 ;
        RECT 5.520 1318.960 13.700 1319.440 ;
        RECT 2906.300 1318.960 2914.100 1319.440 ;
        RECT 5.520 1313.520 13.700 1314.000 ;
        RECT 2906.300 1313.520 2914.100 1314.000 ;
        RECT 5.520 1308.080 13.700 1308.560 ;
        RECT 2906.300 1308.080 2914.100 1308.560 ;
        RECT 5.520 1302.640 13.700 1303.120 ;
        RECT 2906.300 1302.640 2914.100 1303.120 ;
        RECT 5.520 1297.200 13.700 1297.680 ;
        RECT 2906.300 1297.200 2914.100 1297.680 ;
        RECT 5.520 1291.760 13.700 1292.240 ;
        RECT 2906.300 1291.760 2914.100 1292.240 ;
        RECT 5.520 1286.320 13.700 1286.800 ;
        RECT 2906.300 1286.320 2914.100 1286.800 ;
        RECT 5.520 1280.880 13.700 1281.360 ;
        RECT 2906.300 1280.880 2914.100 1281.360 ;
        RECT 5.520 1275.440 13.700 1275.920 ;
        RECT 2906.300 1275.440 2914.100 1275.920 ;
        RECT 5.520 1270.000 13.700 1270.480 ;
        RECT 2906.300 1270.000 2914.100 1270.480 ;
        RECT 5.520 1264.560 13.700 1265.040 ;
        RECT 2906.300 1264.560 2914.100 1265.040 ;
        RECT 5.520 1259.120 13.700 1259.600 ;
        RECT 2906.300 1259.120 2914.100 1259.600 ;
        RECT 5.520 1253.680 13.700 1254.160 ;
        RECT 2906.300 1253.680 2914.100 1254.160 ;
        RECT 5.520 1248.240 13.700 1248.720 ;
        RECT 2906.300 1248.240 2914.100 1248.720 ;
        RECT 5.520 1242.800 13.700 1243.280 ;
        RECT 2906.300 1242.800 2914.100 1243.280 ;
        RECT 5.520 1237.360 13.700 1237.840 ;
        RECT 2906.300 1237.360 2914.100 1237.840 ;
        RECT 5.520 1231.920 13.700 1232.400 ;
        RECT 2906.300 1231.920 2914.100 1232.400 ;
        RECT 5.520 1226.480 13.700 1226.960 ;
        RECT 2906.300 1226.480 2914.100 1226.960 ;
        RECT 5.520 1221.040 13.700 1221.520 ;
        RECT 2906.300 1221.040 2914.100 1221.520 ;
        RECT 5.520 1215.600 13.700 1216.080 ;
        RECT 2906.300 1215.600 2914.100 1216.080 ;
        RECT 5.520 1210.160 13.700 1210.640 ;
        RECT 2906.300 1210.160 2914.100 1210.640 ;
        RECT 5.520 1204.720 13.700 1205.200 ;
        RECT 2906.300 1204.720 2914.100 1205.200 ;
        RECT 5.520 1199.280 13.700 1199.760 ;
        RECT 2906.300 1199.280 2914.100 1199.760 ;
        RECT 5.520 1193.840 13.700 1194.320 ;
        RECT 2906.300 1193.840 2914.100 1194.320 ;
        RECT 5.520 1188.400 13.700 1188.880 ;
        RECT 2906.300 1188.400 2914.100 1188.880 ;
        RECT 5.520 1182.960 13.700 1183.440 ;
        RECT 2906.300 1182.960 2914.100 1183.440 ;
        RECT 5.520 1177.520 13.700 1178.000 ;
        RECT 2906.300 1177.520 2914.100 1178.000 ;
        RECT 5.520 1172.080 13.700 1172.560 ;
        RECT 2906.300 1172.080 2914.100 1172.560 ;
        RECT 5.520 1166.640 13.700 1167.120 ;
        RECT 2906.300 1166.640 2914.100 1167.120 ;
        RECT 5.520 1161.200 13.700 1161.680 ;
        RECT 2906.300 1161.200 2914.100 1161.680 ;
        RECT 5.520 1155.760 13.700 1156.240 ;
        RECT 2906.300 1155.760 2914.100 1156.240 ;
        RECT 5.520 1150.320 13.700 1150.800 ;
        RECT 2906.300 1150.320 2914.100 1150.800 ;
        RECT 5.520 1144.880 13.700 1145.360 ;
        RECT 2906.300 1144.880 2914.100 1145.360 ;
        RECT 5.520 1139.440 13.700 1139.920 ;
        RECT 2906.300 1139.440 2914.100 1139.920 ;
        RECT 5.520 1134.000 13.700 1134.480 ;
        RECT 2906.300 1134.000 2914.100 1134.480 ;
        RECT 5.520 1128.560 13.700 1129.040 ;
        RECT 2906.300 1128.560 2914.100 1129.040 ;
        RECT 5.520 1123.120 13.700 1123.600 ;
        RECT 2906.300 1123.120 2914.100 1123.600 ;
        RECT 5.520 1117.680 13.700 1118.160 ;
        RECT 2906.300 1117.680 2914.100 1118.160 ;
        RECT 5.520 1112.240 13.700 1112.720 ;
        RECT 2906.300 1112.240 2914.100 1112.720 ;
        RECT 5.520 1106.800 13.700 1107.280 ;
        RECT 2906.300 1106.800 2914.100 1107.280 ;
        RECT 5.520 1101.360 13.700 1101.840 ;
        RECT 2906.300 1101.360 2914.100 1101.840 ;
        RECT 5.520 1095.920 13.700 1096.400 ;
        RECT 2906.300 1095.920 2914.100 1096.400 ;
        RECT 5.520 1090.480 13.700 1090.960 ;
        RECT 2906.300 1090.480 2914.100 1090.960 ;
        RECT 5.520 1085.040 13.700 1085.520 ;
        RECT 2906.300 1085.040 2914.100 1085.520 ;
        RECT 5.520 1079.600 13.700 1080.080 ;
        RECT 2906.300 1079.600 2914.100 1080.080 ;
        RECT 5.520 1074.160 13.700 1074.640 ;
        RECT 2906.300 1074.160 2914.100 1074.640 ;
        RECT 5.520 1068.720 13.700 1069.200 ;
        RECT 2906.300 1068.720 2914.100 1069.200 ;
        RECT 5.520 1063.280 13.700 1063.760 ;
        RECT 2906.300 1063.280 2914.100 1063.760 ;
        RECT 5.520 1057.840 13.700 1058.320 ;
        RECT 2906.300 1057.840 2914.100 1058.320 ;
        RECT 5.520 1052.400 13.700 1052.880 ;
        RECT 2906.300 1052.400 2914.100 1052.880 ;
        RECT 5.520 1046.960 13.700 1047.440 ;
        RECT 2906.300 1046.960 2914.100 1047.440 ;
        RECT 5.520 1041.520 13.700 1042.000 ;
        RECT 2906.300 1041.520 2914.100 1042.000 ;
        RECT 5.520 1036.080 13.700 1036.560 ;
        RECT 2906.300 1036.080 2914.100 1036.560 ;
        RECT 5.520 1030.640 13.700 1031.120 ;
        RECT 2906.300 1030.640 2914.100 1031.120 ;
        RECT 5.520 1025.200 13.700 1025.680 ;
        RECT 2906.300 1025.200 2914.100 1025.680 ;
        RECT 5.520 1019.760 13.700 1020.240 ;
        RECT 2906.300 1019.760 2914.100 1020.240 ;
        RECT 5.520 1014.320 13.700 1014.800 ;
        RECT 2906.300 1014.320 2914.100 1014.800 ;
        RECT 5.520 1008.880 13.700 1009.360 ;
        RECT 2906.300 1008.880 2914.100 1009.360 ;
        RECT 5.520 1003.440 13.700 1003.920 ;
        RECT 2906.300 1003.440 2914.100 1003.920 ;
        RECT 5.520 998.000 13.700 998.480 ;
        RECT 2906.300 998.000 2914.100 998.480 ;
        RECT 5.520 992.560 13.700 993.040 ;
        RECT 2906.300 992.560 2914.100 993.040 ;
        RECT 5.520 987.120 13.700 987.600 ;
        RECT 2906.300 987.120 2914.100 987.600 ;
        RECT 5.520 981.680 13.700 982.160 ;
        RECT 2906.300 981.680 2914.100 982.160 ;
        RECT 5.520 976.240 13.700 976.720 ;
        RECT 2906.300 976.240 2914.100 976.720 ;
        RECT 5.520 970.800 13.700 971.280 ;
        RECT 2906.300 970.800 2914.100 971.280 ;
        RECT 5.520 965.360 13.700 965.840 ;
        RECT 2906.300 965.360 2914.100 965.840 ;
        RECT 5.520 959.920 13.700 960.400 ;
        RECT 2906.300 959.920 2914.100 960.400 ;
        RECT 5.520 954.480 13.700 954.960 ;
        RECT 2906.300 954.480 2914.100 954.960 ;
        RECT 5.520 949.040 13.700 949.520 ;
        RECT 2906.300 949.040 2914.100 949.520 ;
        RECT 5.520 943.600 13.700 944.080 ;
        RECT 2906.300 943.600 2914.100 944.080 ;
        RECT 5.520 938.160 13.700 938.640 ;
        RECT 2906.300 938.160 2914.100 938.640 ;
        RECT 5.520 932.720 13.700 933.200 ;
        RECT 2906.300 932.720 2914.100 933.200 ;
        RECT 5.520 927.280 13.700 927.760 ;
        RECT 2906.300 927.280 2914.100 927.760 ;
        RECT 5.520 921.840 13.700 922.320 ;
        RECT 2906.300 921.840 2914.100 922.320 ;
        RECT 5.520 916.400 13.700 916.880 ;
        RECT 2906.300 916.400 2914.100 916.880 ;
        RECT 5.520 910.960 13.700 911.440 ;
        RECT 2906.300 910.960 2914.100 911.440 ;
        RECT 5.520 905.520 13.700 906.000 ;
        RECT 2906.300 905.520 2914.100 906.000 ;
        RECT 5.520 900.080 13.700 900.560 ;
        RECT 2906.300 900.080 2914.100 900.560 ;
        RECT 5.520 894.640 13.700 895.120 ;
        RECT 2906.300 894.640 2914.100 895.120 ;
        RECT 5.520 889.200 13.700 889.680 ;
        RECT 2906.300 889.200 2914.100 889.680 ;
        RECT 5.520 883.760 13.700 884.240 ;
        RECT 2906.300 883.760 2914.100 884.240 ;
        RECT 5.520 878.320 13.700 878.800 ;
        RECT 2906.300 878.320 2914.100 878.800 ;
        RECT 5.520 872.880 13.700 873.360 ;
        RECT 2906.300 872.880 2914.100 873.360 ;
        RECT 5.520 867.440 13.700 867.920 ;
        RECT 2906.300 867.440 2914.100 867.920 ;
        RECT 5.520 862.000 13.700 862.480 ;
        RECT 2906.300 862.000 2914.100 862.480 ;
        RECT 5.520 856.560 13.700 857.040 ;
        RECT 2906.300 856.560 2914.100 857.040 ;
        RECT 5.520 851.120 13.700 851.600 ;
        RECT 2906.300 851.120 2914.100 851.600 ;
        RECT 5.520 845.680 13.700 846.160 ;
        RECT 2906.300 845.680 2914.100 846.160 ;
        RECT 5.520 840.240 13.700 840.720 ;
        RECT 2906.300 840.240 2914.100 840.720 ;
        RECT 5.520 834.800 13.700 835.280 ;
        RECT 2906.300 834.800 2914.100 835.280 ;
        RECT 5.520 829.360 13.700 829.840 ;
        RECT 2906.300 829.360 2914.100 829.840 ;
        RECT 5.520 823.920 13.700 824.400 ;
        RECT 2906.300 823.920 2914.100 824.400 ;
        RECT 5.520 818.480 13.700 818.960 ;
        RECT 2906.300 818.480 2914.100 818.960 ;
        RECT 5.520 813.040 13.700 813.520 ;
        RECT 2906.300 813.040 2914.100 813.520 ;
        RECT 5.520 807.600 13.700 808.080 ;
        RECT 2906.300 807.600 2914.100 808.080 ;
        RECT 5.520 802.160 13.700 802.640 ;
        RECT 2906.300 802.160 2914.100 802.640 ;
        RECT 5.520 796.720 13.700 797.200 ;
        RECT 2906.300 796.720 2914.100 797.200 ;
        RECT 5.520 791.280 13.700 791.760 ;
        RECT 2906.300 791.280 2914.100 791.760 ;
        RECT 5.520 785.840 13.700 786.320 ;
        RECT 2906.300 785.840 2914.100 786.320 ;
        RECT 5.520 780.400 13.700 780.880 ;
        RECT 2906.300 780.400 2914.100 780.880 ;
        RECT 5.520 774.960 13.700 775.440 ;
        RECT 2906.300 774.960 2914.100 775.440 ;
        RECT 5.520 769.520 13.700 770.000 ;
        RECT 2906.300 769.520 2914.100 770.000 ;
        RECT 5.520 764.080 13.700 764.560 ;
        RECT 2906.300 764.080 2914.100 764.560 ;
        RECT 5.520 758.640 13.700 759.120 ;
        RECT 2906.300 758.640 2914.100 759.120 ;
        RECT 5.520 753.200 13.700 753.680 ;
        RECT 2906.300 753.200 2914.100 753.680 ;
        RECT 5.520 747.760 13.700 748.240 ;
        RECT 2906.300 747.760 2914.100 748.240 ;
        RECT 5.520 742.320 13.700 742.800 ;
        RECT 2906.300 742.320 2914.100 742.800 ;
        RECT 5.520 736.880 13.700 737.360 ;
        RECT 2906.300 736.880 2914.100 737.360 ;
        RECT 5.520 731.440 13.700 731.920 ;
        RECT 2906.300 731.440 2914.100 731.920 ;
        RECT 5.520 726.000 13.700 726.480 ;
        RECT 2906.300 726.000 2914.100 726.480 ;
        RECT 5.520 720.560 13.700 721.040 ;
        RECT 2906.300 720.560 2914.100 721.040 ;
        RECT 5.520 715.120 13.700 715.600 ;
        RECT 2906.300 715.120 2914.100 715.600 ;
        RECT 5.520 709.680 13.700 710.160 ;
        RECT 2906.300 709.680 2914.100 710.160 ;
        RECT 5.520 704.240 13.700 704.720 ;
        RECT 2906.300 704.240 2914.100 704.720 ;
        RECT 5.520 698.800 13.700 699.280 ;
        RECT 2906.300 698.800 2914.100 699.280 ;
        RECT 5.520 693.360 13.700 693.840 ;
        RECT 2906.300 693.360 2914.100 693.840 ;
        RECT 5.520 687.920 13.700 688.400 ;
        RECT 2906.300 687.920 2914.100 688.400 ;
        RECT 5.520 682.480 13.700 682.960 ;
        RECT 2906.300 682.480 2914.100 682.960 ;
        RECT 5.520 677.040 13.700 677.520 ;
        RECT 2906.300 677.040 2914.100 677.520 ;
        RECT 5.520 671.600 13.700 672.080 ;
        RECT 2906.300 671.600 2914.100 672.080 ;
        RECT 5.520 666.160 13.700 666.640 ;
        RECT 2906.300 666.160 2914.100 666.640 ;
        RECT 5.520 660.720 13.700 661.200 ;
        RECT 2906.300 660.720 2914.100 661.200 ;
        RECT 5.520 655.280 13.700 655.760 ;
        RECT 2906.300 655.280 2914.100 655.760 ;
        RECT 5.520 649.840 13.700 650.320 ;
        RECT 2906.300 649.840 2914.100 650.320 ;
        RECT 5.520 644.400 13.700 644.880 ;
        RECT 2906.300 644.400 2914.100 644.880 ;
        RECT 5.520 638.960 13.700 639.440 ;
        RECT 2906.300 638.960 2914.100 639.440 ;
        RECT 5.520 633.520 13.700 634.000 ;
        RECT 2906.300 633.520 2914.100 634.000 ;
        RECT 5.520 628.080 13.700 628.560 ;
        RECT 2906.300 628.080 2914.100 628.560 ;
        RECT 5.520 622.640 13.700 623.120 ;
        RECT 2906.300 622.640 2914.100 623.120 ;
        RECT 5.520 617.200 13.700 617.680 ;
        RECT 2906.300 617.200 2914.100 617.680 ;
        RECT 5.520 611.760 13.700 612.240 ;
        RECT 2906.300 611.760 2914.100 612.240 ;
        RECT 5.520 606.320 13.700 606.800 ;
        RECT 2906.300 606.320 2914.100 606.800 ;
        RECT 5.520 600.880 13.700 601.360 ;
        RECT 2906.300 600.880 2914.100 601.360 ;
        RECT 5.520 595.440 13.700 595.920 ;
        RECT 2906.300 595.440 2914.100 595.920 ;
        RECT 5.520 590.000 13.700 590.480 ;
        RECT 2906.300 590.000 2914.100 590.480 ;
        RECT 5.520 584.560 13.700 585.040 ;
        RECT 2906.300 584.560 2914.100 585.040 ;
        RECT 5.520 579.120 13.700 579.600 ;
        RECT 2906.300 579.120 2914.100 579.600 ;
        RECT 5.520 573.680 13.700 574.160 ;
        RECT 2906.300 573.680 2914.100 574.160 ;
        RECT 5.520 568.240 13.700 568.720 ;
        RECT 2906.300 568.240 2914.100 568.720 ;
        RECT 5.520 562.800 13.700 563.280 ;
        RECT 2906.300 562.800 2914.100 563.280 ;
        RECT 5.520 557.360 13.700 557.840 ;
        RECT 2906.300 557.360 2914.100 557.840 ;
        RECT 5.520 551.920 13.700 552.400 ;
        RECT 2906.300 551.920 2914.100 552.400 ;
        RECT 5.520 546.480 13.700 546.960 ;
        RECT 2906.300 546.480 2914.100 546.960 ;
        RECT 5.520 541.040 13.700 541.520 ;
        RECT 2906.300 541.040 2914.100 541.520 ;
        RECT 5.520 535.600 13.700 536.080 ;
        RECT 2906.300 535.600 2914.100 536.080 ;
        RECT 5.520 530.160 13.700 530.640 ;
        RECT 2906.300 530.160 2914.100 530.640 ;
        RECT 5.520 524.720 13.700 525.200 ;
        RECT 2906.300 524.720 2914.100 525.200 ;
        RECT 5.520 519.280 13.700 519.760 ;
        RECT 2906.300 519.280 2914.100 519.760 ;
        RECT 5.520 513.840 13.700 514.320 ;
        RECT 2906.300 513.840 2914.100 514.320 ;
        RECT 5.520 508.400 13.700 508.880 ;
        RECT 2906.300 508.400 2914.100 508.880 ;
        RECT 5.520 502.960 13.700 503.440 ;
        RECT 2906.300 502.960 2914.100 503.440 ;
        RECT 5.520 497.520 13.700 498.000 ;
        RECT 2906.300 497.520 2914.100 498.000 ;
        RECT 5.520 492.080 13.700 492.560 ;
        RECT 2906.300 492.080 2914.100 492.560 ;
        RECT 5.520 486.640 13.700 487.120 ;
        RECT 2906.300 486.640 2914.100 487.120 ;
        RECT 5.520 481.200 13.700 481.680 ;
        RECT 2906.300 481.200 2914.100 481.680 ;
        RECT 5.520 475.760 13.700 476.240 ;
        RECT 2906.300 475.760 2914.100 476.240 ;
        RECT 5.520 470.320 13.700 470.800 ;
        RECT 2906.300 470.320 2914.100 470.800 ;
        RECT 5.520 464.880 13.700 465.360 ;
        RECT 2906.300 464.880 2914.100 465.360 ;
        RECT 5.520 459.440 13.700 459.920 ;
        RECT 2906.300 459.440 2914.100 459.920 ;
        RECT 5.520 454.000 13.700 454.480 ;
        RECT 2906.300 454.000 2914.100 454.480 ;
        RECT 5.520 448.560 13.700 449.040 ;
        RECT 2906.300 448.560 2914.100 449.040 ;
        RECT 5.520 443.120 13.700 443.600 ;
        RECT 2906.300 443.120 2914.100 443.600 ;
        RECT 5.520 437.680 13.700 438.160 ;
        RECT 2906.300 437.680 2914.100 438.160 ;
        RECT 5.520 432.240 13.700 432.720 ;
        RECT 2906.300 432.240 2914.100 432.720 ;
        RECT 5.520 426.800 13.700 427.280 ;
        RECT 2906.300 426.800 2914.100 427.280 ;
        RECT 5.520 421.360 13.700 421.840 ;
        RECT 2906.300 421.360 2914.100 421.840 ;
        RECT 5.520 415.920 13.700 416.400 ;
        RECT 2906.300 415.920 2914.100 416.400 ;
        RECT 5.520 410.480 13.700 410.960 ;
        RECT 2906.300 410.480 2914.100 410.960 ;
        RECT 5.520 405.040 13.700 405.520 ;
        RECT 2906.300 405.040 2914.100 405.520 ;
        RECT 5.520 399.600 13.700 400.080 ;
        RECT 2906.300 399.600 2914.100 400.080 ;
        RECT 5.520 394.160 13.700 394.640 ;
        RECT 2906.300 394.160 2914.100 394.640 ;
        RECT 5.520 388.720 13.700 389.200 ;
        RECT 2906.300 388.720 2914.100 389.200 ;
        RECT 5.520 383.280 13.700 383.760 ;
        RECT 2906.300 383.280 2914.100 383.760 ;
        RECT 5.520 377.840 13.700 378.320 ;
        RECT 2906.300 377.840 2914.100 378.320 ;
        RECT 5.520 372.400 13.700 372.880 ;
        RECT 2906.300 372.400 2914.100 372.880 ;
        RECT 5.520 366.960 13.700 367.440 ;
        RECT 2906.300 366.960 2914.100 367.440 ;
        RECT 5.520 361.520 13.700 362.000 ;
        RECT 2906.300 361.520 2914.100 362.000 ;
        RECT 5.520 356.080 13.700 356.560 ;
        RECT 2906.300 356.080 2914.100 356.560 ;
        RECT 5.520 350.640 13.700 351.120 ;
        RECT 2906.300 350.640 2914.100 351.120 ;
        RECT 5.520 345.200 13.700 345.680 ;
        RECT 2906.300 345.200 2914.100 345.680 ;
        RECT 5.520 339.760 13.700 340.240 ;
        RECT 2906.300 339.760 2914.100 340.240 ;
        RECT 5.520 334.320 13.700 334.800 ;
        RECT 2906.300 334.320 2914.100 334.800 ;
        RECT 5.520 328.880 13.700 329.360 ;
        RECT 2906.300 328.880 2914.100 329.360 ;
        RECT 5.520 323.440 13.700 323.920 ;
        RECT 2906.300 323.440 2914.100 323.920 ;
        RECT 5.520 318.000 13.700 318.480 ;
        RECT 2906.300 318.000 2914.100 318.480 ;
        RECT 5.520 312.560 13.700 313.040 ;
        RECT 2906.300 312.560 2914.100 313.040 ;
        RECT 5.520 307.120 13.700 307.600 ;
        RECT 2906.300 307.120 2914.100 307.600 ;
        RECT 5.520 301.680 13.700 302.160 ;
        RECT 2906.300 301.680 2914.100 302.160 ;
        RECT 5.520 296.240 13.700 296.720 ;
        RECT 2906.300 296.240 2914.100 296.720 ;
        RECT 5.520 290.800 13.700 291.280 ;
        RECT 2906.300 290.800 2914.100 291.280 ;
        RECT 5.520 285.360 13.700 285.840 ;
        RECT 2906.300 285.360 2914.100 285.840 ;
        RECT 5.520 279.920 13.700 280.400 ;
        RECT 2906.300 279.920 2914.100 280.400 ;
        RECT 5.520 274.480 13.700 274.960 ;
        RECT 2906.300 274.480 2914.100 274.960 ;
        RECT 5.520 269.040 13.700 269.520 ;
        RECT 2906.300 269.040 2914.100 269.520 ;
        RECT 5.520 263.600 13.700 264.080 ;
        RECT 2906.300 263.600 2914.100 264.080 ;
        RECT 5.520 258.160 13.700 258.640 ;
        RECT 2906.300 258.160 2914.100 258.640 ;
        RECT 5.520 252.720 13.700 253.200 ;
        RECT 2906.300 252.720 2914.100 253.200 ;
        RECT 5.520 247.280 13.700 247.760 ;
        RECT 2906.300 247.280 2914.100 247.760 ;
        RECT 5.520 241.840 13.700 242.320 ;
        RECT 2906.300 241.840 2914.100 242.320 ;
        RECT 5.520 236.400 13.700 236.880 ;
        RECT 2906.300 236.400 2914.100 236.880 ;
        RECT 5.520 230.960 13.700 231.440 ;
        RECT 2906.300 230.960 2914.100 231.440 ;
        RECT 5.520 225.520 13.700 226.000 ;
        RECT 2906.300 225.520 2914.100 226.000 ;
        RECT 5.520 220.080 13.700 220.560 ;
        RECT 2906.300 220.080 2914.100 220.560 ;
        RECT 5.520 214.640 13.700 215.120 ;
        RECT 2906.300 214.640 2914.100 215.120 ;
        RECT 5.520 209.200 13.700 209.680 ;
        RECT 2906.300 209.200 2914.100 209.680 ;
        RECT 5.520 203.760 13.700 204.240 ;
        RECT 2906.300 203.760 2914.100 204.240 ;
        RECT 5.520 198.320 13.700 198.800 ;
        RECT 2906.300 198.320 2914.100 198.800 ;
        RECT 5.520 192.880 13.700 193.360 ;
        RECT 2906.300 192.880 2914.100 193.360 ;
        RECT 5.520 187.440 13.700 187.920 ;
        RECT 2906.300 187.440 2914.100 187.920 ;
        RECT 5.520 182.000 13.700 182.480 ;
        RECT 2906.300 182.000 2914.100 182.480 ;
        RECT 5.520 176.560 13.700 177.040 ;
        RECT 2906.300 176.560 2914.100 177.040 ;
        RECT 5.520 171.120 13.700 171.600 ;
        RECT 2906.300 171.120 2914.100 171.600 ;
        RECT 5.520 165.680 13.700 166.160 ;
        RECT 2906.300 165.680 2914.100 166.160 ;
        RECT 5.520 160.240 13.700 160.720 ;
        RECT 2906.300 160.240 2914.100 160.720 ;
        RECT 5.520 154.800 13.700 155.280 ;
        RECT 2906.300 154.800 2914.100 155.280 ;
        RECT 5.520 149.360 13.700 149.840 ;
        RECT 2906.300 149.360 2914.100 149.840 ;
        RECT 5.520 143.920 13.700 144.400 ;
        RECT 2906.300 143.920 2914.100 144.400 ;
        RECT 5.520 138.480 13.700 138.960 ;
        RECT 2906.300 138.480 2914.100 138.960 ;
        RECT 5.520 133.040 13.700 133.520 ;
        RECT 2906.300 133.040 2914.100 133.520 ;
        RECT 5.520 127.600 13.700 128.080 ;
        RECT 2906.300 127.600 2914.100 128.080 ;
        RECT 5.520 122.160 13.700 122.640 ;
        RECT 2906.300 122.160 2914.100 122.640 ;
        RECT 5.520 116.720 13.700 117.200 ;
        RECT 2906.300 116.720 2914.100 117.200 ;
        RECT 5.520 111.280 13.700 111.760 ;
        RECT 2906.300 111.280 2914.100 111.760 ;
        RECT 5.520 105.840 13.700 106.320 ;
        RECT 2906.300 105.840 2914.100 106.320 ;
        RECT 5.520 100.400 13.700 100.880 ;
        RECT 2906.300 100.400 2914.100 100.880 ;
        RECT 5.520 94.960 13.700 95.440 ;
        RECT 2906.300 94.960 2914.100 95.440 ;
        RECT 5.520 89.520 13.700 90.000 ;
        RECT 2906.300 89.520 2914.100 90.000 ;
        RECT 5.520 84.080 13.700 84.560 ;
        RECT 2906.300 84.080 2914.100 84.560 ;
        RECT 5.520 78.640 13.700 79.120 ;
        RECT 2906.300 78.640 2914.100 79.120 ;
        RECT 5.520 73.200 13.700 73.680 ;
        RECT 2906.300 73.200 2914.100 73.680 ;
        RECT 5.520 67.760 13.700 68.240 ;
        RECT 2906.300 67.760 2914.100 68.240 ;
        RECT 5.520 62.320 13.700 62.800 ;
        RECT 2906.300 62.320 2914.100 62.800 ;
        RECT 5.520 56.880 13.700 57.360 ;
        RECT 2906.300 56.880 2914.100 57.360 ;
        RECT 5.520 51.440 13.700 51.920 ;
        RECT 2906.300 51.440 2914.100 51.920 ;
        RECT 5.520 46.000 13.700 46.480 ;
        RECT 2906.300 46.000 2914.100 46.480 ;
        RECT 5.520 40.560 13.700 41.040 ;
        RECT 2906.300 40.560 2914.100 41.040 ;
        RECT 5.520 35.120 13.700 35.600 ;
        RECT 2906.300 35.120 2914.100 35.600 ;
        RECT 5.520 29.680 13.700 30.160 ;
        RECT 2906.300 29.680 2914.100 30.160 ;
        RECT 5.520 24.240 13.700 24.720 ;
        RECT 2906.300 24.240 2914.100 24.720 ;
        RECT 5.520 18.800 13.700 19.280 ;
        RECT 2906.300 18.800 2914.100 19.280 ;
        RECT 5.520 13.700 13.700 13.840 ;
        RECT 2906.300 13.700 2914.100 13.840 ;
        RECT 5.520 13.360 2914.100 13.700 ;
      LAYER via ;
        RECT 49.110 13.470 49.370 13.700 ;
        RECT 49.430 13.470 49.690 13.700 ;
        RECT 49.750 13.470 50.010 13.700 ;
        RECT 50.070 13.470 50.330 13.700 ;
        RECT 50.390 13.470 50.650 13.700 ;
        RECT 50.710 13.470 50.970 13.700 ;
        RECT 51.030 13.470 51.290 13.700 ;
        RECT 51.350 13.470 51.610 13.700 ;
        RECT 51.670 13.470 51.930 13.700 ;
        RECT 139.110 13.470 139.370 13.700 ;
        RECT 139.430 13.470 139.690 13.700 ;
        RECT 139.750 13.470 140.010 13.700 ;
        RECT 140.070 13.470 140.330 13.700 ;
        RECT 140.390 13.470 140.650 13.700 ;
        RECT 140.710 13.470 140.970 13.700 ;
        RECT 141.030 13.470 141.290 13.700 ;
        RECT 141.350 13.470 141.610 13.700 ;
        RECT 141.670 13.470 141.930 13.700 ;
        RECT 229.110 13.470 229.370 13.700 ;
        RECT 229.430 13.470 229.690 13.700 ;
        RECT 229.750 13.470 230.010 13.700 ;
        RECT 230.070 13.470 230.330 13.700 ;
        RECT 230.390 13.470 230.650 13.700 ;
        RECT 230.710 13.470 230.970 13.700 ;
        RECT 231.030 13.470 231.290 13.700 ;
        RECT 231.350 13.470 231.610 13.700 ;
        RECT 231.670 13.470 231.930 13.700 ;
        RECT 319.110 13.470 319.370 13.700 ;
        RECT 319.430 13.470 319.690 13.700 ;
        RECT 319.750 13.470 320.010 13.700 ;
        RECT 320.070 13.470 320.330 13.700 ;
        RECT 320.390 13.470 320.650 13.700 ;
        RECT 320.710 13.470 320.970 13.700 ;
        RECT 321.030 13.470 321.290 13.700 ;
        RECT 321.350 13.470 321.610 13.700 ;
        RECT 321.670 13.470 321.930 13.700 ;
        RECT 409.110 13.470 409.370 13.700 ;
        RECT 409.430 13.470 409.690 13.700 ;
        RECT 409.750 13.470 410.010 13.700 ;
        RECT 410.070 13.470 410.330 13.700 ;
        RECT 410.390 13.470 410.650 13.700 ;
        RECT 410.710 13.470 410.970 13.700 ;
        RECT 411.030 13.470 411.290 13.700 ;
        RECT 411.350 13.470 411.610 13.700 ;
        RECT 411.670 13.470 411.930 13.700 ;
        RECT 499.110 13.470 499.370 13.700 ;
        RECT 499.430 13.470 499.690 13.700 ;
        RECT 499.750 13.470 500.010 13.700 ;
        RECT 500.070 13.470 500.330 13.700 ;
        RECT 500.390 13.470 500.650 13.700 ;
        RECT 500.710 13.470 500.970 13.700 ;
        RECT 501.030 13.470 501.290 13.700 ;
        RECT 501.350 13.470 501.610 13.700 ;
        RECT 501.670 13.470 501.930 13.700 ;
        RECT 589.110 13.470 589.370 13.700 ;
        RECT 589.430 13.470 589.690 13.700 ;
        RECT 589.750 13.470 590.010 13.700 ;
        RECT 590.070 13.470 590.330 13.700 ;
        RECT 590.390 13.470 590.650 13.700 ;
        RECT 590.710 13.470 590.970 13.700 ;
        RECT 591.030 13.470 591.290 13.700 ;
        RECT 591.350 13.470 591.610 13.700 ;
        RECT 591.670 13.470 591.930 13.700 ;
        RECT 679.110 13.470 679.370 13.700 ;
        RECT 679.430 13.470 679.690 13.700 ;
        RECT 679.750 13.470 680.010 13.700 ;
        RECT 680.070 13.470 680.330 13.700 ;
        RECT 680.390 13.470 680.650 13.700 ;
        RECT 680.710 13.470 680.970 13.700 ;
        RECT 681.030 13.470 681.290 13.700 ;
        RECT 681.350 13.470 681.610 13.700 ;
        RECT 681.670 13.470 681.930 13.700 ;
        RECT 769.110 13.470 769.370 13.700 ;
        RECT 769.430 13.470 769.690 13.700 ;
        RECT 769.750 13.470 770.010 13.700 ;
        RECT 770.070 13.470 770.330 13.700 ;
        RECT 770.390 13.470 770.650 13.700 ;
        RECT 770.710 13.470 770.970 13.700 ;
        RECT 771.030 13.470 771.290 13.700 ;
        RECT 771.350 13.470 771.610 13.700 ;
        RECT 771.670 13.470 771.930 13.700 ;
        RECT 859.110 13.470 859.370 13.700 ;
        RECT 859.430 13.470 859.690 13.700 ;
        RECT 859.750 13.470 860.010 13.700 ;
        RECT 860.070 13.470 860.330 13.700 ;
        RECT 860.390 13.470 860.650 13.700 ;
        RECT 860.710 13.470 860.970 13.700 ;
        RECT 861.030 13.470 861.290 13.700 ;
        RECT 861.350 13.470 861.610 13.700 ;
        RECT 861.670 13.470 861.930 13.700 ;
        RECT 949.110 13.470 949.370 13.700 ;
        RECT 949.430 13.470 949.690 13.700 ;
        RECT 949.750 13.470 950.010 13.700 ;
        RECT 950.070 13.470 950.330 13.700 ;
        RECT 950.390 13.470 950.650 13.700 ;
        RECT 950.710 13.470 950.970 13.700 ;
        RECT 951.030 13.470 951.290 13.700 ;
        RECT 951.350 13.470 951.610 13.700 ;
        RECT 951.670 13.470 951.930 13.700 ;
        RECT 1039.110 13.470 1039.370 13.700 ;
        RECT 1039.430 13.470 1039.690 13.700 ;
        RECT 1039.750 13.470 1040.010 13.700 ;
        RECT 1040.070 13.470 1040.330 13.700 ;
        RECT 1040.390 13.470 1040.650 13.700 ;
        RECT 1040.710 13.470 1040.970 13.700 ;
        RECT 1041.030 13.470 1041.290 13.700 ;
        RECT 1041.350 13.470 1041.610 13.700 ;
        RECT 1041.670 13.470 1041.930 13.700 ;
        RECT 1129.110 13.470 1129.370 13.700 ;
        RECT 1129.430 13.470 1129.690 13.700 ;
        RECT 1129.750 13.470 1130.010 13.700 ;
        RECT 1130.070 13.470 1130.330 13.700 ;
        RECT 1130.390 13.470 1130.650 13.700 ;
        RECT 1130.710 13.470 1130.970 13.700 ;
        RECT 1131.030 13.470 1131.290 13.700 ;
        RECT 1131.350 13.470 1131.610 13.700 ;
        RECT 1131.670 13.470 1131.930 13.700 ;
        RECT 1219.110 13.470 1219.370 13.700 ;
        RECT 1219.430 13.470 1219.690 13.700 ;
        RECT 1219.750 13.470 1220.010 13.700 ;
        RECT 1220.070 13.470 1220.330 13.700 ;
        RECT 1220.390 13.470 1220.650 13.700 ;
        RECT 1220.710 13.470 1220.970 13.700 ;
        RECT 1221.030 13.470 1221.290 13.700 ;
        RECT 1221.350 13.470 1221.610 13.700 ;
        RECT 1221.670 13.470 1221.930 13.700 ;
        RECT 1309.110 13.470 1309.370 13.700 ;
        RECT 1309.430 13.470 1309.690 13.700 ;
        RECT 1309.750 13.470 1310.010 13.700 ;
        RECT 1310.070 13.470 1310.330 13.700 ;
        RECT 1310.390 13.470 1310.650 13.700 ;
        RECT 1310.710 13.470 1310.970 13.700 ;
        RECT 1311.030 13.470 1311.290 13.700 ;
        RECT 1311.350 13.470 1311.610 13.700 ;
        RECT 1311.670 13.470 1311.930 13.700 ;
        RECT 1399.110 13.470 1399.370 13.700 ;
        RECT 1399.430 13.470 1399.690 13.700 ;
        RECT 1399.750 13.470 1400.010 13.700 ;
        RECT 1400.070 13.470 1400.330 13.700 ;
        RECT 1400.390 13.470 1400.650 13.700 ;
        RECT 1400.710 13.470 1400.970 13.700 ;
        RECT 1401.030 13.470 1401.290 13.700 ;
        RECT 1401.350 13.470 1401.610 13.700 ;
        RECT 1401.670 13.470 1401.930 13.700 ;
        RECT 1489.110 13.470 1489.370 13.700 ;
        RECT 1489.430 13.470 1489.690 13.700 ;
        RECT 1489.750 13.470 1490.010 13.700 ;
        RECT 1490.070 13.470 1490.330 13.700 ;
        RECT 1490.390 13.470 1490.650 13.700 ;
        RECT 1490.710 13.470 1490.970 13.700 ;
        RECT 1491.030 13.470 1491.290 13.700 ;
        RECT 1491.350 13.470 1491.610 13.700 ;
        RECT 1491.670 13.470 1491.930 13.700 ;
        RECT 1579.110 13.470 1579.370 13.700 ;
        RECT 1579.430 13.470 1579.690 13.700 ;
        RECT 1579.750 13.470 1580.010 13.700 ;
        RECT 1580.070 13.470 1580.330 13.700 ;
        RECT 1580.390 13.470 1580.650 13.700 ;
        RECT 1580.710 13.470 1580.970 13.700 ;
        RECT 1581.030 13.470 1581.290 13.700 ;
        RECT 1581.350 13.470 1581.610 13.700 ;
        RECT 1581.670 13.470 1581.930 13.700 ;
        RECT 1669.110 13.470 1669.370 13.700 ;
        RECT 1669.430 13.470 1669.690 13.700 ;
        RECT 1669.750 13.470 1670.010 13.700 ;
        RECT 1670.070 13.470 1670.330 13.700 ;
        RECT 1670.390 13.470 1670.650 13.700 ;
        RECT 1670.710 13.470 1670.970 13.700 ;
        RECT 1671.030 13.470 1671.290 13.700 ;
        RECT 1671.350 13.470 1671.610 13.700 ;
        RECT 1671.670 13.470 1671.930 13.700 ;
        RECT 1759.110 13.470 1759.370 13.700 ;
        RECT 1759.430 13.470 1759.690 13.700 ;
        RECT 1759.750 13.470 1760.010 13.700 ;
        RECT 1760.070 13.470 1760.330 13.700 ;
        RECT 1760.390 13.470 1760.650 13.700 ;
        RECT 1760.710 13.470 1760.970 13.700 ;
        RECT 1761.030 13.470 1761.290 13.700 ;
        RECT 1761.350 13.470 1761.610 13.700 ;
        RECT 1761.670 13.470 1761.930 13.700 ;
        RECT 1849.110 13.470 1849.370 13.700 ;
        RECT 1849.430 13.470 1849.690 13.700 ;
        RECT 1849.750 13.470 1850.010 13.700 ;
        RECT 1850.070 13.470 1850.330 13.700 ;
        RECT 1850.390 13.470 1850.650 13.700 ;
        RECT 1850.710 13.470 1850.970 13.700 ;
        RECT 1851.030 13.470 1851.290 13.700 ;
        RECT 1851.350 13.470 1851.610 13.700 ;
        RECT 1851.670 13.470 1851.930 13.700 ;
        RECT 1939.110 13.470 1939.370 13.700 ;
        RECT 1939.430 13.470 1939.690 13.700 ;
        RECT 1939.750 13.470 1940.010 13.700 ;
        RECT 1940.070 13.470 1940.330 13.700 ;
        RECT 1940.390 13.470 1940.650 13.700 ;
        RECT 1940.710 13.470 1940.970 13.700 ;
        RECT 1941.030 13.470 1941.290 13.700 ;
        RECT 1941.350 13.470 1941.610 13.700 ;
        RECT 1941.670 13.470 1941.930 13.700 ;
        RECT 2029.110 13.470 2029.370 13.700 ;
        RECT 2029.430 13.470 2029.690 13.700 ;
        RECT 2029.750 13.470 2030.010 13.700 ;
        RECT 2030.070 13.470 2030.330 13.700 ;
        RECT 2030.390 13.470 2030.650 13.700 ;
        RECT 2030.710 13.470 2030.970 13.700 ;
        RECT 2031.030 13.470 2031.290 13.700 ;
        RECT 2031.350 13.470 2031.610 13.700 ;
        RECT 2031.670 13.470 2031.930 13.700 ;
        RECT 2119.110 13.470 2119.370 13.700 ;
        RECT 2119.430 13.470 2119.690 13.700 ;
        RECT 2119.750 13.470 2120.010 13.700 ;
        RECT 2120.070 13.470 2120.330 13.700 ;
        RECT 2120.390 13.470 2120.650 13.700 ;
        RECT 2120.710 13.470 2120.970 13.700 ;
        RECT 2121.030 13.470 2121.290 13.700 ;
        RECT 2121.350 13.470 2121.610 13.700 ;
        RECT 2121.670 13.470 2121.930 13.700 ;
        RECT 2209.110 13.470 2209.370 13.700 ;
        RECT 2209.430 13.470 2209.690 13.700 ;
        RECT 2209.750 13.470 2210.010 13.700 ;
        RECT 2210.070 13.470 2210.330 13.700 ;
        RECT 2210.390 13.470 2210.650 13.700 ;
        RECT 2210.710 13.470 2210.970 13.700 ;
        RECT 2211.030 13.470 2211.290 13.700 ;
        RECT 2211.350 13.470 2211.610 13.700 ;
        RECT 2211.670 13.470 2211.930 13.700 ;
        RECT 2299.110 13.470 2299.370 13.700 ;
        RECT 2299.430 13.470 2299.690 13.700 ;
        RECT 2299.750 13.470 2300.010 13.700 ;
        RECT 2300.070 13.470 2300.330 13.700 ;
        RECT 2300.390 13.470 2300.650 13.700 ;
        RECT 2300.710 13.470 2300.970 13.700 ;
        RECT 2301.030 13.470 2301.290 13.700 ;
        RECT 2301.350 13.470 2301.610 13.700 ;
        RECT 2301.670 13.470 2301.930 13.700 ;
        RECT 2389.110 13.470 2389.370 13.700 ;
        RECT 2389.430 13.470 2389.690 13.700 ;
        RECT 2389.750 13.470 2390.010 13.700 ;
        RECT 2390.070 13.470 2390.330 13.700 ;
        RECT 2390.390 13.470 2390.650 13.700 ;
        RECT 2390.710 13.470 2390.970 13.700 ;
        RECT 2391.030 13.470 2391.290 13.700 ;
        RECT 2391.350 13.470 2391.610 13.700 ;
        RECT 2391.670 13.470 2391.930 13.700 ;
        RECT 2479.110 13.470 2479.370 13.700 ;
        RECT 2479.430 13.470 2479.690 13.700 ;
        RECT 2479.750 13.470 2480.010 13.700 ;
        RECT 2480.070 13.470 2480.330 13.700 ;
        RECT 2480.390 13.470 2480.650 13.700 ;
        RECT 2480.710 13.470 2480.970 13.700 ;
        RECT 2481.030 13.470 2481.290 13.700 ;
        RECT 2481.350 13.470 2481.610 13.700 ;
        RECT 2481.670 13.470 2481.930 13.700 ;
        RECT 2569.110 13.470 2569.370 13.700 ;
        RECT 2569.430 13.470 2569.690 13.700 ;
        RECT 2569.750 13.470 2570.010 13.700 ;
        RECT 2570.070 13.470 2570.330 13.700 ;
        RECT 2570.390 13.470 2570.650 13.700 ;
        RECT 2570.710 13.470 2570.970 13.700 ;
        RECT 2571.030 13.470 2571.290 13.700 ;
        RECT 2571.350 13.470 2571.610 13.700 ;
        RECT 2571.670 13.470 2571.930 13.700 ;
        RECT 2659.110 13.470 2659.370 13.700 ;
        RECT 2659.430 13.470 2659.690 13.700 ;
        RECT 2659.750 13.470 2660.010 13.700 ;
        RECT 2660.070 13.470 2660.330 13.700 ;
        RECT 2660.390 13.470 2660.650 13.700 ;
        RECT 2660.710 13.470 2660.970 13.700 ;
        RECT 2661.030 13.470 2661.290 13.700 ;
        RECT 2661.350 13.470 2661.610 13.700 ;
        RECT 2661.670 13.470 2661.930 13.700 ;
        RECT 2749.110 13.470 2749.370 13.700 ;
        RECT 2749.430 13.470 2749.690 13.700 ;
        RECT 2749.750 13.470 2750.010 13.700 ;
        RECT 2750.070 13.470 2750.330 13.700 ;
        RECT 2750.390 13.470 2750.650 13.700 ;
        RECT 2750.710 13.470 2750.970 13.700 ;
        RECT 2751.030 13.470 2751.290 13.700 ;
        RECT 2751.350 13.470 2751.610 13.700 ;
        RECT 2751.670 13.470 2751.930 13.700 ;
        RECT 2839.110 13.470 2839.370 13.700 ;
        RECT 2839.430 13.470 2839.690 13.700 ;
        RECT 2839.750 13.470 2840.010 13.700 ;
        RECT 2840.070 13.470 2840.330 13.700 ;
        RECT 2840.390 13.470 2840.650 13.700 ;
        RECT 2840.710 13.470 2840.970 13.700 ;
        RECT 2841.030 13.470 2841.290 13.700 ;
        RECT 2841.350 13.470 2841.610 13.700 ;
        RECT 2841.670 13.470 2841.930 13.700 ;
      LAYER met2 ;
        RECT 49.110 3506.300 51.930 3506.320 ;
        RECT 139.110 3506.300 141.930 3506.320 ;
        RECT 229.110 3506.300 231.930 3506.320 ;
        RECT 319.110 3506.300 321.930 3506.320 ;
        RECT 409.110 3506.300 411.930 3506.320 ;
        RECT 499.110 3506.300 501.930 3506.320 ;
        RECT 589.110 3506.300 591.930 3506.320 ;
        RECT 679.110 3506.300 681.930 3506.320 ;
        RECT 769.110 3506.300 771.930 3506.320 ;
        RECT 859.110 3506.300 861.930 3506.320 ;
        RECT 949.110 3506.300 951.930 3506.320 ;
        RECT 1039.110 3506.300 1041.930 3506.320 ;
        RECT 1129.110 3506.300 1131.930 3506.320 ;
        RECT 1219.110 3506.300 1221.930 3506.320 ;
        RECT 1309.110 3506.300 1311.930 3506.320 ;
        RECT 1399.110 3506.300 1401.930 3506.320 ;
        RECT 1489.110 3506.300 1491.930 3506.320 ;
        RECT 1579.110 3506.300 1581.930 3506.320 ;
        RECT 1669.110 3506.300 1671.930 3506.320 ;
        RECT 1759.110 3506.300 1761.930 3506.320 ;
        RECT 1849.110 3506.300 1851.930 3506.320 ;
        RECT 1939.110 3506.300 1941.930 3506.320 ;
        RECT 2029.110 3506.300 2031.930 3506.320 ;
        RECT 2119.110 3506.300 2121.930 3506.320 ;
        RECT 2209.110 3506.300 2211.930 3506.320 ;
        RECT 2299.110 3506.300 2301.930 3506.320 ;
        RECT 2389.110 3506.300 2391.930 3506.320 ;
        RECT 2479.110 3506.300 2481.930 3506.320 ;
        RECT 2569.110 3506.300 2571.930 3506.320 ;
        RECT 2659.110 3506.300 2661.930 3506.320 ;
        RECT 2749.110 3506.300 2751.930 3506.320 ;
        RECT 2839.110 3506.300 2841.930 3506.320 ;
        RECT 49.110 13.360 51.930 13.700 ;
        RECT 139.110 13.360 141.930 13.700 ;
        RECT 229.110 13.360 231.930 13.700 ;
        RECT 319.110 13.360 321.930 13.700 ;
        RECT 409.110 13.360 411.930 13.700 ;
        RECT 499.110 13.360 501.930 13.700 ;
        RECT 589.110 13.360 591.930 13.700 ;
        RECT 679.110 13.360 681.930 13.700 ;
        RECT 769.110 13.360 771.930 13.700 ;
        RECT 859.110 13.360 861.930 13.700 ;
        RECT 949.110 13.360 951.930 13.700 ;
        RECT 1039.110 13.360 1041.930 13.700 ;
        RECT 1129.110 13.360 1131.930 13.700 ;
        RECT 1219.110 13.360 1221.930 13.700 ;
        RECT 1309.110 13.360 1311.930 13.700 ;
        RECT 1399.110 13.360 1401.930 13.700 ;
        RECT 1489.110 13.360 1491.930 13.700 ;
        RECT 1579.110 13.360 1581.930 13.700 ;
        RECT 1669.110 13.360 1671.930 13.700 ;
        RECT 1759.110 13.360 1761.930 13.700 ;
        RECT 1849.110 13.360 1851.930 13.700 ;
        RECT 1939.110 13.360 1941.930 13.700 ;
        RECT 2029.110 13.360 2031.930 13.700 ;
        RECT 2119.110 13.360 2121.930 13.700 ;
        RECT 2209.110 13.360 2211.930 13.700 ;
        RECT 2299.110 13.360 2301.930 13.700 ;
        RECT 2389.110 13.360 2391.930 13.700 ;
        RECT 2479.110 13.360 2481.930 13.700 ;
        RECT 2569.110 13.360 2571.930 13.700 ;
        RECT 2659.110 13.360 2661.930 13.700 ;
        RECT 2749.110 13.360 2751.930 13.700 ;
        RECT 2839.110 13.360 2841.930 13.700 ;
      LAYER via2 ;
        RECT 49.180 13.460 49.460 13.700 ;
        RECT 49.580 13.460 49.860 13.700 ;
        RECT 49.980 13.460 50.260 13.700 ;
        RECT 50.380 13.460 50.660 13.700 ;
        RECT 50.780 13.460 51.060 13.700 ;
        RECT 51.180 13.460 51.460 13.700 ;
        RECT 51.580 13.460 51.860 13.700 ;
        RECT 139.180 13.460 139.460 13.700 ;
        RECT 139.580 13.460 139.860 13.700 ;
        RECT 139.980 13.460 140.260 13.700 ;
        RECT 140.380 13.460 140.660 13.700 ;
        RECT 140.780 13.460 141.060 13.700 ;
        RECT 141.180 13.460 141.460 13.700 ;
        RECT 141.580 13.460 141.860 13.700 ;
        RECT 229.180 13.460 229.460 13.700 ;
        RECT 229.580 13.460 229.860 13.700 ;
        RECT 229.980 13.460 230.260 13.700 ;
        RECT 230.380 13.460 230.660 13.700 ;
        RECT 230.780 13.460 231.060 13.700 ;
        RECT 231.180 13.460 231.460 13.700 ;
        RECT 231.580 13.460 231.860 13.700 ;
        RECT 319.180 13.460 319.460 13.700 ;
        RECT 319.580 13.460 319.860 13.700 ;
        RECT 319.980 13.460 320.260 13.700 ;
        RECT 320.380 13.460 320.660 13.700 ;
        RECT 320.780 13.460 321.060 13.700 ;
        RECT 321.180 13.460 321.460 13.700 ;
        RECT 321.580 13.460 321.860 13.700 ;
        RECT 409.180 13.460 409.460 13.700 ;
        RECT 409.580 13.460 409.860 13.700 ;
        RECT 409.980 13.460 410.260 13.700 ;
        RECT 410.380 13.460 410.660 13.700 ;
        RECT 410.780 13.460 411.060 13.700 ;
        RECT 411.180 13.460 411.460 13.700 ;
        RECT 411.580 13.460 411.860 13.700 ;
        RECT 499.180 13.460 499.460 13.700 ;
        RECT 499.580 13.460 499.860 13.700 ;
        RECT 499.980 13.460 500.260 13.700 ;
        RECT 500.380 13.460 500.660 13.700 ;
        RECT 500.780 13.460 501.060 13.700 ;
        RECT 501.180 13.460 501.460 13.700 ;
        RECT 501.580 13.460 501.860 13.700 ;
        RECT 589.180 13.460 589.460 13.700 ;
        RECT 589.580 13.460 589.860 13.700 ;
        RECT 589.980 13.460 590.260 13.700 ;
        RECT 590.380 13.460 590.660 13.700 ;
        RECT 590.780 13.460 591.060 13.700 ;
        RECT 591.180 13.460 591.460 13.700 ;
        RECT 591.580 13.460 591.860 13.700 ;
        RECT 679.180 13.460 679.460 13.700 ;
        RECT 679.580 13.460 679.860 13.700 ;
        RECT 679.980 13.460 680.260 13.700 ;
        RECT 680.380 13.460 680.660 13.700 ;
        RECT 680.780 13.460 681.060 13.700 ;
        RECT 681.180 13.460 681.460 13.700 ;
        RECT 681.580 13.460 681.860 13.700 ;
        RECT 769.180 13.460 769.460 13.700 ;
        RECT 769.580 13.460 769.860 13.700 ;
        RECT 769.980 13.460 770.260 13.700 ;
        RECT 770.380 13.460 770.660 13.700 ;
        RECT 770.780 13.460 771.060 13.700 ;
        RECT 771.180 13.460 771.460 13.700 ;
        RECT 771.580 13.460 771.860 13.700 ;
        RECT 859.180 13.460 859.460 13.700 ;
        RECT 859.580 13.460 859.860 13.700 ;
        RECT 859.980 13.460 860.260 13.700 ;
        RECT 860.380 13.460 860.660 13.700 ;
        RECT 860.780 13.460 861.060 13.700 ;
        RECT 861.180 13.460 861.460 13.700 ;
        RECT 861.580 13.460 861.860 13.700 ;
        RECT 949.180 13.460 949.460 13.700 ;
        RECT 949.580 13.460 949.860 13.700 ;
        RECT 949.980 13.460 950.260 13.700 ;
        RECT 950.380 13.460 950.660 13.700 ;
        RECT 950.780 13.460 951.060 13.700 ;
        RECT 951.180 13.460 951.460 13.700 ;
        RECT 951.580 13.460 951.860 13.700 ;
        RECT 1039.180 13.460 1039.460 13.700 ;
        RECT 1039.580 13.460 1039.860 13.700 ;
        RECT 1039.980 13.460 1040.260 13.700 ;
        RECT 1040.380 13.460 1040.660 13.700 ;
        RECT 1040.780 13.460 1041.060 13.700 ;
        RECT 1041.180 13.460 1041.460 13.700 ;
        RECT 1041.580 13.460 1041.860 13.700 ;
        RECT 1129.180 13.460 1129.460 13.700 ;
        RECT 1129.580 13.460 1129.860 13.700 ;
        RECT 1129.980 13.460 1130.260 13.700 ;
        RECT 1130.380 13.460 1130.660 13.700 ;
        RECT 1130.780 13.460 1131.060 13.700 ;
        RECT 1131.180 13.460 1131.460 13.700 ;
        RECT 1131.580 13.460 1131.860 13.700 ;
        RECT 1219.180 13.460 1219.460 13.700 ;
        RECT 1219.580 13.460 1219.860 13.700 ;
        RECT 1219.980 13.460 1220.260 13.700 ;
        RECT 1220.380 13.460 1220.660 13.700 ;
        RECT 1220.780 13.460 1221.060 13.700 ;
        RECT 1221.180 13.460 1221.460 13.700 ;
        RECT 1221.580 13.460 1221.860 13.700 ;
        RECT 1309.180 13.460 1309.460 13.700 ;
        RECT 1309.580 13.460 1309.860 13.700 ;
        RECT 1309.980 13.460 1310.260 13.700 ;
        RECT 1310.380 13.460 1310.660 13.700 ;
        RECT 1310.780 13.460 1311.060 13.700 ;
        RECT 1311.180 13.460 1311.460 13.700 ;
        RECT 1311.580 13.460 1311.860 13.700 ;
        RECT 1399.180 13.460 1399.460 13.700 ;
        RECT 1399.580 13.460 1399.860 13.700 ;
        RECT 1399.980 13.460 1400.260 13.700 ;
        RECT 1400.380 13.460 1400.660 13.700 ;
        RECT 1400.780 13.460 1401.060 13.700 ;
        RECT 1401.180 13.460 1401.460 13.700 ;
        RECT 1401.580 13.460 1401.860 13.700 ;
        RECT 1489.180 13.460 1489.460 13.700 ;
        RECT 1489.580 13.460 1489.860 13.700 ;
        RECT 1489.980 13.460 1490.260 13.700 ;
        RECT 1490.380 13.460 1490.660 13.700 ;
        RECT 1490.780 13.460 1491.060 13.700 ;
        RECT 1491.180 13.460 1491.460 13.700 ;
        RECT 1491.580 13.460 1491.860 13.700 ;
        RECT 1579.180 13.460 1579.460 13.700 ;
        RECT 1579.580 13.460 1579.860 13.700 ;
        RECT 1579.980 13.460 1580.260 13.700 ;
        RECT 1580.380 13.460 1580.660 13.700 ;
        RECT 1580.780 13.460 1581.060 13.700 ;
        RECT 1581.180 13.460 1581.460 13.700 ;
        RECT 1581.580 13.460 1581.860 13.700 ;
        RECT 1669.180 13.460 1669.460 13.700 ;
        RECT 1669.580 13.460 1669.860 13.700 ;
        RECT 1669.980 13.460 1670.260 13.700 ;
        RECT 1670.380 13.460 1670.660 13.700 ;
        RECT 1670.780 13.460 1671.060 13.700 ;
        RECT 1671.180 13.460 1671.460 13.700 ;
        RECT 1671.580 13.460 1671.860 13.700 ;
        RECT 1759.180 13.460 1759.460 13.700 ;
        RECT 1759.580 13.460 1759.860 13.700 ;
        RECT 1759.980 13.460 1760.260 13.700 ;
        RECT 1760.380 13.460 1760.660 13.700 ;
        RECT 1760.780 13.460 1761.060 13.700 ;
        RECT 1761.180 13.460 1761.460 13.700 ;
        RECT 1761.580 13.460 1761.860 13.700 ;
        RECT 1849.180 13.460 1849.460 13.700 ;
        RECT 1849.580 13.460 1849.860 13.700 ;
        RECT 1849.980 13.460 1850.260 13.700 ;
        RECT 1850.380 13.460 1850.660 13.700 ;
        RECT 1850.780 13.460 1851.060 13.700 ;
        RECT 1851.180 13.460 1851.460 13.700 ;
        RECT 1851.580 13.460 1851.860 13.700 ;
        RECT 1939.180 13.460 1939.460 13.700 ;
        RECT 1939.580 13.460 1939.860 13.700 ;
        RECT 1939.980 13.460 1940.260 13.700 ;
        RECT 1940.380 13.460 1940.660 13.700 ;
        RECT 1940.780 13.460 1941.060 13.700 ;
        RECT 1941.180 13.460 1941.460 13.700 ;
        RECT 1941.580 13.460 1941.860 13.700 ;
        RECT 2029.180 13.460 2029.460 13.700 ;
        RECT 2029.580 13.460 2029.860 13.700 ;
        RECT 2029.980 13.460 2030.260 13.700 ;
        RECT 2030.380 13.460 2030.660 13.700 ;
        RECT 2030.780 13.460 2031.060 13.700 ;
        RECT 2031.180 13.460 2031.460 13.700 ;
        RECT 2031.580 13.460 2031.860 13.700 ;
        RECT 2119.180 13.460 2119.460 13.700 ;
        RECT 2119.580 13.460 2119.860 13.700 ;
        RECT 2119.980 13.460 2120.260 13.700 ;
        RECT 2120.380 13.460 2120.660 13.700 ;
        RECT 2120.780 13.460 2121.060 13.700 ;
        RECT 2121.180 13.460 2121.460 13.700 ;
        RECT 2121.580 13.460 2121.860 13.700 ;
        RECT 2209.180 13.460 2209.460 13.700 ;
        RECT 2209.580 13.460 2209.860 13.700 ;
        RECT 2209.980 13.460 2210.260 13.700 ;
        RECT 2210.380 13.460 2210.660 13.700 ;
        RECT 2210.780 13.460 2211.060 13.700 ;
        RECT 2211.180 13.460 2211.460 13.700 ;
        RECT 2211.580 13.460 2211.860 13.700 ;
        RECT 2299.180 13.460 2299.460 13.700 ;
        RECT 2299.580 13.460 2299.860 13.700 ;
        RECT 2299.980 13.460 2300.260 13.700 ;
        RECT 2300.380 13.460 2300.660 13.700 ;
        RECT 2300.780 13.460 2301.060 13.700 ;
        RECT 2301.180 13.460 2301.460 13.700 ;
        RECT 2301.580 13.460 2301.860 13.700 ;
        RECT 2389.180 13.460 2389.460 13.700 ;
        RECT 2389.580 13.460 2389.860 13.700 ;
        RECT 2389.980 13.460 2390.260 13.700 ;
        RECT 2390.380 13.460 2390.660 13.700 ;
        RECT 2390.780 13.460 2391.060 13.700 ;
        RECT 2391.180 13.460 2391.460 13.700 ;
        RECT 2391.580 13.460 2391.860 13.700 ;
        RECT 2479.180 13.460 2479.460 13.700 ;
        RECT 2479.580 13.460 2479.860 13.700 ;
        RECT 2479.980 13.460 2480.260 13.700 ;
        RECT 2480.380 13.460 2480.660 13.700 ;
        RECT 2480.780 13.460 2481.060 13.700 ;
        RECT 2481.180 13.460 2481.460 13.700 ;
        RECT 2481.580 13.460 2481.860 13.700 ;
        RECT 2569.180 13.460 2569.460 13.700 ;
        RECT 2569.580 13.460 2569.860 13.700 ;
        RECT 2569.980 13.460 2570.260 13.700 ;
        RECT 2570.380 13.460 2570.660 13.700 ;
        RECT 2570.780 13.460 2571.060 13.700 ;
        RECT 2571.180 13.460 2571.460 13.700 ;
        RECT 2571.580 13.460 2571.860 13.700 ;
        RECT 2659.180 13.460 2659.460 13.700 ;
        RECT 2659.580 13.460 2659.860 13.700 ;
        RECT 2659.980 13.460 2660.260 13.700 ;
        RECT 2660.380 13.460 2660.660 13.700 ;
        RECT 2660.780 13.460 2661.060 13.700 ;
        RECT 2661.180 13.460 2661.460 13.700 ;
        RECT 2661.580 13.460 2661.860 13.700 ;
        RECT 2749.180 13.460 2749.460 13.700 ;
        RECT 2749.580 13.460 2749.860 13.700 ;
        RECT 2749.980 13.460 2750.260 13.700 ;
        RECT 2750.380 13.460 2750.660 13.700 ;
        RECT 2750.780 13.460 2751.060 13.700 ;
        RECT 2751.180 13.460 2751.460 13.700 ;
        RECT 2751.580 13.460 2751.860 13.700 ;
        RECT 2839.180 13.460 2839.460 13.700 ;
        RECT 2839.580 13.460 2839.860 13.700 ;
        RECT 2839.980 13.460 2840.260 13.700 ;
        RECT 2840.380 13.460 2840.660 13.700 ;
        RECT 2840.780 13.460 2841.060 13.700 ;
        RECT 2841.180 13.460 2841.460 13.700 ;
        RECT 2841.580 13.460 2841.860 13.700 ;
      LAYER met3 ;
        RECT 49.020 13.435 52.020 13.700 ;
        RECT 139.020 13.435 142.020 13.700 ;
        RECT 229.020 13.435 232.020 13.700 ;
        RECT 319.020 13.435 322.020 13.700 ;
        RECT 409.020 13.435 412.020 13.700 ;
        RECT 499.020 13.435 502.020 13.700 ;
        RECT 589.020 13.435 592.020 13.700 ;
        RECT 679.020 13.435 682.020 13.700 ;
        RECT 769.020 13.435 772.020 13.700 ;
        RECT 859.020 13.435 862.020 13.700 ;
        RECT 949.020 13.435 952.020 13.700 ;
        RECT 1039.020 13.435 1042.020 13.700 ;
        RECT 1129.020 13.435 1132.020 13.700 ;
        RECT 1219.020 13.435 1222.020 13.700 ;
        RECT 1309.020 13.435 1312.020 13.700 ;
        RECT 1399.020 13.435 1402.020 13.700 ;
        RECT 1489.020 13.435 1492.020 13.700 ;
        RECT 1579.020 13.435 1582.020 13.700 ;
        RECT 1669.020 13.435 1672.020 13.700 ;
        RECT 1759.020 13.435 1762.020 13.700 ;
        RECT 1849.020 13.435 1852.020 13.700 ;
        RECT 1939.020 13.435 1942.020 13.700 ;
        RECT 2029.020 13.435 2032.020 13.700 ;
        RECT 2119.020 13.435 2122.020 13.700 ;
        RECT 2209.020 13.435 2212.020 13.700 ;
        RECT 2299.020 13.435 2302.020 13.700 ;
        RECT 2389.020 13.435 2392.020 13.700 ;
        RECT 2479.020 13.435 2482.020 13.700 ;
        RECT 2569.020 13.435 2572.020 13.700 ;
        RECT 2659.020 13.435 2662.020 13.700 ;
        RECT 2749.020 13.435 2752.020 13.700 ;
        RECT 2839.020 13.435 2842.020 13.700 ;
      LAYER via3 ;
        RECT 49.160 13.440 49.480 13.700 ;
        RECT 49.560 13.440 49.880 13.700 ;
        RECT 49.960 13.440 50.280 13.700 ;
        RECT 50.360 13.440 50.680 13.700 ;
        RECT 50.760 13.440 51.080 13.700 ;
        RECT 51.160 13.440 51.480 13.700 ;
        RECT 51.560 13.440 51.880 13.700 ;
        RECT 139.160 13.440 139.480 13.700 ;
        RECT 139.560 13.440 139.880 13.700 ;
        RECT 139.960 13.440 140.280 13.700 ;
        RECT 140.360 13.440 140.680 13.700 ;
        RECT 140.760 13.440 141.080 13.700 ;
        RECT 141.160 13.440 141.480 13.700 ;
        RECT 141.560 13.440 141.880 13.700 ;
        RECT 229.160 13.440 229.480 13.700 ;
        RECT 229.560 13.440 229.880 13.700 ;
        RECT 229.960 13.440 230.280 13.700 ;
        RECT 230.360 13.440 230.680 13.700 ;
        RECT 230.760 13.440 231.080 13.700 ;
        RECT 231.160 13.440 231.480 13.700 ;
        RECT 231.560 13.440 231.880 13.700 ;
        RECT 319.160 13.440 319.480 13.700 ;
        RECT 319.560 13.440 319.880 13.700 ;
        RECT 319.960 13.440 320.280 13.700 ;
        RECT 320.360 13.440 320.680 13.700 ;
        RECT 320.760 13.440 321.080 13.700 ;
        RECT 321.160 13.440 321.480 13.700 ;
        RECT 321.560 13.440 321.880 13.700 ;
        RECT 409.160 13.440 409.480 13.700 ;
        RECT 409.560 13.440 409.880 13.700 ;
        RECT 409.960 13.440 410.280 13.700 ;
        RECT 410.360 13.440 410.680 13.700 ;
        RECT 410.760 13.440 411.080 13.700 ;
        RECT 411.160 13.440 411.480 13.700 ;
        RECT 411.560 13.440 411.880 13.700 ;
        RECT 499.160 13.440 499.480 13.700 ;
        RECT 499.560 13.440 499.880 13.700 ;
        RECT 499.960 13.440 500.280 13.700 ;
        RECT 500.360 13.440 500.680 13.700 ;
        RECT 500.760 13.440 501.080 13.700 ;
        RECT 501.160 13.440 501.480 13.700 ;
        RECT 501.560 13.440 501.880 13.700 ;
        RECT 589.160 13.440 589.480 13.700 ;
        RECT 589.560 13.440 589.880 13.700 ;
        RECT 589.960 13.440 590.280 13.700 ;
        RECT 590.360 13.440 590.680 13.700 ;
        RECT 590.760 13.440 591.080 13.700 ;
        RECT 591.160 13.440 591.480 13.700 ;
        RECT 591.560 13.440 591.880 13.700 ;
        RECT 679.160 13.440 679.480 13.700 ;
        RECT 679.560 13.440 679.880 13.700 ;
        RECT 679.960 13.440 680.280 13.700 ;
        RECT 680.360 13.440 680.680 13.700 ;
        RECT 680.760 13.440 681.080 13.700 ;
        RECT 681.160 13.440 681.480 13.700 ;
        RECT 681.560 13.440 681.880 13.700 ;
        RECT 769.160 13.440 769.480 13.700 ;
        RECT 769.560 13.440 769.880 13.700 ;
        RECT 769.960 13.440 770.280 13.700 ;
        RECT 770.360 13.440 770.680 13.700 ;
        RECT 770.760 13.440 771.080 13.700 ;
        RECT 771.160 13.440 771.480 13.700 ;
        RECT 771.560 13.440 771.880 13.700 ;
        RECT 859.160 13.440 859.480 13.700 ;
        RECT 859.560 13.440 859.880 13.700 ;
        RECT 859.960 13.440 860.280 13.700 ;
        RECT 860.360 13.440 860.680 13.700 ;
        RECT 860.760 13.440 861.080 13.700 ;
        RECT 861.160 13.440 861.480 13.700 ;
        RECT 861.560 13.440 861.880 13.700 ;
        RECT 949.160 13.440 949.480 13.700 ;
        RECT 949.560 13.440 949.880 13.700 ;
        RECT 949.960 13.440 950.280 13.700 ;
        RECT 950.360 13.440 950.680 13.700 ;
        RECT 950.760 13.440 951.080 13.700 ;
        RECT 951.160 13.440 951.480 13.700 ;
        RECT 951.560 13.440 951.880 13.700 ;
        RECT 1039.160 13.440 1039.480 13.700 ;
        RECT 1039.560 13.440 1039.880 13.700 ;
        RECT 1039.960 13.440 1040.280 13.700 ;
        RECT 1040.360 13.440 1040.680 13.700 ;
        RECT 1040.760 13.440 1041.080 13.700 ;
        RECT 1041.160 13.440 1041.480 13.700 ;
        RECT 1041.560 13.440 1041.880 13.700 ;
        RECT 1129.160 13.440 1129.480 13.700 ;
        RECT 1129.560 13.440 1129.880 13.700 ;
        RECT 1129.960 13.440 1130.280 13.700 ;
        RECT 1130.360 13.440 1130.680 13.700 ;
        RECT 1130.760 13.440 1131.080 13.700 ;
        RECT 1131.160 13.440 1131.480 13.700 ;
        RECT 1131.560 13.440 1131.880 13.700 ;
        RECT 1219.160 13.440 1219.480 13.700 ;
        RECT 1219.560 13.440 1219.880 13.700 ;
        RECT 1219.960 13.440 1220.280 13.700 ;
        RECT 1220.360 13.440 1220.680 13.700 ;
        RECT 1220.760 13.440 1221.080 13.700 ;
        RECT 1221.160 13.440 1221.480 13.700 ;
        RECT 1221.560 13.440 1221.880 13.700 ;
        RECT 1309.160 13.440 1309.480 13.700 ;
        RECT 1309.560 13.440 1309.880 13.700 ;
        RECT 1309.960 13.440 1310.280 13.700 ;
        RECT 1310.360 13.440 1310.680 13.700 ;
        RECT 1310.760 13.440 1311.080 13.700 ;
        RECT 1311.160 13.440 1311.480 13.700 ;
        RECT 1311.560 13.440 1311.880 13.700 ;
        RECT 1399.160 13.440 1399.480 13.700 ;
        RECT 1399.560 13.440 1399.880 13.700 ;
        RECT 1399.960 13.440 1400.280 13.700 ;
        RECT 1400.360 13.440 1400.680 13.700 ;
        RECT 1400.760 13.440 1401.080 13.700 ;
        RECT 1401.160 13.440 1401.480 13.700 ;
        RECT 1401.560 13.440 1401.880 13.700 ;
        RECT 1489.160 13.440 1489.480 13.700 ;
        RECT 1489.560 13.440 1489.880 13.700 ;
        RECT 1489.960 13.440 1490.280 13.700 ;
        RECT 1490.360 13.440 1490.680 13.700 ;
        RECT 1490.760 13.440 1491.080 13.700 ;
        RECT 1491.160 13.440 1491.480 13.700 ;
        RECT 1491.560 13.440 1491.880 13.700 ;
        RECT 1579.160 13.440 1579.480 13.700 ;
        RECT 1579.560 13.440 1579.880 13.700 ;
        RECT 1579.960 13.440 1580.280 13.700 ;
        RECT 1580.360 13.440 1580.680 13.700 ;
        RECT 1580.760 13.440 1581.080 13.700 ;
        RECT 1581.160 13.440 1581.480 13.700 ;
        RECT 1581.560 13.440 1581.880 13.700 ;
        RECT 1669.160 13.440 1669.480 13.700 ;
        RECT 1669.560 13.440 1669.880 13.700 ;
        RECT 1669.960 13.440 1670.280 13.700 ;
        RECT 1670.360 13.440 1670.680 13.700 ;
        RECT 1670.760 13.440 1671.080 13.700 ;
        RECT 1671.160 13.440 1671.480 13.700 ;
        RECT 1671.560 13.440 1671.880 13.700 ;
        RECT 1759.160 13.440 1759.480 13.700 ;
        RECT 1759.560 13.440 1759.880 13.700 ;
        RECT 1759.960 13.440 1760.280 13.700 ;
        RECT 1760.360 13.440 1760.680 13.700 ;
        RECT 1760.760 13.440 1761.080 13.700 ;
        RECT 1761.160 13.440 1761.480 13.700 ;
        RECT 1761.560 13.440 1761.880 13.700 ;
        RECT 1849.160 13.440 1849.480 13.700 ;
        RECT 1849.560 13.440 1849.880 13.700 ;
        RECT 1849.960 13.440 1850.280 13.700 ;
        RECT 1850.360 13.440 1850.680 13.700 ;
        RECT 1850.760 13.440 1851.080 13.700 ;
        RECT 1851.160 13.440 1851.480 13.700 ;
        RECT 1851.560 13.440 1851.880 13.700 ;
        RECT 1939.160 13.440 1939.480 13.700 ;
        RECT 1939.560 13.440 1939.880 13.700 ;
        RECT 1939.960 13.440 1940.280 13.700 ;
        RECT 1940.360 13.440 1940.680 13.700 ;
        RECT 1940.760 13.440 1941.080 13.700 ;
        RECT 1941.160 13.440 1941.480 13.700 ;
        RECT 1941.560 13.440 1941.880 13.700 ;
        RECT 2029.160 13.440 2029.480 13.700 ;
        RECT 2029.560 13.440 2029.880 13.700 ;
        RECT 2029.960 13.440 2030.280 13.700 ;
        RECT 2030.360 13.440 2030.680 13.700 ;
        RECT 2030.760 13.440 2031.080 13.700 ;
        RECT 2031.160 13.440 2031.480 13.700 ;
        RECT 2031.560 13.440 2031.880 13.700 ;
        RECT 2119.160 13.440 2119.480 13.700 ;
        RECT 2119.560 13.440 2119.880 13.700 ;
        RECT 2119.960 13.440 2120.280 13.700 ;
        RECT 2120.360 13.440 2120.680 13.700 ;
        RECT 2120.760 13.440 2121.080 13.700 ;
        RECT 2121.160 13.440 2121.480 13.700 ;
        RECT 2121.560 13.440 2121.880 13.700 ;
        RECT 2209.160 13.440 2209.480 13.700 ;
        RECT 2209.560 13.440 2209.880 13.700 ;
        RECT 2209.960 13.440 2210.280 13.700 ;
        RECT 2210.360 13.440 2210.680 13.700 ;
        RECT 2210.760 13.440 2211.080 13.700 ;
        RECT 2211.160 13.440 2211.480 13.700 ;
        RECT 2211.560 13.440 2211.880 13.700 ;
        RECT 2299.160 13.440 2299.480 13.700 ;
        RECT 2299.560 13.440 2299.880 13.700 ;
        RECT 2299.960 13.440 2300.280 13.700 ;
        RECT 2300.360 13.440 2300.680 13.700 ;
        RECT 2300.760 13.440 2301.080 13.700 ;
        RECT 2301.160 13.440 2301.480 13.700 ;
        RECT 2301.560 13.440 2301.880 13.700 ;
        RECT 2389.160 13.440 2389.480 13.700 ;
        RECT 2389.560 13.440 2389.880 13.700 ;
        RECT 2389.960 13.440 2390.280 13.700 ;
        RECT 2390.360 13.440 2390.680 13.700 ;
        RECT 2390.760 13.440 2391.080 13.700 ;
        RECT 2391.160 13.440 2391.480 13.700 ;
        RECT 2391.560 13.440 2391.880 13.700 ;
        RECT 2479.160 13.440 2479.480 13.700 ;
        RECT 2479.560 13.440 2479.880 13.700 ;
        RECT 2479.960 13.440 2480.280 13.700 ;
        RECT 2480.360 13.440 2480.680 13.700 ;
        RECT 2480.760 13.440 2481.080 13.700 ;
        RECT 2481.160 13.440 2481.480 13.700 ;
        RECT 2481.560 13.440 2481.880 13.700 ;
        RECT 2569.160 13.440 2569.480 13.700 ;
        RECT 2569.560 13.440 2569.880 13.700 ;
        RECT 2569.960 13.440 2570.280 13.700 ;
        RECT 2570.360 13.440 2570.680 13.700 ;
        RECT 2570.760 13.440 2571.080 13.700 ;
        RECT 2571.160 13.440 2571.480 13.700 ;
        RECT 2571.560 13.440 2571.880 13.700 ;
        RECT 2659.160 13.440 2659.480 13.700 ;
        RECT 2659.560 13.440 2659.880 13.700 ;
        RECT 2659.960 13.440 2660.280 13.700 ;
        RECT 2660.360 13.440 2660.680 13.700 ;
        RECT 2660.760 13.440 2661.080 13.700 ;
        RECT 2661.160 13.440 2661.480 13.700 ;
        RECT 2661.560 13.440 2661.880 13.700 ;
        RECT 2749.160 13.440 2749.480 13.700 ;
        RECT 2749.560 13.440 2749.880 13.700 ;
        RECT 2749.960 13.440 2750.280 13.700 ;
        RECT 2750.360 13.440 2750.680 13.700 ;
        RECT 2750.760 13.440 2751.080 13.700 ;
        RECT 2751.160 13.440 2751.480 13.700 ;
        RECT 2751.560 13.440 2751.880 13.700 ;
        RECT 2839.160 13.440 2839.480 13.700 ;
        RECT 2839.560 13.440 2839.880 13.700 ;
        RECT 2839.960 13.440 2840.280 13.700 ;
        RECT 2840.360 13.440 2840.680 13.700 ;
        RECT 2840.760 13.440 2841.080 13.700 ;
        RECT 2841.160 13.440 2841.480 13.700 ;
        RECT 2841.560 13.440 2841.880 13.700 ;
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 49.020 3506.300 52.020 3529.000 ;
        RECT 139.020 3506.300 142.020 3529.000 ;
        RECT 229.020 3506.300 232.020 3529.000 ;
        RECT 319.020 3506.300 322.020 3529.000 ;
        RECT 409.020 3506.300 412.020 3529.000 ;
        RECT 499.020 3506.300 502.020 3529.000 ;
        RECT 589.020 3506.300 592.020 3529.000 ;
        RECT 679.020 3506.300 682.020 3529.000 ;
        RECT 769.020 3506.300 772.020 3529.000 ;
        RECT 859.020 3506.300 862.020 3529.000 ;
        RECT 949.020 3506.300 952.020 3529.000 ;
        RECT 1039.020 3506.300 1042.020 3529.000 ;
        RECT 1129.020 3506.300 1132.020 3529.000 ;
        RECT 1219.020 3506.300 1222.020 3529.000 ;
        RECT 1309.020 3506.300 1312.020 3529.000 ;
        RECT 1399.020 3506.300 1402.020 3529.000 ;
        RECT 1489.020 3506.300 1492.020 3529.000 ;
        RECT 1579.020 3506.300 1582.020 3529.000 ;
        RECT 1669.020 3506.300 1672.020 3529.000 ;
        RECT 1759.020 3506.300 1762.020 3529.000 ;
        RECT 1849.020 3506.300 1852.020 3529.000 ;
        RECT 1939.020 3506.300 1942.020 3529.000 ;
        RECT 2029.020 3506.300 2032.020 3529.000 ;
        RECT 2119.020 3506.300 2122.020 3529.000 ;
        RECT 2209.020 3506.300 2212.020 3529.000 ;
        RECT 2299.020 3506.300 2302.020 3529.000 ;
        RECT 2389.020 3506.300 2392.020 3529.000 ;
        RECT 2479.020 3506.300 2482.020 3529.000 ;
        RECT 2569.020 3506.300 2572.020 3529.000 ;
        RECT 2659.020 3506.300 2662.020 3529.000 ;
        RECT 2749.020 3506.300 2752.020 3529.000 ;
        RECT 2839.020 3506.300 2842.020 3529.000 ;
        RECT 49.020 -9.320 52.020 13.700 ;
        RECT 139.020 -9.320 142.020 13.700 ;
        RECT 229.020 -9.320 232.020 13.700 ;
        RECT 319.020 -9.320 322.020 13.700 ;
        RECT 409.020 -9.320 412.020 13.700 ;
        RECT 499.020 -9.320 502.020 13.700 ;
        RECT 589.020 -9.320 592.020 13.700 ;
        RECT 679.020 -9.320 682.020 13.700 ;
        RECT 769.020 -9.320 772.020 13.700 ;
        RECT 859.020 -9.320 862.020 13.700 ;
        RECT 949.020 -9.320 952.020 13.700 ;
        RECT 1039.020 -9.320 1042.020 13.700 ;
        RECT 1129.020 -9.320 1132.020 13.700 ;
        RECT 1219.020 -9.320 1222.020 13.700 ;
        RECT 1309.020 -9.320 1312.020 13.700 ;
        RECT 1399.020 -9.320 1402.020 13.700 ;
        RECT 1489.020 -9.320 1492.020 13.700 ;
        RECT 1579.020 -9.320 1582.020 13.700 ;
        RECT 1669.020 -9.320 1672.020 13.700 ;
        RECT 1759.020 -9.320 1762.020 13.700 ;
        RECT 1849.020 -9.320 1852.020 13.700 ;
        RECT 1939.020 -9.320 1942.020 13.700 ;
        RECT 2029.020 -9.320 2032.020 13.700 ;
        RECT 2119.020 -9.320 2122.020 13.700 ;
        RECT 2209.020 -9.320 2212.020 13.700 ;
        RECT 2299.020 -9.320 2302.020 13.700 ;
        RECT 2389.020 -9.320 2392.020 13.700 ;
        RECT 2479.020 -9.320 2482.020 13.700 ;
        RECT 2569.020 -9.320 2572.020 13.700 ;
        RECT 2659.020 -9.320 2662.020 13.700 ;
        RECT 2749.020 -9.320 2752.020 13.700 ;
        RECT 2839.020 -9.320 2842.020 13.700 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 49.930 3527.710 51.110 3528.890 ;
        RECT 49.930 3526.110 51.110 3527.290 ;
        RECT 139.930 3527.710 141.110 3528.890 ;
        RECT 139.930 3526.110 141.110 3527.290 ;
        RECT 229.930 3527.710 231.110 3528.890 ;
        RECT 229.930 3526.110 231.110 3527.290 ;
        RECT 319.930 3527.710 321.110 3528.890 ;
        RECT 319.930 3526.110 321.110 3527.290 ;
        RECT 409.930 3527.710 411.110 3528.890 ;
        RECT 409.930 3526.110 411.110 3527.290 ;
        RECT 499.930 3527.710 501.110 3528.890 ;
        RECT 499.930 3526.110 501.110 3527.290 ;
        RECT 589.930 3527.710 591.110 3528.890 ;
        RECT 589.930 3526.110 591.110 3527.290 ;
        RECT 679.930 3527.710 681.110 3528.890 ;
        RECT 679.930 3526.110 681.110 3527.290 ;
        RECT 769.930 3527.710 771.110 3528.890 ;
        RECT 769.930 3526.110 771.110 3527.290 ;
        RECT 859.930 3527.710 861.110 3528.890 ;
        RECT 859.930 3526.110 861.110 3527.290 ;
        RECT 949.930 3527.710 951.110 3528.890 ;
        RECT 949.930 3526.110 951.110 3527.290 ;
        RECT 1039.930 3527.710 1041.110 3528.890 ;
        RECT 1039.930 3526.110 1041.110 3527.290 ;
        RECT 1129.930 3527.710 1131.110 3528.890 ;
        RECT 1129.930 3526.110 1131.110 3527.290 ;
        RECT 1219.930 3527.710 1221.110 3528.890 ;
        RECT 1219.930 3526.110 1221.110 3527.290 ;
        RECT 1309.930 3527.710 1311.110 3528.890 ;
        RECT 1309.930 3526.110 1311.110 3527.290 ;
        RECT 1399.930 3527.710 1401.110 3528.890 ;
        RECT 1399.930 3526.110 1401.110 3527.290 ;
        RECT 1489.930 3527.710 1491.110 3528.890 ;
        RECT 1489.930 3526.110 1491.110 3527.290 ;
        RECT 1579.930 3527.710 1581.110 3528.890 ;
        RECT 1579.930 3526.110 1581.110 3527.290 ;
        RECT 1669.930 3527.710 1671.110 3528.890 ;
        RECT 1669.930 3526.110 1671.110 3527.290 ;
        RECT 1759.930 3527.710 1761.110 3528.890 ;
        RECT 1759.930 3526.110 1761.110 3527.290 ;
        RECT 1849.930 3527.710 1851.110 3528.890 ;
        RECT 1849.930 3526.110 1851.110 3527.290 ;
        RECT 1939.930 3527.710 1941.110 3528.890 ;
        RECT 1939.930 3526.110 1941.110 3527.290 ;
        RECT 2029.930 3527.710 2031.110 3528.890 ;
        RECT 2029.930 3526.110 2031.110 3527.290 ;
        RECT 2119.930 3527.710 2121.110 3528.890 ;
        RECT 2119.930 3526.110 2121.110 3527.290 ;
        RECT 2209.930 3527.710 2211.110 3528.890 ;
        RECT 2209.930 3526.110 2211.110 3527.290 ;
        RECT 2299.930 3527.710 2301.110 3528.890 ;
        RECT 2299.930 3526.110 2301.110 3527.290 ;
        RECT 2389.930 3527.710 2391.110 3528.890 ;
        RECT 2389.930 3526.110 2391.110 3527.290 ;
        RECT 2479.930 3527.710 2481.110 3528.890 ;
        RECT 2479.930 3526.110 2481.110 3527.290 ;
        RECT 2569.930 3527.710 2571.110 3528.890 ;
        RECT 2569.930 3526.110 2571.110 3527.290 ;
        RECT 2659.930 3527.710 2661.110 3528.890 ;
        RECT 2659.930 3526.110 2661.110 3527.290 ;
        RECT 2749.930 3527.710 2751.110 3528.890 ;
        RECT 2749.930 3526.110 2751.110 3527.290 ;
        RECT 2839.930 3527.710 2841.110 3528.890 ;
        RECT 2839.930 3526.110 2841.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3475.850 -12.590 3477.030 ;
        RECT -13.770 3474.250 -12.590 3475.430 ;
        RECT -13.770 3385.850 -12.590 3387.030 ;
        RECT -13.770 3384.250 -12.590 3385.430 ;
        RECT -13.770 3295.850 -12.590 3297.030 ;
        RECT -13.770 3294.250 -12.590 3295.430 ;
        RECT -13.770 3205.850 -12.590 3207.030 ;
        RECT -13.770 3204.250 -12.590 3205.430 ;
        RECT -13.770 3115.850 -12.590 3117.030 ;
        RECT -13.770 3114.250 -12.590 3115.430 ;
        RECT -13.770 3025.850 -12.590 3027.030 ;
        RECT -13.770 3024.250 -12.590 3025.430 ;
        RECT -13.770 2935.850 -12.590 2937.030 ;
        RECT -13.770 2934.250 -12.590 2935.430 ;
        RECT -13.770 2845.850 -12.590 2847.030 ;
        RECT -13.770 2844.250 -12.590 2845.430 ;
        RECT -13.770 2755.850 -12.590 2757.030 ;
        RECT -13.770 2754.250 -12.590 2755.430 ;
        RECT -13.770 2665.850 -12.590 2667.030 ;
        RECT -13.770 2664.250 -12.590 2665.430 ;
        RECT -13.770 2575.850 -12.590 2577.030 ;
        RECT -13.770 2574.250 -12.590 2575.430 ;
        RECT -13.770 2485.850 -12.590 2487.030 ;
        RECT -13.770 2484.250 -12.590 2485.430 ;
        RECT -13.770 2395.850 -12.590 2397.030 ;
        RECT -13.770 2394.250 -12.590 2395.430 ;
        RECT -13.770 2305.850 -12.590 2307.030 ;
        RECT -13.770 2304.250 -12.590 2305.430 ;
        RECT -13.770 2215.850 -12.590 2217.030 ;
        RECT -13.770 2214.250 -12.590 2215.430 ;
        RECT -13.770 2125.850 -12.590 2127.030 ;
        RECT -13.770 2124.250 -12.590 2125.430 ;
        RECT -13.770 2035.850 -12.590 2037.030 ;
        RECT -13.770 2034.250 -12.590 2035.430 ;
        RECT -13.770 1945.850 -12.590 1947.030 ;
        RECT -13.770 1944.250 -12.590 1945.430 ;
        RECT -13.770 1855.850 -12.590 1857.030 ;
        RECT -13.770 1854.250 -12.590 1855.430 ;
        RECT -13.770 1765.850 -12.590 1767.030 ;
        RECT -13.770 1764.250 -12.590 1765.430 ;
        RECT -13.770 1675.850 -12.590 1677.030 ;
        RECT -13.770 1674.250 -12.590 1675.430 ;
        RECT -13.770 1585.850 -12.590 1587.030 ;
        RECT -13.770 1584.250 -12.590 1585.430 ;
        RECT -13.770 1495.850 -12.590 1497.030 ;
        RECT -13.770 1494.250 -12.590 1495.430 ;
        RECT -13.770 1405.850 -12.590 1407.030 ;
        RECT -13.770 1404.250 -12.590 1405.430 ;
        RECT -13.770 1315.850 -12.590 1317.030 ;
        RECT -13.770 1314.250 -12.590 1315.430 ;
        RECT -13.770 1225.850 -12.590 1227.030 ;
        RECT -13.770 1224.250 -12.590 1225.430 ;
        RECT -13.770 1135.850 -12.590 1137.030 ;
        RECT -13.770 1134.250 -12.590 1135.430 ;
        RECT -13.770 1045.850 -12.590 1047.030 ;
        RECT -13.770 1044.250 -12.590 1045.430 ;
        RECT -13.770 955.850 -12.590 957.030 ;
        RECT -13.770 954.250 -12.590 955.430 ;
        RECT -13.770 865.850 -12.590 867.030 ;
        RECT -13.770 864.250 -12.590 865.430 ;
        RECT -13.770 775.850 -12.590 777.030 ;
        RECT -13.770 774.250 -12.590 775.430 ;
        RECT -13.770 685.850 -12.590 687.030 ;
        RECT -13.770 684.250 -12.590 685.430 ;
        RECT -13.770 595.850 -12.590 597.030 ;
        RECT -13.770 594.250 -12.590 595.430 ;
        RECT -13.770 505.850 -12.590 507.030 ;
        RECT -13.770 504.250 -12.590 505.430 ;
        RECT -13.770 415.850 -12.590 417.030 ;
        RECT -13.770 414.250 -12.590 415.430 ;
        RECT -13.770 325.850 -12.590 327.030 ;
        RECT -13.770 324.250 -12.590 325.430 ;
        RECT -13.770 235.850 -12.590 237.030 ;
        RECT -13.770 234.250 -12.590 235.430 ;
        RECT -13.770 145.850 -12.590 147.030 ;
        RECT -13.770 144.250 -12.590 145.430 ;
        RECT -13.770 55.850 -12.590 57.030 ;
        RECT -13.770 54.250 -12.590 55.430 ;
        RECT 2932.210 3475.850 2933.390 3477.030 ;
        RECT 2932.210 3474.250 2933.390 3475.430 ;
        RECT 2932.210 3385.850 2933.390 3387.030 ;
        RECT 2932.210 3384.250 2933.390 3385.430 ;
        RECT 2932.210 3295.850 2933.390 3297.030 ;
        RECT 2932.210 3294.250 2933.390 3295.430 ;
        RECT 2932.210 3205.850 2933.390 3207.030 ;
        RECT 2932.210 3204.250 2933.390 3205.430 ;
        RECT 2932.210 3115.850 2933.390 3117.030 ;
        RECT 2932.210 3114.250 2933.390 3115.430 ;
        RECT 2932.210 3025.850 2933.390 3027.030 ;
        RECT 2932.210 3024.250 2933.390 3025.430 ;
        RECT 2932.210 2935.850 2933.390 2937.030 ;
        RECT 2932.210 2934.250 2933.390 2935.430 ;
        RECT 2932.210 2845.850 2933.390 2847.030 ;
        RECT 2932.210 2844.250 2933.390 2845.430 ;
        RECT 2932.210 2755.850 2933.390 2757.030 ;
        RECT 2932.210 2754.250 2933.390 2755.430 ;
        RECT 2932.210 2665.850 2933.390 2667.030 ;
        RECT 2932.210 2664.250 2933.390 2665.430 ;
        RECT 2932.210 2575.850 2933.390 2577.030 ;
        RECT 2932.210 2574.250 2933.390 2575.430 ;
        RECT 2932.210 2485.850 2933.390 2487.030 ;
        RECT 2932.210 2484.250 2933.390 2485.430 ;
        RECT 2932.210 2395.850 2933.390 2397.030 ;
        RECT 2932.210 2394.250 2933.390 2395.430 ;
        RECT 2932.210 2305.850 2933.390 2307.030 ;
        RECT 2932.210 2304.250 2933.390 2305.430 ;
        RECT 2932.210 2215.850 2933.390 2217.030 ;
        RECT 2932.210 2214.250 2933.390 2215.430 ;
        RECT 2932.210 2125.850 2933.390 2127.030 ;
        RECT 2932.210 2124.250 2933.390 2125.430 ;
        RECT 2932.210 2035.850 2933.390 2037.030 ;
        RECT 2932.210 2034.250 2933.390 2035.430 ;
        RECT 2932.210 1945.850 2933.390 1947.030 ;
        RECT 2932.210 1944.250 2933.390 1945.430 ;
        RECT 2932.210 1855.850 2933.390 1857.030 ;
        RECT 2932.210 1854.250 2933.390 1855.430 ;
        RECT 2932.210 1765.850 2933.390 1767.030 ;
        RECT 2932.210 1764.250 2933.390 1765.430 ;
        RECT 2932.210 1675.850 2933.390 1677.030 ;
        RECT 2932.210 1674.250 2933.390 1675.430 ;
        RECT 2932.210 1585.850 2933.390 1587.030 ;
        RECT 2932.210 1584.250 2933.390 1585.430 ;
        RECT 2932.210 1495.850 2933.390 1497.030 ;
        RECT 2932.210 1494.250 2933.390 1495.430 ;
        RECT 2932.210 1405.850 2933.390 1407.030 ;
        RECT 2932.210 1404.250 2933.390 1405.430 ;
        RECT 2932.210 1315.850 2933.390 1317.030 ;
        RECT 2932.210 1314.250 2933.390 1315.430 ;
        RECT 2932.210 1225.850 2933.390 1227.030 ;
        RECT 2932.210 1224.250 2933.390 1225.430 ;
        RECT 2932.210 1135.850 2933.390 1137.030 ;
        RECT 2932.210 1134.250 2933.390 1135.430 ;
        RECT 2932.210 1045.850 2933.390 1047.030 ;
        RECT 2932.210 1044.250 2933.390 1045.430 ;
        RECT 2932.210 955.850 2933.390 957.030 ;
        RECT 2932.210 954.250 2933.390 955.430 ;
        RECT 2932.210 865.850 2933.390 867.030 ;
        RECT 2932.210 864.250 2933.390 865.430 ;
        RECT 2932.210 775.850 2933.390 777.030 ;
        RECT 2932.210 774.250 2933.390 775.430 ;
        RECT 2932.210 685.850 2933.390 687.030 ;
        RECT 2932.210 684.250 2933.390 685.430 ;
        RECT 2932.210 595.850 2933.390 597.030 ;
        RECT 2932.210 594.250 2933.390 595.430 ;
        RECT 2932.210 505.850 2933.390 507.030 ;
        RECT 2932.210 504.250 2933.390 505.430 ;
        RECT 2932.210 415.850 2933.390 417.030 ;
        RECT 2932.210 414.250 2933.390 415.430 ;
        RECT 2932.210 325.850 2933.390 327.030 ;
        RECT 2932.210 324.250 2933.390 325.430 ;
        RECT 2932.210 235.850 2933.390 237.030 ;
        RECT 2932.210 234.250 2933.390 235.430 ;
        RECT 2932.210 145.850 2933.390 147.030 ;
        RECT 2932.210 144.250 2933.390 145.430 ;
        RECT 2932.210 55.850 2933.390 57.030 ;
        RECT 2932.210 54.250 2933.390 55.430 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 49.930 -7.610 51.110 -6.430 ;
        RECT 49.930 -9.210 51.110 -8.030 ;
        RECT 139.930 -7.610 141.110 -6.430 ;
        RECT 139.930 -9.210 141.110 -8.030 ;
        RECT 229.930 -7.610 231.110 -6.430 ;
        RECT 229.930 -9.210 231.110 -8.030 ;
        RECT 319.930 -7.610 321.110 -6.430 ;
        RECT 319.930 -9.210 321.110 -8.030 ;
        RECT 409.930 -7.610 411.110 -6.430 ;
        RECT 409.930 -9.210 411.110 -8.030 ;
        RECT 499.930 -7.610 501.110 -6.430 ;
        RECT 499.930 -9.210 501.110 -8.030 ;
        RECT 589.930 -7.610 591.110 -6.430 ;
        RECT 589.930 -9.210 591.110 -8.030 ;
        RECT 679.930 -7.610 681.110 -6.430 ;
        RECT 679.930 -9.210 681.110 -8.030 ;
        RECT 769.930 -7.610 771.110 -6.430 ;
        RECT 769.930 -9.210 771.110 -8.030 ;
        RECT 859.930 -7.610 861.110 -6.430 ;
        RECT 859.930 -9.210 861.110 -8.030 ;
        RECT 949.930 -7.610 951.110 -6.430 ;
        RECT 949.930 -9.210 951.110 -8.030 ;
        RECT 1039.930 -7.610 1041.110 -6.430 ;
        RECT 1039.930 -9.210 1041.110 -8.030 ;
        RECT 1129.930 -7.610 1131.110 -6.430 ;
        RECT 1129.930 -9.210 1131.110 -8.030 ;
        RECT 1219.930 -7.610 1221.110 -6.430 ;
        RECT 1219.930 -9.210 1221.110 -8.030 ;
        RECT 1309.930 -7.610 1311.110 -6.430 ;
        RECT 1309.930 -9.210 1311.110 -8.030 ;
        RECT 1399.930 -7.610 1401.110 -6.430 ;
        RECT 1399.930 -9.210 1401.110 -8.030 ;
        RECT 1489.930 -7.610 1491.110 -6.430 ;
        RECT 1489.930 -9.210 1491.110 -8.030 ;
        RECT 1579.930 -7.610 1581.110 -6.430 ;
        RECT 1579.930 -9.210 1581.110 -8.030 ;
        RECT 1669.930 -7.610 1671.110 -6.430 ;
        RECT 1669.930 -9.210 1671.110 -8.030 ;
        RECT 1759.930 -7.610 1761.110 -6.430 ;
        RECT 1759.930 -9.210 1761.110 -8.030 ;
        RECT 1849.930 -7.610 1851.110 -6.430 ;
        RECT 1849.930 -9.210 1851.110 -8.030 ;
        RECT 1939.930 -7.610 1941.110 -6.430 ;
        RECT 1939.930 -9.210 1941.110 -8.030 ;
        RECT 2029.930 -7.610 2031.110 -6.430 ;
        RECT 2029.930 -9.210 2031.110 -8.030 ;
        RECT 2119.930 -7.610 2121.110 -6.430 ;
        RECT 2119.930 -9.210 2121.110 -8.030 ;
        RECT 2209.930 -7.610 2211.110 -6.430 ;
        RECT 2209.930 -9.210 2211.110 -8.030 ;
        RECT 2299.930 -7.610 2301.110 -6.430 ;
        RECT 2299.930 -9.210 2301.110 -8.030 ;
        RECT 2389.930 -7.610 2391.110 -6.430 ;
        RECT 2389.930 -9.210 2391.110 -8.030 ;
        RECT 2479.930 -7.610 2481.110 -6.430 ;
        RECT 2479.930 -9.210 2481.110 -8.030 ;
        RECT 2569.930 -7.610 2571.110 -6.430 ;
        RECT 2569.930 -9.210 2571.110 -8.030 ;
        RECT 2659.930 -7.610 2661.110 -6.430 ;
        RECT 2659.930 -9.210 2661.110 -8.030 ;
        RECT 2749.930 -7.610 2751.110 -6.430 ;
        RECT 2749.930 -9.210 2751.110 -8.030 ;
        RECT 2839.930 -7.610 2841.110 -6.430 ;
        RECT 2839.930 -9.210 2841.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 49.020 3529.000 52.020 3529.010 ;
        RECT 139.020 3529.000 142.020 3529.010 ;
        RECT 229.020 3529.000 232.020 3529.010 ;
        RECT 319.020 3529.000 322.020 3529.010 ;
        RECT 409.020 3529.000 412.020 3529.010 ;
        RECT 499.020 3529.000 502.020 3529.010 ;
        RECT 589.020 3529.000 592.020 3529.010 ;
        RECT 679.020 3529.000 682.020 3529.010 ;
        RECT 769.020 3529.000 772.020 3529.010 ;
        RECT 859.020 3529.000 862.020 3529.010 ;
        RECT 949.020 3529.000 952.020 3529.010 ;
        RECT 1039.020 3529.000 1042.020 3529.010 ;
        RECT 1129.020 3529.000 1132.020 3529.010 ;
        RECT 1219.020 3529.000 1222.020 3529.010 ;
        RECT 1309.020 3529.000 1312.020 3529.010 ;
        RECT 1399.020 3529.000 1402.020 3529.010 ;
        RECT 1489.020 3529.000 1492.020 3529.010 ;
        RECT 1579.020 3529.000 1582.020 3529.010 ;
        RECT 1669.020 3529.000 1672.020 3529.010 ;
        RECT 1759.020 3529.000 1762.020 3529.010 ;
        RECT 1849.020 3529.000 1852.020 3529.010 ;
        RECT 1939.020 3529.000 1942.020 3529.010 ;
        RECT 2029.020 3529.000 2032.020 3529.010 ;
        RECT 2119.020 3529.000 2122.020 3529.010 ;
        RECT 2209.020 3529.000 2212.020 3529.010 ;
        RECT 2299.020 3529.000 2302.020 3529.010 ;
        RECT 2389.020 3529.000 2392.020 3529.010 ;
        RECT 2479.020 3529.000 2482.020 3529.010 ;
        RECT 2569.020 3529.000 2572.020 3529.010 ;
        RECT 2659.020 3529.000 2662.020 3529.010 ;
        RECT 2749.020 3529.000 2752.020 3529.010 ;
        RECT 2839.020 3529.000 2842.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 49.020 3525.990 52.020 3526.000 ;
        RECT 139.020 3525.990 142.020 3526.000 ;
        RECT 229.020 3525.990 232.020 3526.000 ;
        RECT 319.020 3525.990 322.020 3526.000 ;
        RECT 409.020 3525.990 412.020 3526.000 ;
        RECT 499.020 3525.990 502.020 3526.000 ;
        RECT 589.020 3525.990 592.020 3526.000 ;
        RECT 679.020 3525.990 682.020 3526.000 ;
        RECT 769.020 3525.990 772.020 3526.000 ;
        RECT 859.020 3525.990 862.020 3526.000 ;
        RECT 949.020 3525.990 952.020 3526.000 ;
        RECT 1039.020 3525.990 1042.020 3526.000 ;
        RECT 1129.020 3525.990 1132.020 3526.000 ;
        RECT 1219.020 3525.990 1222.020 3526.000 ;
        RECT 1309.020 3525.990 1312.020 3526.000 ;
        RECT 1399.020 3525.990 1402.020 3526.000 ;
        RECT 1489.020 3525.990 1492.020 3526.000 ;
        RECT 1579.020 3525.990 1582.020 3526.000 ;
        RECT 1669.020 3525.990 1672.020 3526.000 ;
        RECT 1759.020 3525.990 1762.020 3526.000 ;
        RECT 1849.020 3525.990 1852.020 3526.000 ;
        RECT 1939.020 3525.990 1942.020 3526.000 ;
        RECT 2029.020 3525.990 2032.020 3526.000 ;
        RECT 2119.020 3525.990 2122.020 3526.000 ;
        RECT 2209.020 3525.990 2212.020 3526.000 ;
        RECT 2299.020 3525.990 2302.020 3526.000 ;
        RECT 2389.020 3525.990 2392.020 3526.000 ;
        RECT 2479.020 3525.990 2482.020 3526.000 ;
        RECT 2569.020 3525.990 2572.020 3526.000 ;
        RECT 2659.020 3525.990 2662.020 3526.000 ;
        RECT 2749.020 3525.990 2752.020 3526.000 ;
        RECT 2839.020 3525.990 2842.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3477.140 -11.680 3477.150 ;
        RECT 2931.300 3477.140 2934.300 3477.150 ;
        RECT -14.680 3474.140 13.700 3477.140 ;
        RECT 2906.300 3474.140 2934.300 3477.140 ;
        RECT -14.680 3474.130 -11.680 3474.140 ;
        RECT 2931.300 3474.130 2934.300 3474.140 ;
        RECT -14.680 3387.140 -11.680 3387.150 ;
        RECT 2931.300 3387.140 2934.300 3387.150 ;
        RECT -14.680 3384.140 13.700 3387.140 ;
        RECT 2906.300 3384.140 2934.300 3387.140 ;
        RECT -14.680 3384.130 -11.680 3384.140 ;
        RECT 2931.300 3384.130 2934.300 3384.140 ;
        RECT -14.680 3297.140 -11.680 3297.150 ;
        RECT 2931.300 3297.140 2934.300 3297.150 ;
        RECT -14.680 3294.140 13.700 3297.140 ;
        RECT 2906.300 3294.140 2934.300 3297.140 ;
        RECT -14.680 3294.130 -11.680 3294.140 ;
        RECT 2931.300 3294.130 2934.300 3294.140 ;
        RECT -14.680 3207.140 -11.680 3207.150 ;
        RECT 2931.300 3207.140 2934.300 3207.150 ;
        RECT -14.680 3204.140 13.700 3207.140 ;
        RECT 2906.300 3204.140 2934.300 3207.140 ;
        RECT -14.680 3204.130 -11.680 3204.140 ;
        RECT 2931.300 3204.130 2934.300 3204.140 ;
        RECT -14.680 3117.140 -11.680 3117.150 ;
        RECT 2931.300 3117.140 2934.300 3117.150 ;
        RECT -14.680 3114.140 13.700 3117.140 ;
        RECT 2906.300 3114.140 2934.300 3117.140 ;
        RECT -14.680 3114.130 -11.680 3114.140 ;
        RECT 2931.300 3114.130 2934.300 3114.140 ;
        RECT -14.680 3027.140 -11.680 3027.150 ;
        RECT 2931.300 3027.140 2934.300 3027.150 ;
        RECT -14.680 3024.140 13.700 3027.140 ;
        RECT 2906.300 3024.140 2934.300 3027.140 ;
        RECT -14.680 3024.130 -11.680 3024.140 ;
        RECT 2931.300 3024.130 2934.300 3024.140 ;
        RECT -14.680 2937.140 -11.680 2937.150 ;
        RECT 2931.300 2937.140 2934.300 2937.150 ;
        RECT -14.680 2934.140 13.700 2937.140 ;
        RECT 2906.300 2934.140 2934.300 2937.140 ;
        RECT -14.680 2934.130 -11.680 2934.140 ;
        RECT 2931.300 2934.130 2934.300 2934.140 ;
        RECT -14.680 2847.140 -11.680 2847.150 ;
        RECT 2931.300 2847.140 2934.300 2847.150 ;
        RECT -14.680 2844.140 13.700 2847.140 ;
        RECT 2906.300 2844.140 2934.300 2847.140 ;
        RECT -14.680 2844.130 -11.680 2844.140 ;
        RECT 2931.300 2844.130 2934.300 2844.140 ;
        RECT -14.680 2757.140 -11.680 2757.150 ;
        RECT 2931.300 2757.140 2934.300 2757.150 ;
        RECT -14.680 2754.140 13.700 2757.140 ;
        RECT 2906.300 2754.140 2934.300 2757.140 ;
        RECT -14.680 2754.130 -11.680 2754.140 ;
        RECT 2931.300 2754.130 2934.300 2754.140 ;
        RECT -14.680 2667.140 -11.680 2667.150 ;
        RECT 2931.300 2667.140 2934.300 2667.150 ;
        RECT -14.680 2664.140 13.700 2667.140 ;
        RECT 2906.300 2664.140 2934.300 2667.140 ;
        RECT -14.680 2664.130 -11.680 2664.140 ;
        RECT 2931.300 2664.130 2934.300 2664.140 ;
        RECT -14.680 2577.140 -11.680 2577.150 ;
        RECT 2931.300 2577.140 2934.300 2577.150 ;
        RECT -14.680 2574.140 13.700 2577.140 ;
        RECT 2906.300 2574.140 2934.300 2577.140 ;
        RECT -14.680 2574.130 -11.680 2574.140 ;
        RECT 2931.300 2574.130 2934.300 2574.140 ;
        RECT -14.680 2487.140 -11.680 2487.150 ;
        RECT 2931.300 2487.140 2934.300 2487.150 ;
        RECT -14.680 2484.140 13.700 2487.140 ;
        RECT 2906.300 2484.140 2934.300 2487.140 ;
        RECT -14.680 2484.130 -11.680 2484.140 ;
        RECT 2931.300 2484.130 2934.300 2484.140 ;
        RECT -14.680 2397.140 -11.680 2397.150 ;
        RECT 2931.300 2397.140 2934.300 2397.150 ;
        RECT -14.680 2394.140 13.700 2397.140 ;
        RECT 2906.300 2394.140 2934.300 2397.140 ;
        RECT -14.680 2394.130 -11.680 2394.140 ;
        RECT 2931.300 2394.130 2934.300 2394.140 ;
        RECT -14.680 2307.140 -11.680 2307.150 ;
        RECT 2931.300 2307.140 2934.300 2307.150 ;
        RECT -14.680 2304.140 13.700 2307.140 ;
        RECT 2906.300 2304.140 2934.300 2307.140 ;
        RECT -14.680 2304.130 -11.680 2304.140 ;
        RECT 2931.300 2304.130 2934.300 2304.140 ;
        RECT -14.680 2217.140 -11.680 2217.150 ;
        RECT 2931.300 2217.140 2934.300 2217.150 ;
        RECT -14.680 2214.140 13.700 2217.140 ;
        RECT 2906.300 2214.140 2934.300 2217.140 ;
        RECT -14.680 2214.130 -11.680 2214.140 ;
        RECT 2931.300 2214.130 2934.300 2214.140 ;
        RECT -14.680 2127.140 -11.680 2127.150 ;
        RECT 2931.300 2127.140 2934.300 2127.150 ;
        RECT -14.680 2124.140 13.700 2127.140 ;
        RECT 2906.300 2124.140 2934.300 2127.140 ;
        RECT -14.680 2124.130 -11.680 2124.140 ;
        RECT 2931.300 2124.130 2934.300 2124.140 ;
        RECT -14.680 2037.140 -11.680 2037.150 ;
        RECT 2931.300 2037.140 2934.300 2037.150 ;
        RECT -14.680 2034.140 13.700 2037.140 ;
        RECT 2906.300 2034.140 2934.300 2037.140 ;
        RECT -14.680 2034.130 -11.680 2034.140 ;
        RECT 2931.300 2034.130 2934.300 2034.140 ;
        RECT -14.680 1947.140 -11.680 1947.150 ;
        RECT 2931.300 1947.140 2934.300 1947.150 ;
        RECT -14.680 1944.140 13.700 1947.140 ;
        RECT 2906.300 1944.140 2934.300 1947.140 ;
        RECT -14.680 1944.130 -11.680 1944.140 ;
        RECT 2931.300 1944.130 2934.300 1944.140 ;
        RECT -14.680 1857.140 -11.680 1857.150 ;
        RECT 2931.300 1857.140 2934.300 1857.150 ;
        RECT -14.680 1854.140 13.700 1857.140 ;
        RECT 2906.300 1854.140 2934.300 1857.140 ;
        RECT -14.680 1854.130 -11.680 1854.140 ;
        RECT 2931.300 1854.130 2934.300 1854.140 ;
        RECT -14.680 1767.140 -11.680 1767.150 ;
        RECT 2931.300 1767.140 2934.300 1767.150 ;
        RECT -14.680 1764.140 13.700 1767.140 ;
        RECT 2906.300 1764.140 2934.300 1767.140 ;
        RECT -14.680 1764.130 -11.680 1764.140 ;
        RECT 2931.300 1764.130 2934.300 1764.140 ;
        RECT -14.680 1677.140 -11.680 1677.150 ;
        RECT 2931.300 1677.140 2934.300 1677.150 ;
        RECT -14.680 1674.140 13.700 1677.140 ;
        RECT 2906.300 1674.140 2934.300 1677.140 ;
        RECT -14.680 1674.130 -11.680 1674.140 ;
        RECT 2931.300 1674.130 2934.300 1674.140 ;
        RECT -14.680 1587.140 -11.680 1587.150 ;
        RECT 2931.300 1587.140 2934.300 1587.150 ;
        RECT -14.680 1584.140 13.700 1587.140 ;
        RECT 2906.300 1584.140 2934.300 1587.140 ;
        RECT -14.680 1584.130 -11.680 1584.140 ;
        RECT 2931.300 1584.130 2934.300 1584.140 ;
        RECT -14.680 1497.140 -11.680 1497.150 ;
        RECT 2931.300 1497.140 2934.300 1497.150 ;
        RECT -14.680 1494.140 13.700 1497.140 ;
        RECT 2906.300 1494.140 2934.300 1497.140 ;
        RECT -14.680 1494.130 -11.680 1494.140 ;
        RECT 2931.300 1494.130 2934.300 1494.140 ;
        RECT -14.680 1407.140 -11.680 1407.150 ;
        RECT 2931.300 1407.140 2934.300 1407.150 ;
        RECT -14.680 1404.140 13.700 1407.140 ;
        RECT 2906.300 1404.140 2934.300 1407.140 ;
        RECT -14.680 1404.130 -11.680 1404.140 ;
        RECT 2931.300 1404.130 2934.300 1404.140 ;
        RECT -14.680 1317.140 -11.680 1317.150 ;
        RECT 2931.300 1317.140 2934.300 1317.150 ;
        RECT -14.680 1314.140 13.700 1317.140 ;
        RECT 2906.300 1314.140 2934.300 1317.140 ;
        RECT -14.680 1314.130 -11.680 1314.140 ;
        RECT 2931.300 1314.130 2934.300 1314.140 ;
        RECT -14.680 1227.140 -11.680 1227.150 ;
        RECT 2931.300 1227.140 2934.300 1227.150 ;
        RECT -14.680 1224.140 13.700 1227.140 ;
        RECT 2906.300 1224.140 2934.300 1227.140 ;
        RECT -14.680 1224.130 -11.680 1224.140 ;
        RECT 2931.300 1224.130 2934.300 1224.140 ;
        RECT -14.680 1137.140 -11.680 1137.150 ;
        RECT 2931.300 1137.140 2934.300 1137.150 ;
        RECT -14.680 1134.140 13.700 1137.140 ;
        RECT 2906.300 1134.140 2934.300 1137.140 ;
        RECT -14.680 1134.130 -11.680 1134.140 ;
        RECT 2931.300 1134.130 2934.300 1134.140 ;
        RECT -14.680 1047.140 -11.680 1047.150 ;
        RECT 2931.300 1047.140 2934.300 1047.150 ;
        RECT -14.680 1044.140 13.700 1047.140 ;
        RECT 2906.300 1044.140 2934.300 1047.140 ;
        RECT -14.680 1044.130 -11.680 1044.140 ;
        RECT 2931.300 1044.130 2934.300 1044.140 ;
        RECT -14.680 957.140 -11.680 957.150 ;
        RECT 2931.300 957.140 2934.300 957.150 ;
        RECT -14.680 954.140 13.700 957.140 ;
        RECT 2906.300 954.140 2934.300 957.140 ;
        RECT -14.680 954.130 -11.680 954.140 ;
        RECT 2931.300 954.130 2934.300 954.140 ;
        RECT -14.680 867.140 -11.680 867.150 ;
        RECT 2931.300 867.140 2934.300 867.150 ;
        RECT -14.680 864.140 13.700 867.140 ;
        RECT 2906.300 864.140 2934.300 867.140 ;
        RECT -14.680 864.130 -11.680 864.140 ;
        RECT 2931.300 864.130 2934.300 864.140 ;
        RECT -14.680 777.140 -11.680 777.150 ;
        RECT 2931.300 777.140 2934.300 777.150 ;
        RECT -14.680 774.140 13.700 777.140 ;
        RECT 2906.300 774.140 2934.300 777.140 ;
        RECT -14.680 774.130 -11.680 774.140 ;
        RECT 2931.300 774.130 2934.300 774.140 ;
        RECT -14.680 687.140 -11.680 687.150 ;
        RECT 2931.300 687.140 2934.300 687.150 ;
        RECT -14.680 684.140 13.700 687.140 ;
        RECT 2906.300 684.140 2934.300 687.140 ;
        RECT -14.680 684.130 -11.680 684.140 ;
        RECT 2931.300 684.130 2934.300 684.140 ;
        RECT -14.680 597.140 -11.680 597.150 ;
        RECT 2931.300 597.140 2934.300 597.150 ;
        RECT -14.680 594.140 13.700 597.140 ;
        RECT 2906.300 594.140 2934.300 597.140 ;
        RECT -14.680 594.130 -11.680 594.140 ;
        RECT 2931.300 594.130 2934.300 594.140 ;
        RECT -14.680 507.140 -11.680 507.150 ;
        RECT 2931.300 507.140 2934.300 507.150 ;
        RECT -14.680 504.140 13.700 507.140 ;
        RECT 2906.300 504.140 2934.300 507.140 ;
        RECT -14.680 504.130 -11.680 504.140 ;
        RECT 2931.300 504.130 2934.300 504.140 ;
        RECT -14.680 417.140 -11.680 417.150 ;
        RECT 2931.300 417.140 2934.300 417.150 ;
        RECT -14.680 414.140 13.700 417.140 ;
        RECT 2906.300 414.140 2934.300 417.140 ;
        RECT -14.680 414.130 -11.680 414.140 ;
        RECT 2931.300 414.130 2934.300 414.140 ;
        RECT -14.680 327.140 -11.680 327.150 ;
        RECT 2931.300 327.140 2934.300 327.150 ;
        RECT -14.680 324.140 13.700 327.140 ;
        RECT 2906.300 324.140 2934.300 327.140 ;
        RECT -14.680 324.130 -11.680 324.140 ;
        RECT 2931.300 324.130 2934.300 324.140 ;
        RECT -14.680 237.140 -11.680 237.150 ;
        RECT 2931.300 237.140 2934.300 237.150 ;
        RECT -14.680 234.140 13.700 237.140 ;
        RECT 2906.300 234.140 2934.300 237.140 ;
        RECT -14.680 234.130 -11.680 234.140 ;
        RECT 2931.300 234.130 2934.300 234.140 ;
        RECT -14.680 147.140 -11.680 147.150 ;
        RECT 2931.300 147.140 2934.300 147.150 ;
        RECT -14.680 144.140 13.700 147.140 ;
        RECT 2906.300 144.140 2934.300 147.140 ;
        RECT -14.680 144.130 -11.680 144.140 ;
        RECT 2931.300 144.130 2934.300 144.140 ;
        RECT -14.680 57.140 -11.680 57.150 ;
        RECT 2931.300 57.140 2934.300 57.150 ;
        RECT -14.680 54.140 13.700 57.140 ;
        RECT 2906.300 54.140 2934.300 57.140 ;
        RECT -14.680 54.130 -11.680 54.140 ;
        RECT 2931.300 54.130 2934.300 54.140 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 49.020 -6.320 52.020 -6.310 ;
        RECT 139.020 -6.320 142.020 -6.310 ;
        RECT 229.020 -6.320 232.020 -6.310 ;
        RECT 319.020 -6.320 322.020 -6.310 ;
        RECT 409.020 -6.320 412.020 -6.310 ;
        RECT 499.020 -6.320 502.020 -6.310 ;
        RECT 589.020 -6.320 592.020 -6.310 ;
        RECT 679.020 -6.320 682.020 -6.310 ;
        RECT 769.020 -6.320 772.020 -6.310 ;
        RECT 859.020 -6.320 862.020 -6.310 ;
        RECT 949.020 -6.320 952.020 -6.310 ;
        RECT 1039.020 -6.320 1042.020 -6.310 ;
        RECT 1129.020 -6.320 1132.020 -6.310 ;
        RECT 1219.020 -6.320 1222.020 -6.310 ;
        RECT 1309.020 -6.320 1312.020 -6.310 ;
        RECT 1399.020 -6.320 1402.020 -6.310 ;
        RECT 1489.020 -6.320 1492.020 -6.310 ;
        RECT 1579.020 -6.320 1582.020 -6.310 ;
        RECT 1669.020 -6.320 1672.020 -6.310 ;
        RECT 1759.020 -6.320 1762.020 -6.310 ;
        RECT 1849.020 -6.320 1852.020 -6.310 ;
        RECT 1939.020 -6.320 1942.020 -6.310 ;
        RECT 2029.020 -6.320 2032.020 -6.310 ;
        RECT 2119.020 -6.320 2122.020 -6.310 ;
        RECT 2209.020 -6.320 2212.020 -6.310 ;
        RECT 2299.020 -6.320 2302.020 -6.310 ;
        RECT 2389.020 -6.320 2392.020 -6.310 ;
        RECT 2479.020 -6.320 2482.020 -6.310 ;
        RECT 2569.020 -6.320 2572.020 -6.310 ;
        RECT 2659.020 -6.320 2662.020 -6.310 ;
        RECT 2749.020 -6.320 2752.020 -6.310 ;
        RECT 2839.020 -6.320 2842.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 49.020 -9.330 52.020 -9.320 ;
        RECT 139.020 -9.330 142.020 -9.320 ;
        RECT 229.020 -9.330 232.020 -9.320 ;
        RECT 319.020 -9.330 322.020 -9.320 ;
        RECT 409.020 -9.330 412.020 -9.320 ;
        RECT 499.020 -9.330 502.020 -9.320 ;
        RECT 589.020 -9.330 592.020 -9.320 ;
        RECT 679.020 -9.330 682.020 -9.320 ;
        RECT 769.020 -9.330 772.020 -9.320 ;
        RECT 859.020 -9.330 862.020 -9.320 ;
        RECT 949.020 -9.330 952.020 -9.320 ;
        RECT 1039.020 -9.330 1042.020 -9.320 ;
        RECT 1129.020 -9.330 1132.020 -9.320 ;
        RECT 1219.020 -9.330 1222.020 -9.320 ;
        RECT 1309.020 -9.330 1312.020 -9.320 ;
        RECT 1399.020 -9.330 1402.020 -9.320 ;
        RECT 1489.020 -9.330 1492.020 -9.320 ;
        RECT 1579.020 -9.330 1582.020 -9.320 ;
        RECT 1669.020 -9.330 1672.020 -9.320 ;
        RECT 1759.020 -9.330 1762.020 -9.320 ;
        RECT 1849.020 -9.330 1852.020 -9.320 ;
        RECT 1939.020 -9.330 1942.020 -9.320 ;
        RECT 2029.020 -9.330 2032.020 -9.320 ;
        RECT 2119.020 -9.330 2122.020 -9.320 ;
        RECT 2209.020 -9.330 2212.020 -9.320 ;
        RECT 2299.020 -9.330 2302.020 -9.320 ;
        RECT 2389.020 -9.330 2392.020 -9.320 ;
        RECT 2479.020 -9.330 2482.020 -9.320 ;
        RECT 2569.020 -9.330 2572.020 -9.320 ;
        RECT 2659.020 -9.330 2662.020 -9.320 ;
        RECT 2749.020 -9.330 2752.020 -9.320 ;
        RECT 2839.020 -9.330 2842.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2902.020 3517.600 2905.020 3538.400 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2740.020 3517.600 2743.020 3547.800 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2758.020 3517.600 2761.020 3557.200 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met4 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
    END
  END vssa2
  OBS
      LAYER nwell ;
        RECT 5.330 3507.385 7.090 3508.990 ;
        RECT 2912.530 3507.385 2914.290 3508.990 ;
      LAYER pwell ;
        RECT 5.665 3505.995 5.835 3506.165 ;
        RECT 9.805 3505.995 9.975 3506.165 ;
        RECT 11.185 3505.995 11.355 3506.165 ;
        RECT 2909.185 3505.995 2909.355 3506.165 ;
        RECT 2910.565 3505.995 2910.735 3506.165 ;
        RECT 2913.785 3505.995 2913.955 3506.165 ;
      LAYER nwell ;
        RECT 5.330 3501.945 7.090 3504.775 ;
        RECT 9.470 3503.170 12.610 3504.775 ;
        RECT 2912.530 3501.945 2914.290 3504.775 ;
      LAYER pwell ;
        RECT 5.665 3500.555 5.835 3500.725 ;
        RECT 2913.785 3500.555 2913.955 3500.725 ;
      LAYER nwell ;
        RECT 5.330 3496.505 7.090 3499.335 ;
        RECT 2912.530 3496.505 2914.290 3499.335 ;
      LAYER pwell ;
        RECT 5.665 3495.115 5.835 3495.285 ;
        RECT 2913.785 3495.115 2913.955 3495.285 ;
      LAYER nwell ;
        RECT 5.330 3491.065 7.090 3493.895 ;
        RECT 2912.530 3491.065 2914.290 3493.895 ;
      LAYER pwell ;
        RECT 5.665 3489.675 5.835 3489.845 ;
        RECT 2913.785 3489.675 2913.955 3489.845 ;
      LAYER nwell ;
        RECT 5.330 3485.625 7.090 3488.455 ;
        RECT 2912.530 3485.625 2914.290 3488.455 ;
      LAYER pwell ;
        RECT 5.665 3484.235 5.835 3484.405 ;
        RECT 2913.785 3484.235 2913.955 3484.405 ;
      LAYER nwell ;
        RECT 5.330 3480.185 7.090 3483.015 ;
        RECT 2912.530 3480.185 2914.290 3483.015 ;
      LAYER pwell ;
        RECT 5.665 3478.795 5.835 3478.965 ;
        RECT 2913.785 3478.795 2913.955 3478.965 ;
      LAYER nwell ;
        RECT 5.330 3474.745 7.090 3477.575 ;
        RECT 2912.530 3474.745 2914.290 3477.575 ;
      LAYER pwell ;
        RECT 5.665 3473.355 5.835 3473.525 ;
        RECT 2913.785 3473.355 2913.955 3473.525 ;
      LAYER nwell ;
        RECT 5.330 3469.305 7.090 3472.135 ;
        RECT 2912.530 3469.305 2914.290 3472.135 ;
      LAYER pwell ;
        RECT 5.665 3467.915 5.835 3468.085 ;
        RECT 2913.785 3467.915 2913.955 3468.085 ;
      LAYER nwell ;
        RECT 5.330 3463.865 7.090 3466.695 ;
        RECT 2912.530 3463.865 2914.290 3466.695 ;
      LAYER pwell ;
        RECT 5.665 3462.475 5.835 3462.645 ;
        RECT 2913.785 3462.475 2913.955 3462.645 ;
      LAYER nwell ;
        RECT 5.330 3458.425 7.090 3461.255 ;
        RECT 2912.530 3458.425 2914.290 3461.255 ;
      LAYER pwell ;
        RECT 5.665 3457.035 5.835 3457.205 ;
        RECT 2913.785 3457.035 2913.955 3457.205 ;
      LAYER nwell ;
        RECT 5.330 3452.985 7.090 3455.815 ;
        RECT 2912.530 3452.985 2914.290 3455.815 ;
      LAYER pwell ;
        RECT 5.665 3451.595 5.835 3451.765 ;
        RECT 2913.785 3451.595 2913.955 3451.765 ;
      LAYER nwell ;
        RECT 5.330 3447.545 7.090 3450.375 ;
        RECT 2912.530 3447.545 2914.290 3450.375 ;
      LAYER pwell ;
        RECT 5.665 3446.155 5.835 3446.325 ;
        RECT 2913.785 3446.155 2913.955 3446.325 ;
      LAYER nwell ;
        RECT 5.330 3442.105 7.090 3444.935 ;
        RECT 2912.530 3442.105 2914.290 3444.935 ;
      LAYER pwell ;
        RECT 5.665 3440.715 5.835 3440.885 ;
        RECT 2913.785 3440.715 2913.955 3440.885 ;
      LAYER nwell ;
        RECT 5.330 3436.665 7.090 3439.495 ;
        RECT 2912.530 3436.665 2914.290 3439.495 ;
      LAYER pwell ;
        RECT 5.665 3435.275 5.835 3435.445 ;
        RECT 2913.785 3435.275 2913.955 3435.445 ;
      LAYER nwell ;
        RECT 5.330 3431.225 7.090 3434.055 ;
        RECT 2912.530 3431.225 2914.290 3434.055 ;
      LAYER pwell ;
        RECT 5.665 3429.835 5.835 3430.005 ;
        RECT 2913.785 3429.835 2913.955 3430.005 ;
      LAYER nwell ;
        RECT 5.330 3425.785 7.090 3428.615 ;
        RECT 2912.530 3425.785 2914.290 3428.615 ;
      LAYER pwell ;
        RECT 5.665 3424.395 5.835 3424.565 ;
        RECT 2913.785 3424.395 2913.955 3424.565 ;
      LAYER nwell ;
        RECT 5.330 3420.345 7.090 3423.175 ;
        RECT 2912.530 3420.345 2914.290 3423.175 ;
      LAYER pwell ;
        RECT 5.665 3418.955 5.835 3419.125 ;
        RECT 2913.785 3418.955 2913.955 3419.125 ;
      LAYER nwell ;
        RECT 5.330 3414.905 7.090 3417.735 ;
        RECT 2912.530 3414.905 2914.290 3417.735 ;
      LAYER pwell ;
        RECT 5.665 3413.515 5.835 3413.685 ;
        RECT 2913.785 3413.515 2913.955 3413.685 ;
      LAYER nwell ;
        RECT 5.330 3409.465 7.090 3412.295 ;
        RECT 2912.530 3409.465 2914.290 3412.295 ;
      LAYER pwell ;
        RECT 5.665 3408.075 5.835 3408.245 ;
        RECT 2913.785 3408.075 2913.955 3408.245 ;
      LAYER nwell ;
        RECT 5.330 3404.025 7.090 3406.855 ;
        RECT 2912.530 3404.025 2914.290 3406.855 ;
      LAYER pwell ;
        RECT 5.665 3402.635 5.835 3402.805 ;
        RECT 2909.185 3402.635 2909.355 3402.805 ;
        RECT 2913.785 3402.635 2913.955 3402.805 ;
      LAYER nwell ;
        RECT 5.330 3398.585 7.090 3401.415 ;
        RECT 2912.530 3398.585 2914.290 3401.415 ;
      LAYER pwell ;
        RECT 5.665 3397.195 5.835 3397.365 ;
        RECT 2913.785 3397.195 2913.955 3397.365 ;
      LAYER nwell ;
        RECT 5.330 3393.145 7.090 3395.975 ;
        RECT 2912.530 3393.145 2914.290 3395.975 ;
      LAYER pwell ;
        RECT 5.665 3391.755 5.835 3391.925 ;
        RECT 2913.785 3391.755 2913.955 3391.925 ;
      LAYER nwell ;
        RECT 5.330 3387.705 7.090 3390.535 ;
        RECT 2912.530 3387.705 2914.290 3390.535 ;
      LAYER pwell ;
        RECT 5.665 3386.315 5.835 3386.485 ;
        RECT 2913.785 3386.315 2913.955 3386.485 ;
      LAYER nwell ;
        RECT 5.330 3382.265 7.090 3385.095 ;
        RECT 2912.530 3382.265 2914.290 3385.095 ;
      LAYER pwell ;
        RECT 5.665 3380.875 5.835 3381.045 ;
        RECT 2913.785 3380.875 2913.955 3381.045 ;
      LAYER nwell ;
        RECT 5.330 3376.825 7.090 3379.655 ;
        RECT 2912.530 3376.825 2914.290 3379.655 ;
      LAYER pwell ;
        RECT 5.665 3375.435 5.835 3375.605 ;
        RECT 2913.785 3375.435 2913.955 3375.605 ;
      LAYER nwell ;
        RECT 5.330 3371.385 7.090 3374.215 ;
        RECT 2912.530 3371.385 2914.290 3374.215 ;
      LAYER pwell ;
        RECT 5.665 3369.995 5.835 3370.165 ;
        RECT 2913.785 3369.995 2913.955 3370.165 ;
      LAYER nwell ;
        RECT 5.330 3365.945 7.090 3368.775 ;
        RECT 2912.530 3365.945 2914.290 3368.775 ;
      LAYER pwell ;
        RECT 5.665 3364.555 5.835 3364.725 ;
        RECT 2910.565 3364.555 2910.735 3364.725 ;
        RECT 2913.785 3364.555 2913.955 3364.725 ;
      LAYER nwell ;
        RECT 5.330 3360.505 7.090 3363.335 ;
        RECT 2912.530 3360.505 2914.290 3363.335 ;
      LAYER pwell ;
        RECT 5.665 3359.115 5.835 3359.285 ;
        RECT 2913.785 3359.115 2913.955 3359.285 ;
      LAYER nwell ;
        RECT 5.330 3355.065 7.090 3357.895 ;
        RECT 2912.530 3355.065 2914.290 3357.895 ;
      LAYER pwell ;
        RECT 5.665 3353.675 5.835 3353.845 ;
        RECT 2913.785 3353.675 2913.955 3353.845 ;
      LAYER nwell ;
        RECT 5.330 3349.625 7.090 3352.455 ;
        RECT 2912.530 3349.625 2914.290 3352.455 ;
      LAYER pwell ;
        RECT 5.665 3348.235 5.835 3348.405 ;
        RECT 2913.785 3348.235 2913.955 3348.405 ;
      LAYER nwell ;
        RECT 5.330 3344.185 7.090 3347.015 ;
        RECT 2912.530 3344.185 2914.290 3347.015 ;
      LAYER pwell ;
        RECT 5.665 3342.795 5.835 3342.965 ;
        RECT 2913.785 3342.795 2913.955 3342.965 ;
      LAYER nwell ;
        RECT 5.330 3338.745 7.090 3341.575 ;
        RECT 2912.530 3338.745 2914.290 3341.575 ;
      LAYER pwell ;
        RECT 5.665 3337.355 5.835 3337.525 ;
        RECT 2913.785 3337.355 2913.955 3337.525 ;
      LAYER nwell ;
        RECT 5.330 3333.305 7.090 3336.135 ;
        RECT 2912.530 3333.305 2914.290 3336.135 ;
      LAYER pwell ;
        RECT 5.665 3331.915 5.835 3332.085 ;
        RECT 2913.785 3331.915 2913.955 3332.085 ;
      LAYER nwell ;
        RECT 5.330 3327.865 7.090 3330.695 ;
        RECT 2912.530 3327.865 2914.290 3330.695 ;
      LAYER pwell ;
        RECT 5.665 3326.475 5.835 3326.645 ;
        RECT 2913.785 3326.475 2913.955 3326.645 ;
      LAYER nwell ;
        RECT 5.330 3322.425 7.090 3325.255 ;
        RECT 2912.530 3322.425 2914.290 3325.255 ;
      LAYER pwell ;
        RECT 5.665 3321.035 5.835 3321.205 ;
        RECT 2913.785 3321.035 2913.955 3321.205 ;
      LAYER nwell ;
        RECT 5.330 3316.985 7.090 3319.815 ;
        RECT 2912.530 3316.985 2914.290 3319.815 ;
      LAYER pwell ;
        RECT 5.665 3315.595 5.835 3315.765 ;
        RECT 2913.785 3315.595 2913.955 3315.765 ;
      LAYER nwell ;
        RECT 5.330 3311.545 7.090 3314.375 ;
        RECT 2912.530 3311.545 2914.290 3314.375 ;
      LAYER pwell ;
        RECT 5.665 3310.155 5.835 3310.325 ;
        RECT 2913.785 3310.155 2913.955 3310.325 ;
      LAYER nwell ;
        RECT 5.330 3306.105 7.090 3308.935 ;
        RECT 2912.530 3306.105 2914.290 3308.935 ;
      LAYER pwell ;
        RECT 5.665 3304.715 5.835 3304.885 ;
        RECT 2913.785 3304.715 2913.955 3304.885 ;
      LAYER nwell ;
        RECT 5.330 3300.665 7.090 3303.495 ;
        RECT 2912.530 3300.665 2914.290 3303.495 ;
      LAYER pwell ;
        RECT 5.665 3299.275 5.835 3299.445 ;
        RECT 2913.785 3299.275 2913.955 3299.445 ;
      LAYER nwell ;
        RECT 5.330 3295.225 7.090 3298.055 ;
        RECT 2912.530 3295.225 2914.290 3298.055 ;
      LAYER pwell ;
        RECT 5.665 3293.835 5.835 3294.005 ;
        RECT 2913.785 3293.835 2913.955 3294.005 ;
      LAYER nwell ;
        RECT 5.330 3289.785 7.090 3292.615 ;
        RECT 2912.530 3289.785 2914.290 3292.615 ;
      LAYER pwell ;
        RECT 5.665 3288.395 5.835 3288.565 ;
        RECT 2913.785 3288.395 2913.955 3288.565 ;
      LAYER nwell ;
        RECT 5.330 3284.345 7.090 3287.175 ;
        RECT 2912.530 3284.345 2914.290 3287.175 ;
      LAYER pwell ;
        RECT 5.665 3282.955 5.835 3283.125 ;
        RECT 2913.785 3282.955 2913.955 3283.125 ;
      LAYER nwell ;
        RECT 5.330 3278.905 7.090 3281.735 ;
        RECT 2912.530 3278.905 2914.290 3281.735 ;
      LAYER pwell ;
        RECT 5.665 3277.515 5.835 3277.685 ;
        RECT 2913.785 3277.515 2913.955 3277.685 ;
      LAYER nwell ;
        RECT 5.330 3273.465 7.090 3276.295 ;
        RECT 2912.530 3273.465 2914.290 3276.295 ;
      LAYER pwell ;
        RECT 5.665 3272.075 5.835 3272.245 ;
        RECT 2913.785 3272.075 2913.955 3272.245 ;
      LAYER nwell ;
        RECT 5.330 3268.025 7.090 3270.855 ;
        RECT 2912.530 3268.025 2914.290 3270.855 ;
      LAYER pwell ;
        RECT 5.665 3266.635 5.835 3266.805 ;
        RECT 2913.785 3266.635 2913.955 3266.805 ;
      LAYER nwell ;
        RECT 5.330 3262.585 7.090 3265.415 ;
        RECT 2912.530 3262.585 2914.290 3265.415 ;
      LAYER pwell ;
        RECT 5.665 3261.195 5.835 3261.365 ;
        RECT 2913.785 3261.195 2913.955 3261.365 ;
      LAYER nwell ;
        RECT 5.330 3257.145 7.090 3259.975 ;
        RECT 2912.530 3257.145 2914.290 3259.975 ;
      LAYER pwell ;
        RECT 5.665 3255.755 5.835 3255.925 ;
        RECT 2913.785 3255.755 2913.955 3255.925 ;
      LAYER nwell ;
        RECT 5.330 3251.705 7.090 3254.535 ;
        RECT 2912.530 3251.705 2914.290 3254.535 ;
      LAYER pwell ;
        RECT 5.665 3250.315 5.835 3250.485 ;
        RECT 2913.785 3250.315 2913.955 3250.485 ;
      LAYER nwell ;
        RECT 5.330 3246.265 7.090 3249.095 ;
        RECT 2912.530 3246.265 2914.290 3249.095 ;
      LAYER pwell ;
        RECT 5.665 3244.875 5.835 3245.045 ;
        RECT 2913.785 3244.875 2913.955 3245.045 ;
      LAYER nwell ;
        RECT 5.330 3240.825 7.090 3243.655 ;
        RECT 2912.530 3240.825 2914.290 3243.655 ;
      LAYER pwell ;
        RECT 5.665 3239.435 5.835 3239.605 ;
        RECT 2913.785 3239.435 2913.955 3239.605 ;
      LAYER nwell ;
        RECT 5.330 3235.385 7.090 3238.215 ;
        RECT 2912.530 3235.385 2914.290 3238.215 ;
      LAYER pwell ;
        RECT 5.665 3233.995 5.835 3234.165 ;
        RECT 2913.785 3233.995 2913.955 3234.165 ;
      LAYER nwell ;
        RECT 5.330 3229.945 7.090 3232.775 ;
        RECT 2912.530 3229.945 2914.290 3232.775 ;
      LAYER pwell ;
        RECT 5.665 3228.555 5.835 3228.725 ;
        RECT 2913.785 3228.555 2913.955 3228.725 ;
      LAYER nwell ;
        RECT 5.330 3224.505 7.090 3227.335 ;
        RECT 8.550 3224.505 10.310 3226.110 ;
        RECT 2912.530 3224.505 2914.290 3227.335 ;
      LAYER pwell ;
        RECT 5.665 3223.115 5.835 3223.285 ;
        RECT 8.885 3223.115 9.055 3223.285 ;
        RECT 2913.785 3223.115 2913.955 3223.285 ;
      LAYER nwell ;
        RECT 5.330 3219.065 7.090 3221.895 ;
        RECT 2912.530 3219.065 2914.290 3221.895 ;
      LAYER pwell ;
        RECT 5.665 3217.675 5.835 3217.845 ;
        RECT 2913.785 3217.675 2913.955 3217.845 ;
      LAYER nwell ;
        RECT 5.330 3213.625 7.090 3216.455 ;
        RECT 2912.530 3213.625 2914.290 3216.455 ;
      LAYER pwell ;
        RECT 5.665 3212.235 5.835 3212.405 ;
        RECT 2913.785 3212.235 2913.955 3212.405 ;
      LAYER nwell ;
        RECT 5.330 3208.185 7.090 3211.015 ;
        RECT 2912.530 3208.185 2914.290 3211.015 ;
      LAYER pwell ;
        RECT 5.665 3206.795 5.835 3206.965 ;
        RECT 2913.785 3206.795 2913.955 3206.965 ;
      LAYER nwell ;
        RECT 5.330 3202.745 7.090 3205.575 ;
        RECT 2912.530 3202.745 2914.290 3205.575 ;
      LAYER pwell ;
        RECT 5.665 3201.355 5.835 3201.525 ;
        RECT 2910.565 3201.355 2910.735 3201.525 ;
        RECT 2913.785 3201.355 2913.955 3201.525 ;
      LAYER nwell ;
        RECT 5.330 3197.305 7.090 3200.135 ;
        RECT 2912.530 3197.305 2914.290 3200.135 ;
      LAYER pwell ;
        RECT 5.665 3195.915 5.835 3196.085 ;
        RECT 2913.785 3195.915 2913.955 3196.085 ;
      LAYER nwell ;
        RECT 5.330 3191.865 7.090 3194.695 ;
        RECT 2912.530 3191.865 2914.290 3194.695 ;
      LAYER pwell ;
        RECT 5.665 3190.475 5.835 3190.645 ;
        RECT 2913.785 3190.475 2913.955 3190.645 ;
      LAYER nwell ;
        RECT 5.330 3186.425 7.090 3189.255 ;
        RECT 2912.530 3186.425 2914.290 3189.255 ;
      LAYER pwell ;
        RECT 5.665 3185.035 5.835 3185.205 ;
        RECT 2913.785 3185.035 2913.955 3185.205 ;
      LAYER nwell ;
        RECT 5.330 3180.985 7.090 3183.815 ;
        RECT 2912.530 3180.985 2914.290 3183.815 ;
      LAYER pwell ;
        RECT 5.665 3179.595 5.835 3179.765 ;
        RECT 2913.785 3179.595 2913.955 3179.765 ;
      LAYER nwell ;
        RECT 5.330 3175.545 7.090 3178.375 ;
        RECT 2912.530 3175.545 2914.290 3178.375 ;
      LAYER pwell ;
        RECT 5.665 3174.155 5.835 3174.325 ;
        RECT 2913.785 3174.155 2913.955 3174.325 ;
      LAYER nwell ;
        RECT 5.330 3170.105 7.090 3172.935 ;
        RECT 2912.530 3170.105 2914.290 3172.935 ;
      LAYER pwell ;
        RECT 5.665 3168.715 5.835 3168.885 ;
        RECT 2913.785 3168.715 2913.955 3168.885 ;
      LAYER nwell ;
        RECT 5.330 3164.665 7.090 3167.495 ;
        RECT 2912.530 3164.665 2914.290 3167.495 ;
      LAYER pwell ;
        RECT 5.665 3163.275 5.835 3163.445 ;
        RECT 2913.785 3163.275 2913.955 3163.445 ;
      LAYER nwell ;
        RECT 5.330 3159.225 7.090 3162.055 ;
        RECT 2912.530 3159.225 2914.290 3162.055 ;
      LAYER pwell ;
        RECT 5.665 3157.835 5.835 3158.005 ;
        RECT 2913.785 3157.835 2913.955 3158.005 ;
      LAYER nwell ;
        RECT 5.330 3153.785 7.090 3156.615 ;
        RECT 2912.530 3153.785 2914.290 3156.615 ;
      LAYER pwell ;
        RECT 5.665 3152.395 5.835 3152.565 ;
        RECT 2913.785 3152.395 2913.955 3152.565 ;
      LAYER nwell ;
        RECT 5.330 3148.345 7.090 3151.175 ;
        RECT 2912.530 3148.345 2914.290 3151.175 ;
      LAYER pwell ;
        RECT 5.665 3146.955 5.835 3147.125 ;
        RECT 2913.785 3146.955 2913.955 3147.125 ;
      LAYER nwell ;
        RECT 5.330 3142.905 7.090 3145.735 ;
        RECT 2912.530 3142.905 2914.290 3145.735 ;
      LAYER pwell ;
        RECT 5.665 3141.515 5.835 3141.685 ;
        RECT 2913.785 3141.515 2913.955 3141.685 ;
      LAYER nwell ;
        RECT 5.330 3137.465 7.090 3140.295 ;
        RECT 2912.530 3137.465 2914.290 3140.295 ;
      LAYER pwell ;
        RECT 5.665 3136.075 5.835 3136.245 ;
        RECT 2913.785 3136.075 2913.955 3136.245 ;
      LAYER nwell ;
        RECT 5.330 3132.025 7.090 3134.855 ;
        RECT 2912.530 3132.025 2914.290 3134.855 ;
      LAYER pwell ;
        RECT 5.665 3130.635 5.835 3130.805 ;
        RECT 2913.785 3130.635 2913.955 3130.805 ;
      LAYER nwell ;
        RECT 5.330 3126.585 7.090 3129.415 ;
        RECT 2912.530 3126.585 2914.290 3129.415 ;
      LAYER pwell ;
        RECT 5.665 3125.195 5.835 3125.365 ;
        RECT 2913.785 3125.195 2913.955 3125.365 ;
      LAYER nwell ;
        RECT 5.330 3121.145 7.090 3123.975 ;
        RECT 2912.530 3121.145 2914.290 3123.975 ;
      LAYER pwell ;
        RECT 5.665 3119.755 5.835 3119.925 ;
        RECT 2913.785 3119.755 2913.955 3119.925 ;
      LAYER nwell ;
        RECT 5.330 3115.705 7.090 3118.535 ;
        RECT 2912.530 3115.705 2914.290 3118.535 ;
      LAYER pwell ;
        RECT 5.665 3114.315 5.835 3114.485 ;
        RECT 2913.785 3114.315 2913.955 3114.485 ;
      LAYER nwell ;
        RECT 5.330 3110.265 7.090 3113.095 ;
        RECT 2912.530 3110.265 2914.290 3113.095 ;
      LAYER pwell ;
        RECT 5.665 3108.875 5.835 3109.045 ;
        RECT 2913.785 3108.875 2913.955 3109.045 ;
      LAYER nwell ;
        RECT 5.330 3104.825 7.090 3107.655 ;
        RECT 2912.530 3104.825 2914.290 3107.655 ;
      LAYER pwell ;
        RECT 5.665 3103.435 5.835 3103.605 ;
        RECT 2913.785 3103.435 2913.955 3103.605 ;
      LAYER nwell ;
        RECT 5.330 3099.385 7.090 3102.215 ;
        RECT 2912.530 3099.385 2914.290 3102.215 ;
      LAYER pwell ;
        RECT 5.665 3097.995 5.835 3098.165 ;
        RECT 2909.185 3097.995 2909.355 3098.165 ;
        RECT 2913.785 3097.995 2913.955 3098.165 ;
      LAYER nwell ;
        RECT 5.330 3093.945 7.090 3096.775 ;
        RECT 2912.530 3093.945 2914.290 3096.775 ;
      LAYER pwell ;
        RECT 5.665 3092.555 5.835 3092.725 ;
        RECT 2913.785 3092.555 2913.955 3092.725 ;
      LAYER nwell ;
        RECT 5.330 3088.505 7.090 3091.335 ;
        RECT 2912.530 3088.505 2914.290 3091.335 ;
      LAYER pwell ;
        RECT 5.665 3087.115 5.835 3087.285 ;
        RECT 2913.785 3087.115 2913.955 3087.285 ;
      LAYER nwell ;
        RECT 5.330 3083.065 7.090 3085.895 ;
        RECT 2912.530 3083.065 2914.290 3085.895 ;
      LAYER pwell ;
        RECT 5.665 3081.675 5.835 3081.845 ;
        RECT 2913.785 3081.675 2913.955 3081.845 ;
      LAYER nwell ;
        RECT 5.330 3077.625 7.090 3080.455 ;
        RECT 2912.530 3077.625 2914.290 3080.455 ;
      LAYER pwell ;
        RECT 5.665 3076.235 5.835 3076.405 ;
        RECT 2913.785 3076.235 2913.955 3076.405 ;
      LAYER nwell ;
        RECT 5.330 3072.185 7.090 3075.015 ;
        RECT 2912.530 3072.185 2914.290 3075.015 ;
      LAYER pwell ;
        RECT 5.665 3070.795 5.835 3070.965 ;
        RECT 2913.785 3070.795 2913.955 3070.965 ;
      LAYER nwell ;
        RECT 5.330 3066.745 7.090 3069.575 ;
        RECT 2912.530 3066.745 2914.290 3069.575 ;
      LAYER pwell ;
        RECT 5.665 3065.355 5.835 3065.525 ;
        RECT 2913.785 3065.355 2913.955 3065.525 ;
      LAYER nwell ;
        RECT 5.330 3061.305 7.090 3064.135 ;
        RECT 2912.530 3061.305 2914.290 3064.135 ;
      LAYER pwell ;
        RECT 5.665 3059.915 5.835 3060.085 ;
        RECT 2913.785 3059.915 2913.955 3060.085 ;
      LAYER nwell ;
        RECT 5.330 3055.865 7.090 3058.695 ;
        RECT 2912.530 3055.865 2914.290 3058.695 ;
      LAYER pwell ;
        RECT 5.665 3054.475 5.835 3054.645 ;
        RECT 2913.785 3054.475 2913.955 3054.645 ;
      LAYER nwell ;
        RECT 5.330 3050.425 7.090 3053.255 ;
        RECT 2912.530 3050.425 2914.290 3053.255 ;
      LAYER pwell ;
        RECT 5.665 3049.035 5.835 3049.205 ;
        RECT 2913.785 3049.035 2913.955 3049.205 ;
      LAYER nwell ;
        RECT 5.330 3044.985 7.090 3047.815 ;
        RECT 2912.530 3044.985 2914.290 3047.815 ;
      LAYER pwell ;
        RECT 5.665 3043.595 5.835 3043.765 ;
        RECT 2913.785 3043.595 2913.955 3043.765 ;
      LAYER nwell ;
        RECT 5.330 3039.545 7.090 3042.375 ;
        RECT 2912.530 3039.545 2914.290 3042.375 ;
      LAYER pwell ;
        RECT 5.665 3038.155 5.835 3038.325 ;
        RECT 2913.785 3038.155 2913.955 3038.325 ;
      LAYER nwell ;
        RECT 5.330 3034.105 7.090 3036.935 ;
        RECT 2912.530 3034.105 2914.290 3036.935 ;
      LAYER pwell ;
        RECT 5.665 3032.715 5.835 3032.885 ;
        RECT 2913.785 3032.715 2913.955 3032.885 ;
      LAYER nwell ;
        RECT 5.330 3028.665 7.090 3031.495 ;
        RECT 2912.530 3028.665 2914.290 3031.495 ;
      LAYER pwell ;
        RECT 5.665 3027.275 5.835 3027.445 ;
        RECT 2913.785 3027.275 2913.955 3027.445 ;
      LAYER nwell ;
        RECT 5.330 3023.225 7.090 3026.055 ;
        RECT 2912.530 3023.225 2914.290 3026.055 ;
      LAYER pwell ;
        RECT 5.665 3021.835 5.835 3022.005 ;
        RECT 2913.785 3021.835 2913.955 3022.005 ;
      LAYER nwell ;
        RECT 5.330 3017.785 7.090 3020.615 ;
        RECT 2912.530 3017.785 2914.290 3020.615 ;
      LAYER pwell ;
        RECT 5.665 3016.395 5.835 3016.565 ;
        RECT 2913.785 3016.395 2913.955 3016.565 ;
      LAYER nwell ;
        RECT 5.330 3012.345 7.090 3015.175 ;
        RECT 8.550 3012.345 10.310 3013.950 ;
        RECT 2912.530 3012.345 2914.290 3015.175 ;
      LAYER pwell ;
        RECT 5.665 3010.955 5.835 3011.125 ;
        RECT 8.885 3010.955 9.055 3011.125 ;
        RECT 2913.785 3010.955 2913.955 3011.125 ;
      LAYER nwell ;
        RECT 5.330 3006.905 7.090 3009.735 ;
        RECT 2912.530 3006.905 2914.290 3009.735 ;
      LAYER pwell ;
        RECT 5.665 3005.515 5.835 3005.685 ;
        RECT 2913.785 3005.515 2913.955 3005.685 ;
      LAYER nwell ;
        RECT 5.330 3001.465 7.090 3004.295 ;
        RECT 2912.530 3001.465 2914.290 3004.295 ;
      LAYER pwell ;
        RECT 5.665 3000.075 5.835 3000.245 ;
        RECT 2913.785 3000.075 2913.955 3000.245 ;
      LAYER nwell ;
        RECT 5.330 2996.025 7.090 2998.855 ;
        RECT 2912.530 2996.025 2914.290 2998.855 ;
      LAYER pwell ;
        RECT 5.665 2994.635 5.835 2994.805 ;
        RECT 2913.785 2994.635 2913.955 2994.805 ;
      LAYER nwell ;
        RECT 5.330 2990.585 7.090 2993.415 ;
        RECT 2912.530 2990.585 2914.290 2993.415 ;
      LAYER pwell ;
        RECT 5.665 2989.195 5.835 2989.365 ;
        RECT 2913.785 2989.195 2913.955 2989.365 ;
      LAYER nwell ;
        RECT 5.330 2985.145 7.090 2987.975 ;
        RECT 2912.530 2985.145 2914.290 2987.975 ;
      LAYER pwell ;
        RECT 5.665 2983.755 5.835 2983.925 ;
        RECT 2913.785 2983.755 2913.955 2983.925 ;
      LAYER nwell ;
        RECT 5.330 2979.705 7.090 2982.535 ;
        RECT 2912.530 2979.705 2914.290 2982.535 ;
      LAYER pwell ;
        RECT 5.665 2978.315 5.835 2978.485 ;
        RECT 2913.785 2978.315 2913.955 2978.485 ;
      LAYER nwell ;
        RECT 5.330 2974.265 7.090 2977.095 ;
        RECT 2912.530 2974.265 2914.290 2977.095 ;
      LAYER pwell ;
        RECT 5.665 2972.875 5.835 2973.045 ;
        RECT 8.885 2972.875 9.055 2973.045 ;
        RECT 2913.785 2972.875 2913.955 2973.045 ;
      LAYER nwell ;
        RECT 5.330 2968.825 7.090 2971.655 ;
        RECT 8.550 2970.050 10.310 2971.655 ;
        RECT 2912.530 2968.825 2914.290 2971.655 ;
      LAYER pwell ;
        RECT 5.665 2967.435 5.835 2967.605 ;
        RECT 2913.785 2967.435 2913.955 2967.605 ;
      LAYER nwell ;
        RECT 5.330 2963.385 7.090 2966.215 ;
        RECT 2912.530 2963.385 2914.290 2966.215 ;
      LAYER pwell ;
        RECT 5.665 2961.995 5.835 2962.165 ;
        RECT 2913.785 2961.995 2913.955 2962.165 ;
      LAYER nwell ;
        RECT 5.330 2957.945 7.090 2960.775 ;
        RECT 2912.530 2957.945 2914.290 2960.775 ;
      LAYER pwell ;
        RECT 5.665 2956.555 5.835 2956.725 ;
        RECT 8.885 2956.555 9.055 2956.725 ;
        RECT 2913.785 2956.555 2913.955 2956.725 ;
      LAYER nwell ;
        RECT 5.330 2952.505 7.090 2955.335 ;
        RECT 8.550 2953.730 10.310 2955.335 ;
        RECT 2912.530 2952.505 2914.290 2955.335 ;
      LAYER pwell ;
        RECT 5.665 2951.115 5.835 2951.285 ;
        RECT 2913.785 2951.115 2913.955 2951.285 ;
      LAYER nwell ;
        RECT 5.330 2947.065 7.090 2949.895 ;
        RECT 2912.530 2947.065 2914.290 2949.895 ;
      LAYER pwell ;
        RECT 5.665 2945.675 5.835 2945.845 ;
        RECT 2913.785 2945.675 2913.955 2945.845 ;
      LAYER nwell ;
        RECT 5.330 2941.625 7.090 2944.455 ;
        RECT 2912.530 2941.625 2914.290 2944.455 ;
      LAYER pwell ;
        RECT 5.665 2940.235 5.835 2940.405 ;
        RECT 2913.785 2940.235 2913.955 2940.405 ;
      LAYER nwell ;
        RECT 5.330 2936.185 7.090 2939.015 ;
        RECT 2912.530 2936.185 2914.290 2939.015 ;
      LAYER pwell ;
        RECT 5.665 2934.795 5.835 2934.965 ;
        RECT 2913.785 2934.795 2913.955 2934.965 ;
      LAYER nwell ;
        RECT 5.330 2930.745 7.090 2933.575 ;
        RECT 2912.530 2930.745 2914.290 2933.575 ;
      LAYER pwell ;
        RECT 5.665 2929.355 5.835 2929.525 ;
        RECT 2913.785 2929.355 2913.955 2929.525 ;
      LAYER nwell ;
        RECT 5.330 2925.305 7.090 2928.135 ;
        RECT 2912.530 2925.305 2914.290 2928.135 ;
      LAYER pwell ;
        RECT 5.665 2923.915 5.835 2924.085 ;
        RECT 2913.785 2923.915 2913.955 2924.085 ;
      LAYER nwell ;
        RECT 5.330 2919.865 7.090 2922.695 ;
        RECT 2912.530 2919.865 2914.290 2922.695 ;
      LAYER pwell ;
        RECT 5.665 2918.475 5.835 2918.645 ;
        RECT 2913.785 2918.475 2913.955 2918.645 ;
      LAYER nwell ;
        RECT 5.330 2914.425 7.090 2917.255 ;
        RECT 2912.530 2914.425 2914.290 2917.255 ;
      LAYER pwell ;
        RECT 5.665 2913.035 5.835 2913.205 ;
        RECT 2910.565 2913.035 2910.735 2913.205 ;
        RECT 2913.785 2913.035 2913.955 2913.205 ;
      LAYER nwell ;
        RECT 5.330 2908.985 7.090 2911.815 ;
        RECT 2912.530 2908.985 2914.290 2911.815 ;
      LAYER pwell ;
        RECT 5.665 2907.595 5.835 2907.765 ;
        RECT 2913.785 2907.595 2913.955 2907.765 ;
      LAYER nwell ;
        RECT 5.330 2903.545 7.090 2906.375 ;
        RECT 2912.530 2903.545 2914.290 2906.375 ;
      LAYER pwell ;
        RECT 5.665 2902.155 5.835 2902.325 ;
        RECT 2913.785 2902.155 2913.955 2902.325 ;
      LAYER nwell ;
        RECT 5.330 2898.105 7.090 2900.935 ;
        RECT 2912.530 2898.105 2914.290 2900.935 ;
      LAYER pwell ;
        RECT 5.665 2896.715 5.835 2896.885 ;
        RECT 2913.785 2896.715 2913.955 2896.885 ;
      LAYER nwell ;
        RECT 5.330 2892.665 7.090 2895.495 ;
        RECT 2912.530 2892.665 2914.290 2895.495 ;
      LAYER pwell ;
        RECT 5.665 2891.275 5.835 2891.445 ;
        RECT 2913.785 2891.275 2913.955 2891.445 ;
      LAYER nwell ;
        RECT 5.330 2887.225 7.090 2890.055 ;
        RECT 2912.530 2887.225 2914.290 2890.055 ;
      LAYER pwell ;
        RECT 5.665 2885.835 5.835 2886.005 ;
        RECT 8.885 2885.835 9.055 2886.005 ;
        RECT 2913.785 2885.835 2913.955 2886.005 ;
      LAYER nwell ;
        RECT 5.330 2881.785 7.090 2884.615 ;
        RECT 8.550 2883.010 10.310 2884.615 ;
        RECT 2912.530 2881.785 2914.290 2884.615 ;
      LAYER pwell ;
        RECT 5.665 2880.395 5.835 2880.565 ;
        RECT 2913.785 2880.395 2913.955 2880.565 ;
      LAYER nwell ;
        RECT 5.330 2876.345 7.090 2879.175 ;
        RECT 2912.530 2876.345 2914.290 2879.175 ;
      LAYER pwell ;
        RECT 5.665 2874.955 5.835 2875.125 ;
        RECT 2913.785 2874.955 2913.955 2875.125 ;
      LAYER nwell ;
        RECT 5.330 2870.905 7.090 2873.735 ;
        RECT 8.550 2870.905 10.310 2872.510 ;
        RECT 2912.530 2870.905 2914.290 2873.735 ;
      LAYER pwell ;
        RECT 5.665 2869.515 5.835 2869.685 ;
        RECT 8.885 2869.515 9.055 2869.685 ;
        RECT 2913.785 2869.515 2913.955 2869.685 ;
      LAYER nwell ;
        RECT 5.330 2865.465 7.090 2868.295 ;
        RECT 2912.530 2865.465 2914.290 2868.295 ;
      LAYER pwell ;
        RECT 5.665 2864.075 5.835 2864.245 ;
        RECT 2913.785 2864.075 2913.955 2864.245 ;
      LAYER nwell ;
        RECT 5.330 2860.025 7.090 2862.855 ;
        RECT 2912.530 2860.025 2914.290 2862.855 ;
      LAYER pwell ;
        RECT 5.665 2858.635 5.835 2858.805 ;
        RECT 2913.785 2858.635 2913.955 2858.805 ;
      LAYER nwell ;
        RECT 5.330 2854.585 7.090 2857.415 ;
        RECT 2912.530 2854.585 2914.290 2857.415 ;
      LAYER pwell ;
        RECT 5.665 2853.195 5.835 2853.365 ;
        RECT 2913.785 2853.195 2913.955 2853.365 ;
      LAYER nwell ;
        RECT 5.330 2849.145 7.090 2851.975 ;
        RECT 2912.530 2849.145 2914.290 2851.975 ;
      LAYER pwell ;
        RECT 5.665 2847.755 5.835 2847.925 ;
        RECT 2913.785 2847.755 2913.955 2847.925 ;
      LAYER nwell ;
        RECT 5.330 2843.705 7.090 2846.535 ;
        RECT 2912.530 2843.705 2914.290 2846.535 ;
      LAYER pwell ;
        RECT 5.665 2842.315 5.835 2842.485 ;
        RECT 2913.785 2842.315 2913.955 2842.485 ;
      LAYER nwell ;
        RECT 5.330 2838.265 7.090 2841.095 ;
        RECT 2912.530 2838.265 2914.290 2841.095 ;
      LAYER pwell ;
        RECT 5.665 2836.875 5.835 2837.045 ;
        RECT 2913.785 2836.875 2913.955 2837.045 ;
      LAYER nwell ;
        RECT 5.330 2832.825 7.090 2835.655 ;
        RECT 2912.530 2832.825 2914.290 2835.655 ;
      LAYER pwell ;
        RECT 5.665 2831.435 5.835 2831.605 ;
        RECT 2913.785 2831.435 2913.955 2831.605 ;
      LAYER nwell ;
        RECT 5.330 2827.385 7.090 2830.215 ;
        RECT 2912.530 2827.385 2914.290 2830.215 ;
      LAYER pwell ;
        RECT 5.665 2825.995 5.835 2826.165 ;
        RECT 2913.785 2825.995 2913.955 2826.165 ;
      LAYER nwell ;
        RECT 5.330 2821.945 7.090 2824.775 ;
        RECT 2912.530 2821.945 2914.290 2824.775 ;
      LAYER pwell ;
        RECT 5.665 2820.555 5.835 2820.725 ;
        RECT 2913.785 2820.555 2913.955 2820.725 ;
      LAYER nwell ;
        RECT 5.330 2816.505 7.090 2819.335 ;
        RECT 2912.530 2816.505 2914.290 2819.335 ;
      LAYER pwell ;
        RECT 5.665 2815.115 5.835 2815.285 ;
        RECT 2913.785 2815.115 2913.955 2815.285 ;
      LAYER nwell ;
        RECT 5.330 2811.065 7.090 2813.895 ;
        RECT 2912.530 2811.065 2914.290 2813.895 ;
      LAYER pwell ;
        RECT 5.665 2809.675 5.835 2809.845 ;
        RECT 2913.785 2809.675 2913.955 2809.845 ;
      LAYER nwell ;
        RECT 5.330 2805.625 7.090 2808.455 ;
        RECT 2912.530 2805.625 2914.290 2808.455 ;
      LAYER pwell ;
        RECT 5.665 2804.235 5.835 2804.405 ;
        RECT 2913.785 2804.235 2913.955 2804.405 ;
      LAYER nwell ;
        RECT 5.330 2800.185 7.090 2803.015 ;
        RECT 2912.530 2800.185 2914.290 2803.015 ;
      LAYER pwell ;
        RECT 5.665 2798.795 5.835 2798.965 ;
        RECT 2913.785 2798.795 2913.955 2798.965 ;
      LAYER nwell ;
        RECT 5.330 2794.745 7.090 2797.575 ;
        RECT 2912.530 2794.745 2914.290 2797.575 ;
      LAYER pwell ;
        RECT 5.665 2793.355 5.835 2793.525 ;
        RECT 2913.785 2793.355 2913.955 2793.525 ;
      LAYER nwell ;
        RECT 5.330 2789.305 7.090 2792.135 ;
        RECT 2912.530 2789.305 2914.290 2792.135 ;
      LAYER pwell ;
        RECT 5.665 2787.915 5.835 2788.085 ;
        RECT 2913.785 2787.915 2913.955 2788.085 ;
      LAYER nwell ;
        RECT 5.330 2783.865 7.090 2786.695 ;
        RECT 2912.530 2783.865 2914.290 2786.695 ;
      LAYER pwell ;
        RECT 5.665 2782.475 5.835 2782.645 ;
        RECT 2913.785 2782.475 2913.955 2782.645 ;
      LAYER nwell ;
        RECT 5.330 2778.425 7.090 2781.255 ;
        RECT 2912.530 2778.425 2914.290 2781.255 ;
      LAYER pwell ;
        RECT 5.665 2777.035 5.835 2777.205 ;
        RECT 2909.185 2777.035 2909.355 2777.205 ;
        RECT 2913.785 2777.035 2913.955 2777.205 ;
      LAYER nwell ;
        RECT 5.330 2772.985 7.090 2775.815 ;
        RECT 2912.530 2772.985 2914.290 2775.815 ;
      LAYER pwell ;
        RECT 5.665 2771.595 5.835 2771.765 ;
        RECT 2913.785 2771.595 2913.955 2771.765 ;
      LAYER nwell ;
        RECT 5.330 2767.545 7.090 2770.375 ;
        RECT 2912.530 2767.545 2914.290 2770.375 ;
      LAYER pwell ;
        RECT 5.665 2766.155 5.835 2766.325 ;
        RECT 2913.785 2766.155 2913.955 2766.325 ;
      LAYER nwell ;
        RECT 5.330 2762.105 7.090 2764.935 ;
        RECT 2912.530 2762.105 2914.290 2764.935 ;
      LAYER pwell ;
        RECT 5.665 2760.715 5.835 2760.885 ;
        RECT 2913.785 2760.715 2913.955 2760.885 ;
      LAYER nwell ;
        RECT 5.330 2756.665 7.090 2759.495 ;
        RECT 2912.530 2756.665 2914.290 2759.495 ;
      LAYER pwell ;
        RECT 5.665 2755.275 5.835 2755.445 ;
        RECT 2913.785 2755.275 2913.955 2755.445 ;
      LAYER nwell ;
        RECT 5.330 2751.225 7.090 2754.055 ;
        RECT 2912.530 2751.225 2914.290 2754.055 ;
      LAYER pwell ;
        RECT 5.665 2749.835 5.835 2750.005 ;
        RECT 2913.785 2749.835 2913.955 2750.005 ;
      LAYER nwell ;
        RECT 5.330 2745.785 7.090 2748.615 ;
        RECT 2912.530 2745.785 2914.290 2748.615 ;
      LAYER pwell ;
        RECT 5.665 2744.395 5.835 2744.565 ;
        RECT 2913.785 2744.395 2913.955 2744.565 ;
      LAYER nwell ;
        RECT 5.330 2740.345 7.090 2743.175 ;
        RECT 2912.530 2740.345 2914.290 2743.175 ;
      LAYER pwell ;
        RECT 5.665 2738.955 5.835 2739.125 ;
        RECT 2913.785 2738.955 2913.955 2739.125 ;
      LAYER nwell ;
        RECT 5.330 2734.905 7.090 2737.735 ;
        RECT 2912.530 2734.905 2914.290 2737.735 ;
      LAYER pwell ;
        RECT 5.665 2733.515 5.835 2733.685 ;
        RECT 2913.785 2733.515 2913.955 2733.685 ;
      LAYER nwell ;
        RECT 5.330 2729.465 7.090 2732.295 ;
        RECT 2912.530 2729.465 2914.290 2732.295 ;
      LAYER pwell ;
        RECT 5.665 2728.075 5.835 2728.245 ;
        RECT 2913.785 2728.075 2913.955 2728.245 ;
      LAYER nwell ;
        RECT 5.330 2724.025 7.090 2726.855 ;
        RECT 2912.530 2724.025 2914.290 2726.855 ;
      LAYER pwell ;
        RECT 5.665 2722.635 5.835 2722.805 ;
        RECT 2913.785 2722.635 2913.955 2722.805 ;
      LAYER nwell ;
        RECT 5.330 2718.585 7.090 2721.415 ;
        RECT 2912.530 2718.585 2914.290 2721.415 ;
      LAYER pwell ;
        RECT 5.665 2717.195 5.835 2717.365 ;
        RECT 2913.785 2717.195 2913.955 2717.365 ;
      LAYER nwell ;
        RECT 5.330 2713.145 7.090 2715.975 ;
        RECT 2912.530 2713.145 2914.290 2715.975 ;
      LAYER pwell ;
        RECT 5.665 2711.755 5.835 2711.925 ;
        RECT 2913.785 2711.755 2913.955 2711.925 ;
      LAYER nwell ;
        RECT 5.330 2707.705 7.090 2710.535 ;
        RECT 2912.530 2707.705 2914.290 2710.535 ;
      LAYER pwell ;
        RECT 5.665 2706.315 5.835 2706.485 ;
        RECT 2913.785 2706.315 2913.955 2706.485 ;
      LAYER nwell ;
        RECT 5.330 2702.265 7.090 2705.095 ;
        RECT 2912.530 2702.265 2914.290 2705.095 ;
      LAYER pwell ;
        RECT 5.665 2700.875 5.835 2701.045 ;
        RECT 2913.785 2700.875 2913.955 2701.045 ;
      LAYER nwell ;
        RECT 5.330 2696.825 7.090 2699.655 ;
        RECT 2912.530 2696.825 2914.290 2699.655 ;
      LAYER pwell ;
        RECT 5.665 2695.435 5.835 2695.605 ;
        RECT 2913.785 2695.435 2913.955 2695.605 ;
      LAYER nwell ;
        RECT 5.330 2691.385 7.090 2694.215 ;
        RECT 2912.530 2691.385 2914.290 2694.215 ;
      LAYER pwell ;
        RECT 5.665 2689.995 5.835 2690.165 ;
        RECT 2913.785 2689.995 2913.955 2690.165 ;
      LAYER nwell ;
        RECT 5.330 2685.945 7.090 2688.775 ;
        RECT 2912.530 2685.945 2914.290 2688.775 ;
      LAYER pwell ;
        RECT 5.665 2684.555 5.835 2684.725 ;
        RECT 2913.785 2684.555 2913.955 2684.725 ;
      LAYER nwell ;
        RECT 5.330 2680.505 7.090 2683.335 ;
        RECT 2912.530 2680.505 2914.290 2683.335 ;
      LAYER pwell ;
        RECT 5.665 2679.115 5.835 2679.285 ;
        RECT 2913.785 2679.115 2913.955 2679.285 ;
      LAYER nwell ;
        RECT 5.330 2675.065 7.090 2677.895 ;
        RECT 2912.530 2675.065 2914.290 2677.895 ;
      LAYER pwell ;
        RECT 5.665 2673.675 5.835 2673.845 ;
        RECT 2913.785 2673.675 2913.955 2673.845 ;
      LAYER nwell ;
        RECT 5.330 2669.625 7.090 2672.455 ;
        RECT 2912.530 2669.625 2914.290 2672.455 ;
      LAYER pwell ;
        RECT 5.665 2668.235 5.835 2668.405 ;
        RECT 2913.785 2668.235 2913.955 2668.405 ;
      LAYER nwell ;
        RECT 5.330 2664.185 7.090 2667.015 ;
        RECT 2912.530 2664.185 2914.290 2667.015 ;
      LAYER pwell ;
        RECT 5.665 2662.795 5.835 2662.965 ;
        RECT 2913.785 2662.795 2913.955 2662.965 ;
      LAYER nwell ;
        RECT 5.330 2658.745 7.090 2661.575 ;
        RECT 2912.530 2658.745 2914.290 2661.575 ;
      LAYER pwell ;
        RECT 5.665 2657.355 5.835 2657.525 ;
        RECT 2913.785 2657.355 2913.955 2657.525 ;
      LAYER nwell ;
        RECT 5.330 2653.305 7.090 2656.135 ;
        RECT 2912.530 2653.305 2914.290 2656.135 ;
      LAYER pwell ;
        RECT 5.665 2651.915 5.835 2652.085 ;
        RECT 2913.785 2651.915 2913.955 2652.085 ;
      LAYER nwell ;
        RECT 5.330 2647.865 7.090 2650.695 ;
        RECT 2912.530 2647.865 2914.290 2650.695 ;
      LAYER pwell ;
        RECT 5.665 2646.475 5.835 2646.645 ;
        RECT 2913.785 2646.475 2913.955 2646.645 ;
      LAYER nwell ;
        RECT 5.330 2642.425 7.090 2645.255 ;
        RECT 2912.530 2642.425 2914.290 2645.255 ;
      LAYER pwell ;
        RECT 5.665 2641.035 5.835 2641.205 ;
        RECT 2913.785 2641.035 2913.955 2641.205 ;
      LAYER nwell ;
        RECT 5.330 2636.985 7.090 2639.815 ;
        RECT 2912.530 2636.985 2914.290 2639.815 ;
      LAYER pwell ;
        RECT 5.665 2635.595 5.835 2635.765 ;
        RECT 2913.785 2635.595 2913.955 2635.765 ;
      LAYER nwell ;
        RECT 5.330 2631.545 7.090 2634.375 ;
        RECT 2912.530 2631.545 2914.290 2634.375 ;
      LAYER pwell ;
        RECT 5.665 2630.155 5.835 2630.325 ;
        RECT 2909.185 2630.155 2909.355 2630.325 ;
        RECT 2913.785 2630.155 2913.955 2630.325 ;
      LAYER nwell ;
        RECT 5.330 2626.105 7.090 2628.935 ;
        RECT 2908.850 2627.330 2910.610 2628.935 ;
        RECT 2912.530 2626.105 2914.290 2628.935 ;
      LAYER pwell ;
        RECT 5.665 2624.715 5.835 2624.885 ;
        RECT 2913.785 2624.715 2913.955 2624.885 ;
      LAYER nwell ;
        RECT 5.330 2620.665 7.090 2623.495 ;
        RECT 2912.530 2620.665 2914.290 2623.495 ;
      LAYER pwell ;
        RECT 5.665 2619.275 5.835 2619.445 ;
        RECT 2913.785 2619.275 2913.955 2619.445 ;
      LAYER nwell ;
        RECT 5.330 2615.225 7.090 2618.055 ;
        RECT 2912.530 2615.225 2914.290 2618.055 ;
      LAYER pwell ;
        RECT 5.665 2613.835 5.835 2614.005 ;
        RECT 2913.785 2613.835 2913.955 2614.005 ;
      LAYER nwell ;
        RECT 5.330 2609.785 7.090 2612.615 ;
        RECT 2912.530 2609.785 2914.290 2612.615 ;
      LAYER pwell ;
        RECT 5.665 2608.395 5.835 2608.565 ;
        RECT 2913.785 2608.395 2913.955 2608.565 ;
      LAYER nwell ;
        RECT 5.330 2604.345 7.090 2607.175 ;
        RECT 2912.530 2604.345 2914.290 2607.175 ;
      LAYER pwell ;
        RECT 5.665 2602.955 5.835 2603.125 ;
        RECT 2909.185 2602.955 2909.355 2603.125 ;
        RECT 2913.785 2602.955 2913.955 2603.125 ;
      LAYER nwell ;
        RECT 5.330 2598.905 7.090 2601.735 ;
        RECT 2908.850 2600.130 2910.610 2601.735 ;
        RECT 2912.530 2598.905 2914.290 2601.735 ;
      LAYER pwell ;
        RECT 5.665 2597.515 5.835 2597.685 ;
        RECT 2913.785 2597.515 2913.955 2597.685 ;
      LAYER nwell ;
        RECT 5.330 2593.465 7.090 2596.295 ;
        RECT 2912.530 2593.465 2914.290 2596.295 ;
      LAYER pwell ;
        RECT 5.665 2592.075 5.835 2592.245 ;
        RECT 2913.785 2592.075 2913.955 2592.245 ;
      LAYER nwell ;
        RECT 5.330 2588.025 7.090 2590.855 ;
        RECT 2912.530 2588.025 2914.290 2590.855 ;
      LAYER pwell ;
        RECT 5.665 2586.635 5.835 2586.805 ;
        RECT 2913.785 2586.635 2913.955 2586.805 ;
      LAYER nwell ;
        RECT 5.330 2582.585 7.090 2585.415 ;
        RECT 2912.530 2582.585 2914.290 2585.415 ;
      LAYER pwell ;
        RECT 5.665 2581.195 5.835 2581.365 ;
        RECT 2913.785 2581.195 2913.955 2581.365 ;
      LAYER nwell ;
        RECT 5.330 2577.145 7.090 2579.975 ;
        RECT 2912.530 2577.145 2914.290 2579.975 ;
      LAYER pwell ;
        RECT 5.665 2575.755 5.835 2575.925 ;
        RECT 2913.785 2575.755 2913.955 2575.925 ;
      LAYER nwell ;
        RECT 5.330 2571.705 7.090 2574.535 ;
        RECT 2912.530 2571.705 2914.290 2574.535 ;
      LAYER pwell ;
        RECT 5.665 2570.315 5.835 2570.485 ;
        RECT 2913.785 2570.315 2913.955 2570.485 ;
      LAYER nwell ;
        RECT 5.330 2566.265 7.090 2569.095 ;
        RECT 2912.530 2566.265 2914.290 2569.095 ;
      LAYER pwell ;
        RECT 5.665 2564.875 5.835 2565.045 ;
        RECT 2913.785 2564.875 2913.955 2565.045 ;
      LAYER nwell ;
        RECT 5.330 2560.825 7.090 2563.655 ;
        RECT 2912.530 2560.825 2914.290 2563.655 ;
      LAYER pwell ;
        RECT 5.665 2559.435 5.835 2559.605 ;
        RECT 2913.785 2559.435 2913.955 2559.605 ;
      LAYER nwell ;
        RECT 5.330 2555.385 7.090 2558.215 ;
        RECT 2912.530 2555.385 2914.290 2558.215 ;
      LAYER pwell ;
        RECT 5.665 2553.995 5.835 2554.165 ;
        RECT 2913.785 2553.995 2913.955 2554.165 ;
      LAYER nwell ;
        RECT 5.330 2549.945 7.090 2552.775 ;
        RECT 2912.530 2549.945 2914.290 2552.775 ;
      LAYER pwell ;
        RECT 5.665 2548.555 5.835 2548.725 ;
        RECT 2913.785 2548.555 2913.955 2548.725 ;
      LAYER nwell ;
        RECT 5.330 2544.505 7.090 2547.335 ;
        RECT 2912.530 2544.505 2914.290 2547.335 ;
      LAYER pwell ;
        RECT 5.665 2543.115 5.835 2543.285 ;
        RECT 2913.785 2543.115 2913.955 2543.285 ;
      LAYER nwell ;
        RECT 5.330 2539.065 7.090 2541.895 ;
        RECT 2912.530 2539.065 2914.290 2541.895 ;
      LAYER pwell ;
        RECT 5.665 2537.675 5.835 2537.845 ;
        RECT 2913.785 2537.675 2913.955 2537.845 ;
      LAYER nwell ;
        RECT 5.330 2533.625 7.090 2536.455 ;
        RECT 2912.530 2533.625 2914.290 2536.455 ;
      LAYER pwell ;
        RECT 5.665 2532.235 5.835 2532.405 ;
        RECT 2913.785 2532.235 2913.955 2532.405 ;
      LAYER nwell ;
        RECT 5.330 2528.185 7.090 2531.015 ;
        RECT 2912.530 2528.185 2914.290 2531.015 ;
      LAYER pwell ;
        RECT 5.665 2526.795 5.835 2526.965 ;
        RECT 2913.785 2526.795 2913.955 2526.965 ;
      LAYER nwell ;
        RECT 5.330 2522.745 7.090 2525.575 ;
        RECT 2912.530 2522.745 2914.290 2525.575 ;
      LAYER pwell ;
        RECT 5.665 2521.355 5.835 2521.525 ;
        RECT 2913.785 2521.355 2913.955 2521.525 ;
      LAYER nwell ;
        RECT 5.330 2517.305 7.090 2520.135 ;
        RECT 2912.530 2517.305 2914.290 2520.135 ;
      LAYER pwell ;
        RECT 5.665 2515.915 5.835 2516.085 ;
        RECT 2913.785 2515.915 2913.955 2516.085 ;
      LAYER nwell ;
        RECT 5.330 2511.865 7.090 2514.695 ;
        RECT 2912.530 2511.865 2914.290 2514.695 ;
      LAYER pwell ;
        RECT 5.665 2510.475 5.835 2510.645 ;
        RECT 2913.785 2510.475 2913.955 2510.645 ;
      LAYER nwell ;
        RECT 5.330 2506.425 7.090 2509.255 ;
        RECT 2912.530 2506.425 2914.290 2509.255 ;
      LAYER pwell ;
        RECT 5.665 2505.035 5.835 2505.205 ;
        RECT 2913.785 2505.035 2913.955 2505.205 ;
      LAYER nwell ;
        RECT 5.330 2500.985 7.090 2503.815 ;
        RECT 8.550 2500.985 10.310 2502.590 ;
        RECT 2912.530 2500.985 2914.290 2503.815 ;
      LAYER pwell ;
        RECT 5.665 2499.595 5.835 2499.765 ;
        RECT 8.885 2499.595 9.055 2499.765 ;
        RECT 2913.785 2499.595 2913.955 2499.765 ;
      LAYER nwell ;
        RECT 5.330 2495.545 7.090 2498.375 ;
        RECT 2912.530 2495.545 2914.290 2498.375 ;
      LAYER pwell ;
        RECT 5.665 2494.155 5.835 2494.325 ;
        RECT 2913.785 2494.155 2913.955 2494.325 ;
      LAYER nwell ;
        RECT 5.330 2490.105 7.090 2492.935 ;
        RECT 2912.530 2490.105 2914.290 2492.935 ;
      LAYER pwell ;
        RECT 5.665 2488.715 5.835 2488.885 ;
        RECT 2913.785 2488.715 2913.955 2488.885 ;
      LAYER nwell ;
        RECT 5.330 2484.665 7.090 2487.495 ;
        RECT 2912.530 2484.665 2914.290 2487.495 ;
      LAYER pwell ;
        RECT 5.665 2483.275 5.835 2483.445 ;
        RECT 2913.785 2483.275 2913.955 2483.445 ;
      LAYER nwell ;
        RECT 5.330 2479.225 7.090 2482.055 ;
        RECT 2912.530 2479.225 2914.290 2482.055 ;
      LAYER pwell ;
        RECT 5.665 2477.835 5.835 2478.005 ;
        RECT 2913.785 2477.835 2913.955 2478.005 ;
      LAYER nwell ;
        RECT 5.330 2473.785 7.090 2476.615 ;
        RECT 2912.530 2473.785 2914.290 2476.615 ;
      LAYER pwell ;
        RECT 5.665 2472.395 5.835 2472.565 ;
        RECT 2913.785 2472.395 2913.955 2472.565 ;
      LAYER nwell ;
        RECT 5.330 2468.345 7.090 2471.175 ;
        RECT 2912.530 2468.345 2914.290 2471.175 ;
      LAYER pwell ;
        RECT 5.665 2466.955 5.835 2467.125 ;
        RECT 2913.785 2466.955 2913.955 2467.125 ;
      LAYER nwell ;
        RECT 5.330 2462.905 7.090 2465.735 ;
        RECT 2908.850 2462.905 2910.610 2464.510 ;
        RECT 2912.530 2462.905 2914.290 2465.735 ;
      LAYER pwell ;
        RECT 5.665 2461.515 5.835 2461.685 ;
        RECT 2909.185 2461.515 2909.355 2461.685 ;
        RECT 2913.785 2461.515 2913.955 2461.685 ;
      LAYER nwell ;
        RECT 5.330 2457.465 7.090 2460.295 ;
        RECT 2912.530 2457.465 2914.290 2460.295 ;
      LAYER pwell ;
        RECT 5.665 2456.075 5.835 2456.245 ;
        RECT 2913.785 2456.075 2913.955 2456.245 ;
      LAYER nwell ;
        RECT 5.330 2452.025 7.090 2454.855 ;
        RECT 2912.530 2452.025 2914.290 2454.855 ;
      LAYER pwell ;
        RECT 5.665 2450.635 5.835 2450.805 ;
        RECT 2913.785 2450.635 2913.955 2450.805 ;
      LAYER nwell ;
        RECT 5.330 2446.585 7.090 2449.415 ;
        RECT 2912.530 2446.585 2914.290 2449.415 ;
      LAYER pwell ;
        RECT 5.665 2445.195 5.835 2445.365 ;
        RECT 2913.785 2445.195 2913.955 2445.365 ;
      LAYER nwell ;
        RECT 5.330 2441.145 7.090 2443.975 ;
        RECT 2912.530 2441.145 2914.290 2443.975 ;
      LAYER pwell ;
        RECT 5.665 2439.755 5.835 2439.925 ;
        RECT 2913.785 2439.755 2913.955 2439.925 ;
      LAYER nwell ;
        RECT 5.330 2435.705 7.090 2438.535 ;
        RECT 2912.530 2435.705 2914.290 2438.535 ;
      LAYER pwell ;
        RECT 5.665 2434.315 5.835 2434.485 ;
        RECT 2909.185 2434.315 2909.355 2434.485 ;
        RECT 2913.785 2434.315 2913.955 2434.485 ;
      LAYER nwell ;
        RECT 5.330 2430.265 7.090 2433.095 ;
        RECT 2908.850 2431.490 2910.610 2433.095 ;
        RECT 2912.530 2430.265 2914.290 2433.095 ;
      LAYER pwell ;
        RECT 5.665 2428.875 5.835 2429.045 ;
        RECT 2913.785 2428.875 2913.955 2429.045 ;
      LAYER nwell ;
        RECT 5.330 2424.825 7.090 2427.655 ;
        RECT 2912.530 2424.825 2914.290 2427.655 ;
      LAYER pwell ;
        RECT 5.665 2423.435 5.835 2423.605 ;
        RECT 2913.785 2423.435 2913.955 2423.605 ;
      LAYER nwell ;
        RECT 5.330 2419.385 7.090 2422.215 ;
        RECT 2912.530 2419.385 2914.290 2422.215 ;
      LAYER pwell ;
        RECT 5.665 2417.995 5.835 2418.165 ;
        RECT 2913.785 2417.995 2913.955 2418.165 ;
      LAYER nwell ;
        RECT 5.330 2413.945 7.090 2416.775 ;
        RECT 2912.530 2413.945 2914.290 2416.775 ;
      LAYER pwell ;
        RECT 5.665 2412.555 5.835 2412.725 ;
        RECT 2913.785 2412.555 2913.955 2412.725 ;
      LAYER nwell ;
        RECT 5.330 2408.505 7.090 2411.335 ;
        RECT 2912.530 2408.505 2914.290 2411.335 ;
      LAYER pwell ;
        RECT 5.665 2407.115 5.835 2407.285 ;
        RECT 2913.785 2407.115 2913.955 2407.285 ;
      LAYER nwell ;
        RECT 5.330 2403.065 7.090 2405.895 ;
        RECT 2912.530 2403.065 2914.290 2405.895 ;
      LAYER pwell ;
        RECT 5.665 2401.675 5.835 2401.845 ;
        RECT 2913.785 2401.675 2913.955 2401.845 ;
      LAYER nwell ;
        RECT 5.330 2397.625 7.090 2400.455 ;
        RECT 2912.530 2397.625 2914.290 2400.455 ;
      LAYER pwell ;
        RECT 5.665 2396.235 5.835 2396.405 ;
        RECT 2913.785 2396.235 2913.955 2396.405 ;
      LAYER nwell ;
        RECT 5.330 2392.185 7.090 2395.015 ;
        RECT 2912.530 2392.185 2914.290 2395.015 ;
      LAYER pwell ;
        RECT 5.665 2390.795 5.835 2390.965 ;
        RECT 2913.785 2390.795 2913.955 2390.965 ;
      LAYER nwell ;
        RECT 5.330 2386.745 7.090 2389.575 ;
        RECT 2908.850 2386.745 2910.610 2388.350 ;
        RECT 2912.530 2386.745 2914.290 2389.575 ;
      LAYER pwell ;
        RECT 5.665 2385.355 5.835 2385.525 ;
        RECT 2909.185 2385.355 2909.355 2385.525 ;
        RECT 2913.785 2385.355 2913.955 2385.525 ;
      LAYER nwell ;
        RECT 5.330 2381.305 7.090 2384.135 ;
        RECT 8.550 2381.305 10.310 2382.910 ;
        RECT 2912.530 2381.305 2914.290 2384.135 ;
      LAYER pwell ;
        RECT 5.665 2379.915 5.835 2380.085 ;
        RECT 8.885 2379.915 9.055 2380.085 ;
        RECT 2913.785 2379.915 2913.955 2380.085 ;
      LAYER nwell ;
        RECT 5.330 2375.865 7.090 2378.695 ;
        RECT 2912.530 2375.865 2914.290 2378.695 ;
      LAYER pwell ;
        RECT 5.665 2374.475 5.835 2374.645 ;
        RECT 2913.785 2374.475 2913.955 2374.645 ;
      LAYER nwell ;
        RECT 5.330 2370.425 7.090 2373.255 ;
        RECT 2912.530 2370.425 2914.290 2373.255 ;
      LAYER pwell ;
        RECT 5.665 2369.035 5.835 2369.205 ;
        RECT 2913.785 2369.035 2913.955 2369.205 ;
      LAYER nwell ;
        RECT 5.330 2364.985 7.090 2367.815 ;
        RECT 2912.530 2364.985 2914.290 2367.815 ;
      LAYER pwell ;
        RECT 5.665 2363.595 5.835 2363.765 ;
        RECT 2913.785 2363.595 2913.955 2363.765 ;
      LAYER nwell ;
        RECT 5.330 2359.545 7.090 2362.375 ;
        RECT 2912.530 2359.545 2914.290 2362.375 ;
      LAYER pwell ;
        RECT 5.665 2358.155 5.835 2358.325 ;
        RECT 2913.785 2358.155 2913.955 2358.325 ;
      LAYER nwell ;
        RECT 5.330 2354.105 7.090 2356.935 ;
        RECT 2912.530 2354.105 2914.290 2356.935 ;
      LAYER pwell ;
        RECT 5.665 2352.715 5.835 2352.885 ;
        RECT 2913.785 2352.715 2913.955 2352.885 ;
      LAYER nwell ;
        RECT 5.330 2348.665 7.090 2351.495 ;
        RECT 2912.530 2348.665 2914.290 2351.495 ;
      LAYER pwell ;
        RECT 5.665 2347.275 5.835 2347.445 ;
        RECT 2913.785 2347.275 2913.955 2347.445 ;
      LAYER nwell ;
        RECT 5.330 2343.225 7.090 2346.055 ;
        RECT 2912.530 2343.225 2914.290 2346.055 ;
      LAYER pwell ;
        RECT 5.665 2341.835 5.835 2342.005 ;
        RECT 2913.785 2341.835 2913.955 2342.005 ;
      LAYER nwell ;
        RECT 5.330 2337.785 7.090 2340.615 ;
        RECT 2912.530 2337.785 2914.290 2340.615 ;
      LAYER pwell ;
        RECT 5.665 2336.395 5.835 2336.565 ;
        RECT 2913.785 2336.395 2913.955 2336.565 ;
      LAYER nwell ;
        RECT 5.330 2332.345 7.090 2335.175 ;
        RECT 2912.530 2332.345 2914.290 2335.175 ;
      LAYER pwell ;
        RECT 5.665 2330.955 5.835 2331.125 ;
        RECT 2913.785 2330.955 2913.955 2331.125 ;
      LAYER nwell ;
        RECT 5.330 2326.905 7.090 2329.735 ;
        RECT 2912.530 2326.905 2914.290 2329.735 ;
      LAYER pwell ;
        RECT 5.665 2325.515 5.835 2325.685 ;
        RECT 2913.785 2325.515 2913.955 2325.685 ;
      LAYER nwell ;
        RECT 5.330 2321.465 7.090 2324.295 ;
        RECT 2912.530 2321.465 2914.290 2324.295 ;
      LAYER pwell ;
        RECT 5.665 2320.075 5.835 2320.245 ;
        RECT 2913.785 2320.075 2913.955 2320.245 ;
      LAYER nwell ;
        RECT 5.330 2316.025 7.090 2318.855 ;
        RECT 2912.530 2316.025 2914.290 2318.855 ;
      LAYER pwell ;
        RECT 5.665 2314.635 5.835 2314.805 ;
        RECT 2913.785 2314.635 2913.955 2314.805 ;
      LAYER nwell ;
        RECT 5.330 2310.585 7.090 2313.415 ;
        RECT 2912.530 2310.585 2914.290 2313.415 ;
      LAYER pwell ;
        RECT 5.665 2309.195 5.835 2309.365 ;
        RECT 2913.785 2309.195 2913.955 2309.365 ;
      LAYER nwell ;
        RECT 5.330 2305.145 7.090 2307.975 ;
        RECT 2912.530 2305.145 2914.290 2307.975 ;
      LAYER pwell ;
        RECT 5.665 2303.755 5.835 2303.925 ;
        RECT 2913.785 2303.755 2913.955 2303.925 ;
      LAYER nwell ;
        RECT 5.330 2299.705 7.090 2302.535 ;
        RECT 2912.530 2299.705 2914.290 2302.535 ;
      LAYER pwell ;
        RECT 5.665 2298.315 5.835 2298.485 ;
        RECT 2913.785 2298.315 2913.955 2298.485 ;
      LAYER nwell ;
        RECT 5.330 2294.265 7.090 2297.095 ;
        RECT 2912.530 2294.265 2914.290 2297.095 ;
      LAYER pwell ;
        RECT 5.665 2292.875 5.835 2293.045 ;
        RECT 2913.785 2292.875 2913.955 2293.045 ;
      LAYER nwell ;
        RECT 5.330 2288.825 7.090 2291.655 ;
        RECT 2912.530 2288.825 2914.290 2291.655 ;
      LAYER pwell ;
        RECT 5.665 2287.435 5.835 2287.605 ;
        RECT 2913.785 2287.435 2913.955 2287.605 ;
      LAYER nwell ;
        RECT 5.330 2283.385 7.090 2286.215 ;
        RECT 2912.530 2283.385 2914.290 2286.215 ;
      LAYER pwell ;
        RECT 5.665 2281.995 5.835 2282.165 ;
        RECT 2913.785 2281.995 2913.955 2282.165 ;
      LAYER nwell ;
        RECT 5.330 2277.945 7.090 2280.775 ;
        RECT 2912.530 2277.945 2914.290 2280.775 ;
      LAYER pwell ;
        RECT 5.665 2276.555 5.835 2276.725 ;
        RECT 2913.785 2276.555 2913.955 2276.725 ;
      LAYER nwell ;
        RECT 5.330 2272.505 7.090 2275.335 ;
        RECT 2912.530 2272.505 2914.290 2275.335 ;
      LAYER pwell ;
        RECT 5.665 2271.115 5.835 2271.285 ;
        RECT 2913.785 2271.115 2913.955 2271.285 ;
      LAYER nwell ;
        RECT 5.330 2267.065 7.090 2269.895 ;
        RECT 2912.530 2267.065 2914.290 2269.895 ;
      LAYER pwell ;
        RECT 5.665 2265.675 5.835 2265.845 ;
        RECT 2909.185 2265.675 2909.355 2265.845 ;
        RECT 2913.785 2265.675 2913.955 2265.845 ;
      LAYER nwell ;
        RECT 5.330 2261.625 7.090 2264.455 ;
        RECT 2908.850 2262.850 2910.610 2264.455 ;
        RECT 2912.530 2261.625 2914.290 2264.455 ;
      LAYER pwell ;
        RECT 5.665 2260.235 5.835 2260.405 ;
        RECT 2913.785 2260.235 2913.955 2260.405 ;
      LAYER nwell ;
        RECT 5.330 2256.185 7.090 2259.015 ;
        RECT 2912.530 2256.185 2914.290 2259.015 ;
      LAYER pwell ;
        RECT 5.665 2254.795 5.835 2254.965 ;
        RECT 2913.785 2254.795 2913.955 2254.965 ;
      LAYER nwell ;
        RECT 5.330 2250.745 7.090 2253.575 ;
        RECT 2912.530 2250.745 2914.290 2253.575 ;
      LAYER pwell ;
        RECT 5.665 2249.355 5.835 2249.525 ;
        RECT 2913.785 2249.355 2913.955 2249.525 ;
      LAYER nwell ;
        RECT 5.330 2245.305 7.090 2248.135 ;
        RECT 2912.530 2245.305 2914.290 2248.135 ;
      LAYER pwell ;
        RECT 5.665 2243.915 5.835 2244.085 ;
        RECT 2913.785 2243.915 2913.955 2244.085 ;
      LAYER nwell ;
        RECT 5.330 2239.865 7.090 2242.695 ;
        RECT 2912.530 2239.865 2914.290 2242.695 ;
      LAYER pwell ;
        RECT 5.665 2238.475 5.835 2238.645 ;
        RECT 2913.785 2238.475 2913.955 2238.645 ;
      LAYER nwell ;
        RECT 5.330 2234.425 7.090 2237.255 ;
        RECT 2912.530 2234.425 2914.290 2237.255 ;
      LAYER pwell ;
        RECT 5.665 2233.035 5.835 2233.205 ;
        RECT 2913.785 2233.035 2913.955 2233.205 ;
      LAYER nwell ;
        RECT 5.330 2228.985 7.090 2231.815 ;
        RECT 2912.530 2228.985 2914.290 2231.815 ;
      LAYER pwell ;
        RECT 5.665 2227.595 5.835 2227.765 ;
        RECT 2913.785 2227.595 2913.955 2227.765 ;
      LAYER nwell ;
        RECT 5.330 2223.545 7.090 2226.375 ;
        RECT 2912.530 2223.545 2914.290 2226.375 ;
      LAYER pwell ;
        RECT 5.665 2222.155 5.835 2222.325 ;
        RECT 2913.785 2222.155 2913.955 2222.325 ;
      LAYER nwell ;
        RECT 5.330 2218.105 7.090 2220.935 ;
        RECT 2912.530 2218.105 2914.290 2220.935 ;
      LAYER pwell ;
        RECT 5.665 2216.715 5.835 2216.885 ;
        RECT 2913.785 2216.715 2913.955 2216.885 ;
      LAYER nwell ;
        RECT 5.330 2212.665 7.090 2215.495 ;
        RECT 2912.530 2212.665 2914.290 2215.495 ;
      LAYER pwell ;
        RECT 5.665 2211.275 5.835 2211.445 ;
        RECT 2913.785 2211.275 2913.955 2211.445 ;
      LAYER nwell ;
        RECT 5.330 2207.225 7.090 2210.055 ;
        RECT 2912.530 2207.225 2914.290 2210.055 ;
      LAYER pwell ;
        RECT 5.665 2205.835 5.835 2206.005 ;
        RECT 2913.785 2205.835 2913.955 2206.005 ;
      LAYER nwell ;
        RECT 5.330 2201.785 7.090 2204.615 ;
        RECT 2912.530 2201.785 2914.290 2204.615 ;
      LAYER pwell ;
        RECT 5.665 2200.395 5.835 2200.565 ;
        RECT 2913.785 2200.395 2913.955 2200.565 ;
      LAYER nwell ;
        RECT 5.330 2196.345 7.090 2199.175 ;
        RECT 2912.530 2196.345 2914.290 2199.175 ;
      LAYER pwell ;
        RECT 5.665 2194.955 5.835 2195.125 ;
        RECT 2913.785 2194.955 2913.955 2195.125 ;
      LAYER nwell ;
        RECT 5.330 2190.905 7.090 2193.735 ;
        RECT 2912.530 2190.905 2914.290 2193.735 ;
      LAYER pwell ;
        RECT 5.665 2189.515 5.835 2189.685 ;
        RECT 2913.785 2189.515 2913.955 2189.685 ;
      LAYER nwell ;
        RECT 5.330 2185.465 7.090 2188.295 ;
        RECT 2912.530 2185.465 2914.290 2188.295 ;
      LAYER pwell ;
        RECT 5.665 2184.075 5.835 2184.245 ;
        RECT 2913.785 2184.075 2913.955 2184.245 ;
      LAYER nwell ;
        RECT 5.330 2180.025 7.090 2182.855 ;
        RECT 2912.530 2180.025 2914.290 2182.855 ;
      LAYER pwell ;
        RECT 5.665 2178.635 5.835 2178.805 ;
        RECT 2913.785 2178.635 2913.955 2178.805 ;
      LAYER nwell ;
        RECT 5.330 2174.585 7.090 2177.415 ;
        RECT 2912.530 2174.585 2914.290 2177.415 ;
      LAYER pwell ;
        RECT 5.665 2173.195 5.835 2173.365 ;
        RECT 2913.785 2173.195 2913.955 2173.365 ;
      LAYER nwell ;
        RECT 5.330 2169.145 7.090 2171.975 ;
        RECT 2912.530 2169.145 2914.290 2171.975 ;
      LAYER pwell ;
        RECT 5.665 2167.755 5.835 2167.925 ;
        RECT 2913.785 2167.755 2913.955 2167.925 ;
      LAYER nwell ;
        RECT 5.330 2163.705 7.090 2166.535 ;
        RECT 2912.530 2163.705 2914.290 2166.535 ;
      LAYER pwell ;
        RECT 5.665 2162.315 5.835 2162.485 ;
        RECT 2913.785 2162.315 2913.955 2162.485 ;
      LAYER nwell ;
        RECT 5.330 2158.265 7.090 2161.095 ;
        RECT 2912.530 2158.265 2914.290 2161.095 ;
      LAYER pwell ;
        RECT 5.665 2156.875 5.835 2157.045 ;
        RECT 2913.785 2156.875 2913.955 2157.045 ;
      LAYER nwell ;
        RECT 5.330 2152.825 7.090 2155.655 ;
        RECT 2912.530 2152.825 2914.290 2155.655 ;
      LAYER pwell ;
        RECT 5.665 2151.435 5.835 2151.605 ;
        RECT 2913.785 2151.435 2913.955 2151.605 ;
      LAYER nwell ;
        RECT 5.330 2147.385 7.090 2150.215 ;
        RECT 2912.530 2147.385 2914.290 2150.215 ;
      LAYER pwell ;
        RECT 5.665 2145.995 5.835 2146.165 ;
        RECT 2913.785 2145.995 2913.955 2146.165 ;
      LAYER nwell ;
        RECT 5.330 2141.945 7.090 2144.775 ;
        RECT 2912.530 2141.945 2914.290 2144.775 ;
      LAYER pwell ;
        RECT 5.665 2140.555 5.835 2140.725 ;
        RECT 2913.785 2140.555 2913.955 2140.725 ;
      LAYER nwell ;
        RECT 5.330 2136.505 7.090 2139.335 ;
        RECT 2912.530 2136.505 2914.290 2139.335 ;
      LAYER pwell ;
        RECT 5.665 2135.115 5.835 2135.285 ;
        RECT 2913.785 2135.115 2913.955 2135.285 ;
      LAYER nwell ;
        RECT 5.330 2131.065 7.090 2133.895 ;
        RECT 2912.530 2131.065 2914.290 2133.895 ;
      LAYER pwell ;
        RECT 5.665 2129.675 5.835 2129.845 ;
        RECT 2913.785 2129.675 2913.955 2129.845 ;
      LAYER nwell ;
        RECT 5.330 2125.625 7.090 2128.455 ;
        RECT 2912.530 2125.625 2914.290 2128.455 ;
      LAYER pwell ;
        RECT 5.665 2124.235 5.835 2124.405 ;
        RECT 2913.785 2124.235 2913.955 2124.405 ;
      LAYER nwell ;
        RECT 5.330 2120.185 7.090 2123.015 ;
        RECT 2912.530 2120.185 2914.290 2123.015 ;
      LAYER pwell ;
        RECT 5.665 2118.795 5.835 2118.965 ;
        RECT 2909.185 2118.795 2909.355 2118.965 ;
        RECT 2913.785 2118.795 2913.955 2118.965 ;
      LAYER nwell ;
        RECT 5.330 2114.745 7.090 2117.575 ;
        RECT 2908.850 2115.970 2910.610 2117.575 ;
        RECT 2912.530 2114.745 2914.290 2117.575 ;
      LAYER pwell ;
        RECT 5.665 2113.355 5.835 2113.525 ;
        RECT 2913.785 2113.355 2913.955 2113.525 ;
      LAYER nwell ;
        RECT 5.330 2109.305 7.090 2112.135 ;
        RECT 2912.530 2109.305 2914.290 2112.135 ;
      LAYER pwell ;
        RECT 5.665 2107.915 5.835 2108.085 ;
        RECT 2913.785 2107.915 2913.955 2108.085 ;
      LAYER nwell ;
        RECT 5.330 2103.865 7.090 2106.695 ;
        RECT 2912.530 2103.865 2914.290 2106.695 ;
      LAYER pwell ;
        RECT 5.665 2102.475 5.835 2102.645 ;
        RECT 2913.785 2102.475 2913.955 2102.645 ;
      LAYER nwell ;
        RECT 5.330 2098.425 7.090 2101.255 ;
        RECT 2912.530 2098.425 2914.290 2101.255 ;
      LAYER pwell ;
        RECT 5.665 2097.035 5.835 2097.205 ;
        RECT 2913.785 2097.035 2913.955 2097.205 ;
      LAYER nwell ;
        RECT 5.330 2092.985 7.090 2095.815 ;
        RECT 2912.530 2092.985 2914.290 2095.815 ;
      LAYER pwell ;
        RECT 5.665 2091.595 5.835 2091.765 ;
        RECT 2913.785 2091.595 2913.955 2091.765 ;
      LAYER nwell ;
        RECT 5.330 2087.545 7.090 2090.375 ;
        RECT 2912.530 2087.545 2914.290 2090.375 ;
      LAYER pwell ;
        RECT 5.665 2086.155 5.835 2086.325 ;
        RECT 2913.785 2086.155 2913.955 2086.325 ;
      LAYER nwell ;
        RECT 5.330 2082.105 7.090 2084.935 ;
        RECT 2912.530 2082.105 2914.290 2084.935 ;
      LAYER pwell ;
        RECT 5.665 2080.715 5.835 2080.885 ;
        RECT 2913.785 2080.715 2913.955 2080.885 ;
      LAYER nwell ;
        RECT 5.330 2076.665 7.090 2079.495 ;
        RECT 2912.530 2076.665 2914.290 2079.495 ;
      LAYER pwell ;
        RECT 5.665 2075.275 5.835 2075.445 ;
        RECT 2913.785 2075.275 2913.955 2075.445 ;
      LAYER nwell ;
        RECT 5.330 2071.225 7.090 2074.055 ;
        RECT 2912.530 2071.225 2914.290 2074.055 ;
      LAYER pwell ;
        RECT 5.665 2069.835 5.835 2070.005 ;
        RECT 2913.785 2069.835 2913.955 2070.005 ;
      LAYER nwell ;
        RECT 5.330 2065.785 7.090 2068.615 ;
        RECT 2912.530 2065.785 2914.290 2068.615 ;
      LAYER pwell ;
        RECT 5.665 2064.395 5.835 2064.565 ;
        RECT 2913.785 2064.395 2913.955 2064.565 ;
      LAYER nwell ;
        RECT 5.330 2060.345 7.090 2063.175 ;
        RECT 2912.530 2060.345 2914.290 2063.175 ;
      LAYER pwell ;
        RECT 5.665 2058.955 5.835 2059.125 ;
        RECT 2913.785 2058.955 2913.955 2059.125 ;
      LAYER nwell ;
        RECT 5.330 2054.905 7.090 2057.735 ;
        RECT 2912.530 2054.905 2914.290 2057.735 ;
      LAYER pwell ;
        RECT 5.665 2053.515 5.835 2053.685 ;
        RECT 2913.785 2053.515 2913.955 2053.685 ;
      LAYER nwell ;
        RECT 5.330 2049.465 7.090 2052.295 ;
        RECT 2912.530 2049.465 2914.290 2052.295 ;
      LAYER pwell ;
        RECT 5.665 2048.075 5.835 2048.245 ;
        RECT 2913.785 2048.075 2913.955 2048.245 ;
      LAYER nwell ;
        RECT 5.330 2044.025 7.090 2046.855 ;
        RECT 2912.530 2044.025 2914.290 2046.855 ;
      LAYER pwell ;
        RECT 5.665 2042.635 5.835 2042.805 ;
        RECT 2913.785 2042.635 2913.955 2042.805 ;
      LAYER nwell ;
        RECT 5.330 2038.585 7.090 2041.415 ;
        RECT 2912.530 2038.585 2914.290 2041.415 ;
      LAYER pwell ;
        RECT 5.665 2037.195 5.835 2037.365 ;
        RECT 2913.785 2037.195 2913.955 2037.365 ;
      LAYER nwell ;
        RECT 5.330 2033.145 7.090 2035.975 ;
        RECT 2912.530 2033.145 2914.290 2035.975 ;
      LAYER pwell ;
        RECT 5.665 2031.755 5.835 2031.925 ;
        RECT 2913.785 2031.755 2913.955 2031.925 ;
      LAYER nwell ;
        RECT 5.330 2027.705 7.090 2030.535 ;
        RECT 2912.530 2027.705 2914.290 2030.535 ;
      LAYER pwell ;
        RECT 5.665 2026.315 5.835 2026.485 ;
        RECT 2913.785 2026.315 2913.955 2026.485 ;
      LAYER nwell ;
        RECT 5.330 2022.265 7.090 2025.095 ;
        RECT 2912.530 2022.265 2914.290 2025.095 ;
      LAYER pwell ;
        RECT 5.665 2020.875 5.835 2021.045 ;
        RECT 2913.785 2020.875 2913.955 2021.045 ;
      LAYER nwell ;
        RECT 5.330 2016.825 7.090 2019.655 ;
        RECT 2912.530 2016.825 2914.290 2019.655 ;
      LAYER pwell ;
        RECT 5.665 2015.435 5.835 2015.605 ;
        RECT 2913.785 2015.435 2913.955 2015.605 ;
      LAYER nwell ;
        RECT 5.330 2011.385 7.090 2014.215 ;
        RECT 2912.530 2011.385 2914.290 2014.215 ;
      LAYER pwell ;
        RECT 5.665 2009.995 5.835 2010.165 ;
        RECT 2913.785 2009.995 2913.955 2010.165 ;
      LAYER nwell ;
        RECT 5.330 2005.945 7.090 2008.775 ;
        RECT 2912.530 2005.945 2914.290 2008.775 ;
      LAYER pwell ;
        RECT 5.665 2004.555 5.835 2004.725 ;
        RECT 2913.785 2004.555 2913.955 2004.725 ;
      LAYER nwell ;
        RECT 5.330 2000.505 7.090 2003.335 ;
        RECT 2912.530 2000.505 2914.290 2003.335 ;
      LAYER pwell ;
        RECT 5.665 1999.115 5.835 1999.285 ;
        RECT 2913.785 1999.115 2913.955 1999.285 ;
      LAYER nwell ;
        RECT 5.330 1995.065 7.090 1997.895 ;
        RECT 2912.530 1995.065 2914.290 1997.895 ;
      LAYER pwell ;
        RECT 5.665 1993.675 5.835 1993.845 ;
        RECT 2913.785 1993.675 2913.955 1993.845 ;
      LAYER nwell ;
        RECT 5.330 1989.625 7.090 1992.455 ;
        RECT 2912.530 1989.625 2914.290 1992.455 ;
      LAYER pwell ;
        RECT 5.665 1988.235 5.835 1988.405 ;
        RECT 2913.785 1988.235 2913.955 1988.405 ;
      LAYER nwell ;
        RECT 5.330 1984.185 7.090 1987.015 ;
        RECT 8.550 1984.185 10.310 1985.790 ;
        RECT 2912.530 1984.185 2914.290 1987.015 ;
      LAYER pwell ;
        RECT 5.665 1982.795 5.835 1982.965 ;
        RECT 8.885 1982.795 9.055 1982.965 ;
        RECT 2913.785 1982.795 2913.955 1982.965 ;
      LAYER nwell ;
        RECT 5.330 1978.745 7.090 1981.575 ;
        RECT 2912.530 1978.745 2914.290 1981.575 ;
      LAYER pwell ;
        RECT 5.665 1977.355 5.835 1977.525 ;
        RECT 2913.785 1977.355 2913.955 1977.525 ;
      LAYER nwell ;
        RECT 5.330 1973.305 7.090 1976.135 ;
        RECT 2912.530 1973.305 2914.290 1976.135 ;
      LAYER pwell ;
        RECT 5.665 1971.915 5.835 1972.085 ;
        RECT 2913.785 1971.915 2913.955 1972.085 ;
      LAYER nwell ;
        RECT 5.330 1967.865 7.090 1970.695 ;
        RECT 2912.530 1967.865 2914.290 1970.695 ;
      LAYER pwell ;
        RECT 5.665 1966.475 5.835 1966.645 ;
        RECT 2913.785 1966.475 2913.955 1966.645 ;
      LAYER nwell ;
        RECT 5.330 1962.425 7.090 1965.255 ;
        RECT 2912.530 1962.425 2914.290 1965.255 ;
      LAYER pwell ;
        RECT 5.665 1961.035 5.835 1961.205 ;
        RECT 2913.785 1961.035 2913.955 1961.205 ;
      LAYER nwell ;
        RECT 5.330 1956.985 7.090 1959.815 ;
        RECT 2912.530 1956.985 2914.290 1959.815 ;
      LAYER pwell ;
        RECT 5.665 1955.595 5.835 1955.765 ;
        RECT 8.885 1955.595 9.055 1955.765 ;
        RECT 2913.785 1955.595 2913.955 1955.765 ;
      LAYER nwell ;
        RECT 5.330 1951.545 7.090 1954.375 ;
        RECT 8.550 1952.770 10.310 1954.375 ;
        RECT 2912.530 1951.545 2914.290 1954.375 ;
      LAYER pwell ;
        RECT 5.665 1950.155 5.835 1950.325 ;
        RECT 2913.785 1950.155 2913.955 1950.325 ;
      LAYER nwell ;
        RECT 5.330 1946.105 7.090 1948.935 ;
        RECT 2912.530 1946.105 2914.290 1948.935 ;
      LAYER pwell ;
        RECT 5.665 1944.715 5.835 1944.885 ;
        RECT 2913.785 1944.715 2913.955 1944.885 ;
      LAYER nwell ;
        RECT 5.330 1940.665 7.090 1943.495 ;
        RECT 2912.530 1940.665 2914.290 1943.495 ;
      LAYER pwell ;
        RECT 5.665 1939.275 5.835 1939.445 ;
        RECT 2913.785 1939.275 2913.955 1939.445 ;
      LAYER nwell ;
        RECT 5.330 1935.225 7.090 1938.055 ;
        RECT 2908.850 1935.225 2910.610 1936.830 ;
        RECT 2912.530 1935.225 2914.290 1938.055 ;
      LAYER pwell ;
        RECT 5.665 1933.835 5.835 1934.005 ;
        RECT 2909.185 1933.835 2909.355 1934.005 ;
        RECT 2913.785 1933.835 2913.955 1934.005 ;
      LAYER nwell ;
        RECT 5.330 1929.785 7.090 1932.615 ;
        RECT 2912.530 1929.785 2914.290 1932.615 ;
      LAYER pwell ;
        RECT 5.665 1928.395 5.835 1928.565 ;
        RECT 2913.785 1928.395 2913.955 1928.565 ;
      LAYER nwell ;
        RECT 5.330 1924.345 7.090 1927.175 ;
        RECT 2912.530 1924.345 2914.290 1927.175 ;
      LAYER pwell ;
        RECT 5.665 1922.955 5.835 1923.125 ;
        RECT 2913.785 1922.955 2913.955 1923.125 ;
      LAYER nwell ;
        RECT 5.330 1918.905 7.090 1921.735 ;
        RECT 2912.530 1918.905 2914.290 1921.735 ;
      LAYER pwell ;
        RECT 5.665 1917.515 5.835 1917.685 ;
        RECT 2913.785 1917.515 2913.955 1917.685 ;
      LAYER nwell ;
        RECT 5.330 1913.465 7.090 1916.295 ;
        RECT 2912.530 1913.465 2914.290 1916.295 ;
      LAYER pwell ;
        RECT 5.665 1912.075 5.835 1912.245 ;
        RECT 2913.785 1912.075 2913.955 1912.245 ;
      LAYER nwell ;
        RECT 5.330 1908.025 7.090 1910.855 ;
        RECT 2912.530 1908.025 2914.290 1910.855 ;
      LAYER pwell ;
        RECT 5.665 1906.635 5.835 1906.805 ;
        RECT 2913.785 1906.635 2913.955 1906.805 ;
      LAYER nwell ;
        RECT 5.330 1902.585 7.090 1905.415 ;
        RECT 2912.530 1902.585 2914.290 1905.415 ;
      LAYER pwell ;
        RECT 5.665 1901.195 5.835 1901.365 ;
        RECT 2913.785 1901.195 2913.955 1901.365 ;
      LAYER nwell ;
        RECT 5.330 1897.145 7.090 1899.975 ;
        RECT 2912.530 1897.145 2914.290 1899.975 ;
      LAYER pwell ;
        RECT 5.665 1895.755 5.835 1895.925 ;
        RECT 2913.785 1895.755 2913.955 1895.925 ;
      LAYER nwell ;
        RECT 5.330 1891.705 7.090 1894.535 ;
        RECT 2912.530 1891.705 2914.290 1894.535 ;
      LAYER pwell ;
        RECT 5.665 1890.315 5.835 1890.485 ;
        RECT 2913.785 1890.315 2913.955 1890.485 ;
      LAYER nwell ;
        RECT 5.330 1886.265 7.090 1889.095 ;
        RECT 2912.530 1886.265 2914.290 1889.095 ;
      LAYER pwell ;
        RECT 5.665 1884.875 5.835 1885.045 ;
        RECT 2913.785 1884.875 2913.955 1885.045 ;
      LAYER nwell ;
        RECT 5.330 1880.825 7.090 1883.655 ;
        RECT 2912.530 1880.825 2914.290 1883.655 ;
      LAYER pwell ;
        RECT 5.665 1879.435 5.835 1879.605 ;
        RECT 2913.785 1879.435 2913.955 1879.605 ;
      LAYER nwell ;
        RECT 5.330 1875.385 7.090 1878.215 ;
        RECT 2912.530 1875.385 2914.290 1878.215 ;
      LAYER pwell ;
        RECT 5.665 1873.995 5.835 1874.165 ;
        RECT 2913.785 1873.995 2913.955 1874.165 ;
      LAYER nwell ;
        RECT 5.330 1869.945 7.090 1872.775 ;
        RECT 2912.530 1869.945 2914.290 1872.775 ;
      LAYER pwell ;
        RECT 5.665 1868.555 5.835 1868.725 ;
        RECT 2913.785 1868.555 2913.955 1868.725 ;
      LAYER nwell ;
        RECT 5.330 1864.505 7.090 1867.335 ;
        RECT 2912.530 1864.505 2914.290 1867.335 ;
      LAYER pwell ;
        RECT 5.665 1863.115 5.835 1863.285 ;
        RECT 2913.785 1863.115 2913.955 1863.285 ;
      LAYER nwell ;
        RECT 5.330 1859.065 7.090 1861.895 ;
        RECT 2912.530 1859.065 2914.290 1861.895 ;
      LAYER pwell ;
        RECT 5.665 1857.675 5.835 1857.845 ;
        RECT 2913.785 1857.675 2913.955 1857.845 ;
      LAYER nwell ;
        RECT 5.330 1853.625 7.090 1856.455 ;
        RECT 2912.530 1853.625 2914.290 1856.455 ;
      LAYER pwell ;
        RECT 5.665 1852.235 5.835 1852.405 ;
        RECT 2913.785 1852.235 2913.955 1852.405 ;
      LAYER nwell ;
        RECT 5.330 1848.185 7.090 1851.015 ;
        RECT 2912.530 1848.185 2914.290 1851.015 ;
      LAYER pwell ;
        RECT 5.665 1846.795 5.835 1846.965 ;
        RECT 2913.785 1846.795 2913.955 1846.965 ;
      LAYER nwell ;
        RECT 5.330 1842.745 7.090 1845.575 ;
        RECT 2912.530 1842.745 2914.290 1845.575 ;
      LAYER pwell ;
        RECT 5.665 1841.355 5.835 1841.525 ;
        RECT 2913.785 1841.355 2913.955 1841.525 ;
      LAYER nwell ;
        RECT 5.330 1837.305 7.090 1840.135 ;
        RECT 2912.530 1837.305 2914.290 1840.135 ;
      LAYER pwell ;
        RECT 5.665 1835.915 5.835 1836.085 ;
        RECT 2913.785 1835.915 2913.955 1836.085 ;
      LAYER nwell ;
        RECT 5.330 1831.865 7.090 1834.695 ;
        RECT 2912.530 1831.865 2914.290 1834.695 ;
      LAYER pwell ;
        RECT 5.665 1830.475 5.835 1830.645 ;
        RECT 2913.785 1830.475 2913.955 1830.645 ;
      LAYER nwell ;
        RECT 5.330 1826.425 7.090 1829.255 ;
        RECT 2912.530 1826.425 2914.290 1829.255 ;
      LAYER pwell ;
        RECT 5.665 1825.035 5.835 1825.205 ;
        RECT 2913.785 1825.035 2913.955 1825.205 ;
      LAYER nwell ;
        RECT 5.330 1820.985 7.090 1823.815 ;
        RECT 2912.530 1820.985 2914.290 1823.815 ;
      LAYER pwell ;
        RECT 5.665 1819.595 5.835 1819.765 ;
        RECT 2913.785 1819.595 2913.955 1819.765 ;
      LAYER nwell ;
        RECT 5.330 1815.545 7.090 1818.375 ;
        RECT 2912.530 1815.545 2914.290 1818.375 ;
      LAYER pwell ;
        RECT 5.665 1814.155 5.835 1814.325 ;
        RECT 2913.785 1814.155 2913.955 1814.325 ;
      LAYER nwell ;
        RECT 5.330 1810.105 7.090 1812.935 ;
        RECT 2912.530 1810.105 2914.290 1812.935 ;
      LAYER pwell ;
        RECT 5.665 1808.715 5.835 1808.885 ;
        RECT 2913.785 1808.715 2913.955 1808.885 ;
      LAYER nwell ;
        RECT 5.330 1804.665 7.090 1807.495 ;
        RECT 2912.530 1804.665 2914.290 1807.495 ;
      LAYER pwell ;
        RECT 5.665 1803.275 5.835 1803.445 ;
        RECT 2913.785 1803.275 2913.955 1803.445 ;
      LAYER nwell ;
        RECT 5.330 1799.225 7.090 1802.055 ;
        RECT 2912.530 1799.225 2914.290 1802.055 ;
      LAYER pwell ;
        RECT 5.665 1797.835 5.835 1798.005 ;
        RECT 2913.785 1797.835 2913.955 1798.005 ;
      LAYER nwell ;
        RECT 5.330 1793.785 7.090 1796.615 ;
        RECT 2912.530 1793.785 2914.290 1796.615 ;
      LAYER pwell ;
        RECT 5.665 1792.395 5.835 1792.565 ;
        RECT 2913.785 1792.395 2913.955 1792.565 ;
      LAYER nwell ;
        RECT 5.330 1788.345 7.090 1791.175 ;
        RECT 2912.530 1788.345 2914.290 1791.175 ;
      LAYER pwell ;
        RECT 5.665 1786.955 5.835 1787.125 ;
        RECT 2913.785 1786.955 2913.955 1787.125 ;
      LAYER nwell ;
        RECT 5.330 1782.905 7.090 1785.735 ;
        RECT 2912.530 1782.905 2914.290 1785.735 ;
      LAYER pwell ;
        RECT 5.665 1781.515 5.835 1781.685 ;
        RECT 2913.785 1781.515 2913.955 1781.685 ;
      LAYER nwell ;
        RECT 5.330 1777.465 7.090 1780.295 ;
        RECT 8.550 1777.465 10.310 1779.070 ;
        RECT 2912.530 1777.465 2914.290 1780.295 ;
      LAYER pwell ;
        RECT 5.665 1776.075 5.835 1776.245 ;
        RECT 8.885 1776.075 9.055 1776.245 ;
        RECT 2913.785 1776.075 2913.955 1776.245 ;
      LAYER nwell ;
        RECT 5.330 1772.025 7.090 1774.855 ;
        RECT 2912.530 1772.025 2914.290 1774.855 ;
      LAYER pwell ;
        RECT 5.665 1770.635 5.835 1770.805 ;
        RECT 2913.785 1770.635 2913.955 1770.805 ;
      LAYER nwell ;
        RECT 5.330 1766.585 7.090 1769.415 ;
        RECT 2912.530 1766.585 2914.290 1769.415 ;
      LAYER pwell ;
        RECT 5.665 1765.195 5.835 1765.365 ;
        RECT 2913.785 1765.195 2913.955 1765.365 ;
      LAYER nwell ;
        RECT 5.330 1761.145 7.090 1763.975 ;
        RECT 2912.530 1761.145 2914.290 1763.975 ;
      LAYER pwell ;
        RECT 5.665 1759.755 5.835 1759.925 ;
        RECT 2913.785 1759.755 2913.955 1759.925 ;
      LAYER nwell ;
        RECT 5.330 1755.705 7.090 1758.535 ;
        RECT 2912.530 1755.705 2914.290 1758.535 ;
      LAYER pwell ;
        RECT 5.665 1754.315 5.835 1754.485 ;
        RECT 2913.785 1754.315 2913.955 1754.485 ;
      LAYER nwell ;
        RECT 5.330 1750.265 7.090 1753.095 ;
        RECT 2912.530 1750.265 2914.290 1753.095 ;
      LAYER pwell ;
        RECT 5.665 1748.875 5.835 1749.045 ;
        RECT 2913.785 1748.875 2913.955 1749.045 ;
      LAYER nwell ;
        RECT 5.330 1744.825 7.090 1747.655 ;
        RECT 2912.530 1744.825 2914.290 1747.655 ;
      LAYER pwell ;
        RECT 5.665 1743.435 5.835 1743.605 ;
        RECT 2913.785 1743.435 2913.955 1743.605 ;
      LAYER nwell ;
        RECT 5.330 1739.385 7.090 1742.215 ;
        RECT 2912.530 1739.385 2914.290 1742.215 ;
      LAYER pwell ;
        RECT 5.665 1737.995 5.835 1738.165 ;
        RECT 2913.785 1737.995 2913.955 1738.165 ;
      LAYER nwell ;
        RECT 5.330 1733.945 7.090 1736.775 ;
        RECT 2912.530 1733.945 2914.290 1736.775 ;
      LAYER pwell ;
        RECT 5.665 1732.555 5.835 1732.725 ;
        RECT 2913.785 1732.555 2913.955 1732.725 ;
      LAYER nwell ;
        RECT 5.330 1728.505 7.090 1731.335 ;
        RECT 2912.530 1728.505 2914.290 1731.335 ;
      LAYER pwell ;
        RECT 5.665 1727.115 5.835 1727.285 ;
        RECT 2913.785 1727.115 2913.955 1727.285 ;
      LAYER nwell ;
        RECT 5.330 1723.065 7.090 1725.895 ;
        RECT 2912.530 1723.065 2914.290 1725.895 ;
      LAYER pwell ;
        RECT 5.665 1721.675 5.835 1721.845 ;
        RECT 2913.785 1721.675 2913.955 1721.845 ;
      LAYER nwell ;
        RECT 5.330 1717.625 7.090 1720.455 ;
        RECT 2912.530 1717.625 2914.290 1720.455 ;
      LAYER pwell ;
        RECT 5.665 1716.235 5.835 1716.405 ;
        RECT 2913.785 1716.235 2913.955 1716.405 ;
      LAYER nwell ;
        RECT 5.330 1712.185 7.090 1715.015 ;
        RECT 2912.530 1712.185 2914.290 1715.015 ;
      LAYER pwell ;
        RECT 5.665 1710.795 5.835 1710.965 ;
        RECT 2913.785 1710.795 2913.955 1710.965 ;
      LAYER nwell ;
        RECT 5.330 1706.745 7.090 1709.575 ;
        RECT 8.550 1706.745 10.310 1708.350 ;
        RECT 2912.530 1706.745 2914.290 1709.575 ;
      LAYER pwell ;
        RECT 5.665 1705.355 5.835 1705.525 ;
        RECT 8.885 1705.355 9.055 1705.525 ;
        RECT 2913.785 1705.355 2913.955 1705.525 ;
      LAYER nwell ;
        RECT 5.330 1701.305 7.090 1704.135 ;
        RECT 2912.530 1701.305 2914.290 1704.135 ;
      LAYER pwell ;
        RECT 5.665 1699.915 5.835 1700.085 ;
        RECT 2913.785 1699.915 2913.955 1700.085 ;
      LAYER nwell ;
        RECT 5.330 1695.865 7.090 1698.695 ;
        RECT 2912.530 1695.865 2914.290 1698.695 ;
      LAYER pwell ;
        RECT 5.665 1694.475 5.835 1694.645 ;
        RECT 2913.785 1694.475 2913.955 1694.645 ;
      LAYER nwell ;
        RECT 5.330 1690.425 7.090 1693.255 ;
        RECT 2912.530 1690.425 2914.290 1693.255 ;
      LAYER pwell ;
        RECT 5.665 1689.035 5.835 1689.205 ;
        RECT 2913.785 1689.035 2913.955 1689.205 ;
      LAYER nwell ;
        RECT 5.330 1684.985 7.090 1687.815 ;
        RECT 2912.530 1684.985 2914.290 1687.815 ;
      LAYER pwell ;
        RECT 5.665 1683.595 5.835 1683.765 ;
        RECT 2913.785 1683.595 2913.955 1683.765 ;
      LAYER nwell ;
        RECT 5.330 1679.545 7.090 1682.375 ;
        RECT 2912.530 1679.545 2914.290 1682.375 ;
      LAYER pwell ;
        RECT 5.665 1678.155 5.835 1678.325 ;
        RECT 2913.785 1678.155 2913.955 1678.325 ;
      LAYER nwell ;
        RECT 5.330 1674.105 7.090 1676.935 ;
        RECT 2912.530 1674.105 2914.290 1676.935 ;
      LAYER pwell ;
        RECT 5.665 1672.715 5.835 1672.885 ;
        RECT 2909.185 1672.715 2909.355 1672.885 ;
        RECT 2913.785 1672.715 2913.955 1672.885 ;
      LAYER nwell ;
        RECT 5.330 1668.665 7.090 1671.495 ;
        RECT 2908.850 1669.890 2910.610 1671.495 ;
        RECT 2912.530 1668.665 2914.290 1671.495 ;
      LAYER pwell ;
        RECT 5.665 1667.275 5.835 1667.445 ;
        RECT 2913.785 1667.275 2913.955 1667.445 ;
      LAYER nwell ;
        RECT 5.330 1663.225 7.090 1666.055 ;
        RECT 2912.530 1663.225 2914.290 1666.055 ;
      LAYER pwell ;
        RECT 5.665 1661.835 5.835 1662.005 ;
        RECT 2913.785 1661.835 2913.955 1662.005 ;
      LAYER nwell ;
        RECT 5.330 1657.785 7.090 1660.615 ;
        RECT 2912.530 1657.785 2914.290 1660.615 ;
      LAYER pwell ;
        RECT 5.665 1656.395 5.835 1656.565 ;
        RECT 2913.785 1656.395 2913.955 1656.565 ;
      LAYER nwell ;
        RECT 5.330 1652.345 7.090 1655.175 ;
        RECT 2912.530 1652.345 2914.290 1655.175 ;
      LAYER pwell ;
        RECT 5.665 1650.955 5.835 1651.125 ;
        RECT 2913.785 1650.955 2913.955 1651.125 ;
      LAYER nwell ;
        RECT 5.330 1646.905 7.090 1649.735 ;
        RECT 2912.530 1646.905 2914.290 1649.735 ;
      LAYER pwell ;
        RECT 5.665 1645.515 5.835 1645.685 ;
        RECT 2913.785 1645.515 2913.955 1645.685 ;
      LAYER nwell ;
        RECT 5.330 1641.465 7.090 1644.295 ;
        RECT 2912.530 1641.465 2914.290 1644.295 ;
      LAYER pwell ;
        RECT 5.665 1640.075 5.835 1640.245 ;
        RECT 2913.785 1640.075 2913.955 1640.245 ;
      LAYER nwell ;
        RECT 5.330 1636.025 7.090 1638.855 ;
        RECT 2912.530 1636.025 2914.290 1638.855 ;
      LAYER pwell ;
        RECT 5.665 1634.635 5.835 1634.805 ;
        RECT 2913.785 1634.635 2913.955 1634.805 ;
      LAYER nwell ;
        RECT 5.330 1630.585 7.090 1633.415 ;
        RECT 2912.530 1630.585 2914.290 1633.415 ;
      LAYER pwell ;
        RECT 5.665 1629.195 5.835 1629.365 ;
        RECT 2913.785 1629.195 2913.955 1629.365 ;
      LAYER nwell ;
        RECT 5.330 1625.145 7.090 1627.975 ;
        RECT 2912.530 1625.145 2914.290 1627.975 ;
      LAYER pwell ;
        RECT 5.665 1623.755 5.835 1623.925 ;
        RECT 2913.785 1623.755 2913.955 1623.925 ;
      LAYER nwell ;
        RECT 5.330 1619.705 7.090 1622.535 ;
        RECT 2912.530 1619.705 2914.290 1622.535 ;
      LAYER pwell ;
        RECT 5.665 1618.315 5.835 1618.485 ;
        RECT 2913.785 1618.315 2913.955 1618.485 ;
      LAYER nwell ;
        RECT 5.330 1614.265 7.090 1617.095 ;
        RECT 2912.530 1614.265 2914.290 1617.095 ;
      LAYER pwell ;
        RECT 5.665 1612.875 5.835 1613.045 ;
        RECT 2913.785 1612.875 2913.955 1613.045 ;
      LAYER nwell ;
        RECT 5.330 1608.825 7.090 1611.655 ;
        RECT 2912.530 1608.825 2914.290 1611.655 ;
      LAYER pwell ;
        RECT 5.665 1607.435 5.835 1607.605 ;
        RECT 2913.785 1607.435 2913.955 1607.605 ;
      LAYER nwell ;
        RECT 5.330 1603.385 7.090 1606.215 ;
        RECT 2912.530 1603.385 2914.290 1606.215 ;
      LAYER pwell ;
        RECT 5.665 1601.995 5.835 1602.165 ;
        RECT 2913.785 1601.995 2913.955 1602.165 ;
      LAYER nwell ;
        RECT 5.330 1597.945 7.090 1600.775 ;
        RECT 2912.530 1597.945 2914.290 1600.775 ;
      LAYER pwell ;
        RECT 5.665 1596.555 5.835 1596.725 ;
        RECT 2913.785 1596.555 2913.955 1596.725 ;
      LAYER nwell ;
        RECT 5.330 1592.505 7.090 1595.335 ;
        RECT 2912.530 1592.505 2914.290 1595.335 ;
      LAYER pwell ;
        RECT 5.665 1591.115 5.835 1591.285 ;
        RECT 2913.785 1591.115 2913.955 1591.285 ;
      LAYER nwell ;
        RECT 5.330 1587.065 7.090 1589.895 ;
        RECT 2912.530 1587.065 2914.290 1589.895 ;
      LAYER pwell ;
        RECT 5.665 1585.675 5.835 1585.845 ;
        RECT 2913.785 1585.675 2913.955 1585.845 ;
      LAYER nwell ;
        RECT 5.330 1581.625 7.090 1584.455 ;
        RECT 8.550 1581.625 10.310 1583.230 ;
        RECT 2912.530 1581.625 2914.290 1584.455 ;
      LAYER pwell ;
        RECT 5.665 1580.235 5.835 1580.405 ;
        RECT 8.885 1580.235 9.055 1580.405 ;
        RECT 2913.785 1580.235 2913.955 1580.405 ;
      LAYER nwell ;
        RECT 5.330 1576.185 7.090 1579.015 ;
        RECT 2912.530 1576.185 2914.290 1579.015 ;
      LAYER pwell ;
        RECT 5.665 1574.795 5.835 1574.965 ;
        RECT 2913.785 1574.795 2913.955 1574.965 ;
      LAYER nwell ;
        RECT 5.330 1570.745 7.090 1573.575 ;
        RECT 2912.530 1570.745 2914.290 1573.575 ;
      LAYER pwell ;
        RECT 5.665 1569.355 5.835 1569.525 ;
        RECT 2913.785 1569.355 2913.955 1569.525 ;
      LAYER nwell ;
        RECT 5.330 1565.305 7.090 1568.135 ;
        RECT 2912.530 1565.305 2914.290 1568.135 ;
      LAYER pwell ;
        RECT 5.665 1563.915 5.835 1564.085 ;
        RECT 2913.785 1563.915 2913.955 1564.085 ;
      LAYER nwell ;
        RECT 5.330 1559.865 7.090 1562.695 ;
        RECT 2912.530 1559.865 2914.290 1562.695 ;
      LAYER pwell ;
        RECT 5.665 1558.475 5.835 1558.645 ;
        RECT 2913.785 1558.475 2913.955 1558.645 ;
      LAYER nwell ;
        RECT 5.330 1554.425 7.090 1557.255 ;
        RECT 2912.530 1554.425 2914.290 1557.255 ;
      LAYER pwell ;
        RECT 5.665 1553.035 5.835 1553.205 ;
        RECT 2913.785 1553.035 2913.955 1553.205 ;
      LAYER nwell ;
        RECT 5.330 1548.985 7.090 1551.815 ;
        RECT 2912.530 1548.985 2914.290 1551.815 ;
      LAYER pwell ;
        RECT 5.665 1547.595 5.835 1547.765 ;
        RECT 2913.785 1547.595 2913.955 1547.765 ;
      LAYER nwell ;
        RECT 5.330 1543.545 7.090 1546.375 ;
        RECT 2912.530 1543.545 2914.290 1546.375 ;
      LAYER pwell ;
        RECT 5.665 1542.155 5.835 1542.325 ;
        RECT 2913.785 1542.155 2913.955 1542.325 ;
      LAYER nwell ;
        RECT 5.330 1538.105 7.090 1540.935 ;
        RECT 2912.530 1538.105 2914.290 1540.935 ;
      LAYER pwell ;
        RECT 5.665 1536.715 5.835 1536.885 ;
        RECT 2913.785 1536.715 2913.955 1536.885 ;
      LAYER nwell ;
        RECT 5.330 1532.665 7.090 1535.495 ;
        RECT 2912.530 1532.665 2914.290 1535.495 ;
      LAYER pwell ;
        RECT 5.665 1531.275 5.835 1531.445 ;
        RECT 2913.785 1531.275 2913.955 1531.445 ;
      LAYER nwell ;
        RECT 5.330 1527.225 7.090 1530.055 ;
        RECT 2908.850 1527.225 2910.610 1528.830 ;
        RECT 2912.530 1527.225 2914.290 1530.055 ;
      LAYER pwell ;
        RECT 5.665 1525.835 5.835 1526.005 ;
        RECT 2909.185 1525.835 2909.355 1526.005 ;
        RECT 2913.785 1525.835 2913.955 1526.005 ;
      LAYER nwell ;
        RECT 5.330 1521.785 7.090 1524.615 ;
        RECT 2912.530 1521.785 2914.290 1524.615 ;
      LAYER pwell ;
        RECT 5.665 1520.395 5.835 1520.565 ;
        RECT 2913.785 1520.395 2913.955 1520.565 ;
      LAYER nwell ;
        RECT 5.330 1516.345 7.090 1519.175 ;
        RECT 2908.850 1516.345 2910.610 1517.950 ;
        RECT 2912.530 1516.345 2914.290 1519.175 ;
      LAYER pwell ;
        RECT 5.665 1514.955 5.835 1515.125 ;
        RECT 2909.185 1514.955 2909.355 1515.125 ;
        RECT 2913.785 1514.955 2913.955 1515.125 ;
      LAYER nwell ;
        RECT 5.330 1510.905 7.090 1513.735 ;
        RECT 2912.530 1510.905 2914.290 1513.735 ;
      LAYER pwell ;
        RECT 5.665 1509.515 5.835 1509.685 ;
        RECT 2913.785 1509.515 2913.955 1509.685 ;
      LAYER nwell ;
        RECT 5.330 1505.465 7.090 1508.295 ;
        RECT 2912.530 1505.465 2914.290 1508.295 ;
      LAYER pwell ;
        RECT 5.665 1504.075 5.835 1504.245 ;
        RECT 2913.785 1504.075 2913.955 1504.245 ;
      LAYER nwell ;
        RECT 5.330 1500.025 7.090 1502.855 ;
        RECT 2912.530 1500.025 2914.290 1502.855 ;
      LAYER pwell ;
        RECT 5.665 1498.635 5.835 1498.805 ;
        RECT 2913.785 1498.635 2913.955 1498.805 ;
      LAYER nwell ;
        RECT 5.330 1494.585 7.090 1497.415 ;
        RECT 2912.530 1494.585 2914.290 1497.415 ;
      LAYER pwell ;
        RECT 5.665 1493.195 5.835 1493.365 ;
        RECT 2913.785 1493.195 2913.955 1493.365 ;
      LAYER nwell ;
        RECT 5.330 1489.145 7.090 1491.975 ;
        RECT 2912.530 1489.145 2914.290 1491.975 ;
      LAYER pwell ;
        RECT 5.665 1487.755 5.835 1487.925 ;
        RECT 2913.785 1487.755 2913.955 1487.925 ;
      LAYER nwell ;
        RECT 5.330 1483.705 7.090 1486.535 ;
        RECT 2912.530 1483.705 2914.290 1486.535 ;
      LAYER pwell ;
        RECT 5.665 1482.315 5.835 1482.485 ;
        RECT 2913.785 1482.315 2913.955 1482.485 ;
      LAYER nwell ;
        RECT 5.330 1478.265 7.090 1481.095 ;
        RECT 2912.530 1478.265 2914.290 1481.095 ;
      LAYER pwell ;
        RECT 5.665 1476.875 5.835 1477.045 ;
        RECT 2913.785 1476.875 2913.955 1477.045 ;
      LAYER nwell ;
        RECT 5.330 1472.825 7.090 1475.655 ;
        RECT 2908.850 1472.825 2910.610 1474.430 ;
        RECT 2912.530 1472.825 2914.290 1475.655 ;
      LAYER pwell ;
        RECT 5.665 1471.435 5.835 1471.605 ;
        RECT 2909.185 1471.435 2909.355 1471.605 ;
        RECT 2913.785 1471.435 2913.955 1471.605 ;
      LAYER nwell ;
        RECT 5.330 1467.385 7.090 1470.215 ;
        RECT 2912.530 1467.385 2914.290 1470.215 ;
      LAYER pwell ;
        RECT 5.665 1465.995 5.835 1466.165 ;
        RECT 2913.785 1465.995 2913.955 1466.165 ;
      LAYER nwell ;
        RECT 5.330 1461.945 7.090 1464.775 ;
        RECT 2912.530 1461.945 2914.290 1464.775 ;
      LAYER pwell ;
        RECT 5.665 1460.555 5.835 1460.725 ;
        RECT 2913.785 1460.555 2913.955 1460.725 ;
      LAYER nwell ;
        RECT 5.330 1456.505 7.090 1459.335 ;
        RECT 2912.530 1456.505 2914.290 1459.335 ;
      LAYER pwell ;
        RECT 5.665 1455.115 5.835 1455.285 ;
        RECT 2913.785 1455.115 2913.955 1455.285 ;
      LAYER nwell ;
        RECT 5.330 1451.065 7.090 1453.895 ;
        RECT 2912.530 1451.065 2914.290 1453.895 ;
      LAYER pwell ;
        RECT 5.665 1449.675 5.835 1449.845 ;
        RECT 2913.785 1449.675 2913.955 1449.845 ;
      LAYER nwell ;
        RECT 5.330 1445.625 7.090 1448.455 ;
        RECT 2912.530 1445.625 2914.290 1448.455 ;
      LAYER pwell ;
        RECT 5.665 1444.235 5.835 1444.405 ;
        RECT 2913.785 1444.235 2913.955 1444.405 ;
      LAYER nwell ;
        RECT 5.330 1440.185 7.090 1443.015 ;
        RECT 2912.530 1440.185 2914.290 1443.015 ;
      LAYER pwell ;
        RECT 5.665 1438.795 5.835 1438.965 ;
        RECT 2913.785 1438.795 2913.955 1438.965 ;
      LAYER nwell ;
        RECT 5.330 1434.745 7.090 1437.575 ;
        RECT 2912.530 1434.745 2914.290 1437.575 ;
      LAYER pwell ;
        RECT 5.665 1433.355 5.835 1433.525 ;
        RECT 2913.785 1433.355 2913.955 1433.525 ;
      LAYER nwell ;
        RECT 5.330 1429.305 7.090 1432.135 ;
        RECT 2912.530 1429.305 2914.290 1432.135 ;
      LAYER pwell ;
        RECT 5.665 1427.915 5.835 1428.085 ;
        RECT 2913.785 1427.915 2913.955 1428.085 ;
      LAYER nwell ;
        RECT 5.330 1423.865 7.090 1426.695 ;
        RECT 2912.530 1423.865 2914.290 1426.695 ;
      LAYER pwell ;
        RECT 5.665 1422.475 5.835 1422.645 ;
        RECT 2913.785 1422.475 2913.955 1422.645 ;
      LAYER nwell ;
        RECT 5.330 1418.425 7.090 1421.255 ;
        RECT 2912.530 1418.425 2914.290 1421.255 ;
      LAYER pwell ;
        RECT 5.665 1417.035 5.835 1417.205 ;
        RECT 2913.785 1417.035 2913.955 1417.205 ;
      LAYER nwell ;
        RECT 5.330 1412.985 7.090 1415.815 ;
        RECT 2912.530 1412.985 2914.290 1415.815 ;
      LAYER pwell ;
        RECT 5.665 1411.595 5.835 1411.765 ;
        RECT 2913.785 1411.595 2913.955 1411.765 ;
      LAYER nwell ;
        RECT 5.330 1407.545 7.090 1410.375 ;
        RECT 2912.530 1407.545 2914.290 1410.375 ;
      LAYER pwell ;
        RECT 5.665 1406.155 5.835 1406.325 ;
        RECT 2913.785 1406.155 2913.955 1406.325 ;
      LAYER nwell ;
        RECT 5.330 1402.105 7.090 1404.935 ;
        RECT 2912.530 1402.105 2914.290 1404.935 ;
      LAYER pwell ;
        RECT 5.665 1400.715 5.835 1400.885 ;
        RECT 2913.785 1400.715 2913.955 1400.885 ;
      LAYER nwell ;
        RECT 5.330 1396.665 7.090 1399.495 ;
        RECT 2912.530 1396.665 2914.290 1399.495 ;
      LAYER pwell ;
        RECT 5.665 1395.275 5.835 1395.445 ;
        RECT 2913.785 1395.275 2913.955 1395.445 ;
      LAYER nwell ;
        RECT 5.330 1391.225 7.090 1394.055 ;
        RECT 2912.530 1391.225 2914.290 1394.055 ;
      LAYER pwell ;
        RECT 5.665 1389.835 5.835 1390.005 ;
        RECT 2913.785 1389.835 2913.955 1390.005 ;
      LAYER nwell ;
        RECT 5.330 1385.785 7.090 1388.615 ;
        RECT 2912.530 1385.785 2914.290 1388.615 ;
      LAYER pwell ;
        RECT 5.665 1384.395 5.835 1384.565 ;
        RECT 2913.785 1384.395 2913.955 1384.565 ;
      LAYER nwell ;
        RECT 5.330 1380.345 7.090 1383.175 ;
        RECT 2912.530 1380.345 2914.290 1383.175 ;
      LAYER pwell ;
        RECT 5.665 1378.955 5.835 1379.125 ;
        RECT 2913.785 1378.955 2913.955 1379.125 ;
      LAYER nwell ;
        RECT 5.330 1374.905 7.090 1377.735 ;
        RECT 2912.530 1374.905 2914.290 1377.735 ;
      LAYER pwell ;
        RECT 5.665 1373.515 5.835 1373.685 ;
        RECT 2913.785 1373.515 2913.955 1373.685 ;
      LAYER nwell ;
        RECT 5.330 1369.465 7.090 1372.295 ;
        RECT 2912.530 1369.465 2914.290 1372.295 ;
      LAYER pwell ;
        RECT 5.665 1368.075 5.835 1368.245 ;
        RECT 2913.785 1368.075 2913.955 1368.245 ;
      LAYER nwell ;
        RECT 5.330 1364.025 7.090 1366.855 ;
        RECT 2912.530 1364.025 2914.290 1366.855 ;
      LAYER pwell ;
        RECT 5.665 1362.635 5.835 1362.805 ;
        RECT 2913.785 1362.635 2913.955 1362.805 ;
      LAYER nwell ;
        RECT 5.330 1358.585 7.090 1361.415 ;
        RECT 2912.530 1358.585 2914.290 1361.415 ;
      LAYER pwell ;
        RECT 5.665 1357.195 5.835 1357.365 ;
        RECT 2913.785 1357.195 2913.955 1357.365 ;
      LAYER nwell ;
        RECT 5.330 1353.145 7.090 1355.975 ;
        RECT 2912.530 1353.145 2914.290 1355.975 ;
      LAYER pwell ;
        RECT 5.665 1351.755 5.835 1351.925 ;
        RECT 2913.785 1351.755 2913.955 1351.925 ;
      LAYER nwell ;
        RECT 5.330 1347.705 7.090 1350.535 ;
        RECT 2912.530 1347.705 2914.290 1350.535 ;
      LAYER pwell ;
        RECT 5.665 1346.315 5.835 1346.485 ;
        RECT 2913.785 1346.315 2913.955 1346.485 ;
      LAYER nwell ;
        RECT 5.330 1342.265 7.090 1345.095 ;
        RECT 2912.530 1342.265 2914.290 1345.095 ;
      LAYER pwell ;
        RECT 5.665 1340.875 5.835 1341.045 ;
        RECT 2913.785 1340.875 2913.955 1341.045 ;
      LAYER nwell ;
        RECT 5.330 1336.825 7.090 1339.655 ;
        RECT 2912.530 1336.825 2914.290 1339.655 ;
      LAYER pwell ;
        RECT 5.665 1335.435 5.835 1335.605 ;
        RECT 2913.785 1335.435 2913.955 1335.605 ;
      LAYER nwell ;
        RECT 5.330 1331.385 7.090 1334.215 ;
        RECT 2912.530 1331.385 2914.290 1334.215 ;
      LAYER pwell ;
        RECT 5.665 1329.995 5.835 1330.165 ;
        RECT 8.885 1329.995 9.055 1330.165 ;
        RECT 2913.785 1329.995 2913.955 1330.165 ;
      LAYER nwell ;
        RECT 5.330 1325.945 7.090 1328.775 ;
        RECT 8.550 1327.170 10.310 1328.775 ;
        RECT 2912.530 1325.945 2914.290 1328.775 ;
      LAYER pwell ;
        RECT 5.665 1324.555 5.835 1324.725 ;
        RECT 2913.785 1324.555 2913.955 1324.725 ;
      LAYER nwell ;
        RECT 5.330 1320.505 7.090 1323.335 ;
        RECT 2912.530 1320.505 2914.290 1323.335 ;
      LAYER pwell ;
        RECT 5.665 1319.115 5.835 1319.285 ;
        RECT 2913.785 1319.115 2913.955 1319.285 ;
      LAYER nwell ;
        RECT 5.330 1315.065 7.090 1317.895 ;
        RECT 2912.530 1315.065 2914.290 1317.895 ;
      LAYER pwell ;
        RECT 5.665 1313.675 5.835 1313.845 ;
        RECT 2913.785 1313.675 2913.955 1313.845 ;
      LAYER nwell ;
        RECT 5.330 1309.625 7.090 1312.455 ;
        RECT 2912.530 1309.625 2914.290 1312.455 ;
      LAYER pwell ;
        RECT 5.665 1308.235 5.835 1308.405 ;
        RECT 2913.785 1308.235 2913.955 1308.405 ;
      LAYER nwell ;
        RECT 5.330 1304.185 7.090 1307.015 ;
        RECT 2912.530 1304.185 2914.290 1307.015 ;
      LAYER pwell ;
        RECT 5.665 1302.795 5.835 1302.965 ;
        RECT 2909.185 1302.795 2909.355 1302.965 ;
        RECT 2913.785 1302.795 2913.955 1302.965 ;
      LAYER nwell ;
        RECT 5.330 1298.745 7.090 1301.575 ;
        RECT 2908.850 1299.970 2910.610 1301.575 ;
        RECT 2912.530 1298.745 2914.290 1301.575 ;
      LAYER pwell ;
        RECT 5.665 1297.355 5.835 1297.525 ;
        RECT 2913.785 1297.355 2913.955 1297.525 ;
      LAYER nwell ;
        RECT 5.330 1293.305 7.090 1296.135 ;
        RECT 2912.530 1293.305 2914.290 1296.135 ;
      LAYER pwell ;
        RECT 5.665 1291.915 5.835 1292.085 ;
        RECT 2913.785 1291.915 2913.955 1292.085 ;
      LAYER nwell ;
        RECT 5.330 1287.865 7.090 1290.695 ;
        RECT 2912.530 1287.865 2914.290 1290.695 ;
      LAYER pwell ;
        RECT 5.665 1286.475 5.835 1286.645 ;
        RECT 8.885 1286.475 9.055 1286.645 ;
        RECT 2913.785 1286.475 2913.955 1286.645 ;
      LAYER nwell ;
        RECT 5.330 1282.425 7.090 1285.255 ;
        RECT 8.550 1283.650 10.310 1285.255 ;
        RECT 2912.530 1282.425 2914.290 1285.255 ;
      LAYER pwell ;
        RECT 5.665 1281.035 5.835 1281.205 ;
        RECT 2913.785 1281.035 2913.955 1281.205 ;
      LAYER nwell ;
        RECT 5.330 1276.985 7.090 1279.815 ;
        RECT 2912.530 1276.985 2914.290 1279.815 ;
      LAYER pwell ;
        RECT 5.665 1275.595 5.835 1275.765 ;
        RECT 8.885 1275.595 9.055 1275.765 ;
        RECT 2913.785 1275.595 2913.955 1275.765 ;
      LAYER nwell ;
        RECT 5.330 1271.545 7.090 1274.375 ;
        RECT 8.550 1272.770 10.310 1274.375 ;
        RECT 2912.530 1271.545 2914.290 1274.375 ;
      LAYER pwell ;
        RECT 5.665 1270.155 5.835 1270.325 ;
        RECT 2913.785 1270.155 2913.955 1270.325 ;
      LAYER nwell ;
        RECT 5.330 1266.105 7.090 1268.935 ;
        RECT 2908.850 1266.105 2910.610 1267.710 ;
        RECT 2912.530 1266.105 2914.290 1268.935 ;
      LAYER pwell ;
        RECT 5.665 1264.715 5.835 1264.885 ;
        RECT 2909.185 1264.715 2909.355 1264.885 ;
        RECT 2913.785 1264.715 2913.955 1264.885 ;
      LAYER nwell ;
        RECT 5.330 1260.665 7.090 1263.495 ;
        RECT 2912.530 1260.665 2914.290 1263.495 ;
      LAYER pwell ;
        RECT 5.665 1259.275 5.835 1259.445 ;
        RECT 2913.785 1259.275 2913.955 1259.445 ;
      LAYER nwell ;
        RECT 5.330 1255.225 7.090 1258.055 ;
        RECT 2912.530 1255.225 2914.290 1258.055 ;
      LAYER pwell ;
        RECT 5.665 1253.835 5.835 1254.005 ;
        RECT 2913.785 1253.835 2913.955 1254.005 ;
      LAYER nwell ;
        RECT 5.330 1249.785 7.090 1252.615 ;
        RECT 2912.530 1249.785 2914.290 1252.615 ;
      LAYER pwell ;
        RECT 5.665 1248.395 5.835 1248.565 ;
        RECT 2913.785 1248.395 2913.955 1248.565 ;
      LAYER nwell ;
        RECT 5.330 1244.345 7.090 1247.175 ;
        RECT 2912.530 1244.345 2914.290 1247.175 ;
      LAYER pwell ;
        RECT 5.665 1242.955 5.835 1243.125 ;
        RECT 2913.785 1242.955 2913.955 1243.125 ;
      LAYER nwell ;
        RECT 5.330 1238.905 7.090 1241.735 ;
        RECT 2912.530 1238.905 2914.290 1241.735 ;
      LAYER pwell ;
        RECT 5.665 1237.515 5.835 1237.685 ;
        RECT 2913.785 1237.515 2913.955 1237.685 ;
      LAYER nwell ;
        RECT 5.330 1233.465 7.090 1236.295 ;
        RECT 2912.530 1233.465 2914.290 1236.295 ;
      LAYER pwell ;
        RECT 5.665 1232.075 5.835 1232.245 ;
        RECT 2913.785 1232.075 2913.955 1232.245 ;
      LAYER nwell ;
        RECT 5.330 1228.025 7.090 1230.855 ;
        RECT 2912.530 1228.025 2914.290 1230.855 ;
      LAYER pwell ;
        RECT 5.665 1226.635 5.835 1226.805 ;
        RECT 2913.785 1226.635 2913.955 1226.805 ;
      LAYER nwell ;
        RECT 5.330 1222.585 7.090 1225.415 ;
        RECT 2912.530 1222.585 2914.290 1225.415 ;
      LAYER pwell ;
        RECT 5.665 1221.195 5.835 1221.365 ;
        RECT 2913.785 1221.195 2913.955 1221.365 ;
      LAYER nwell ;
        RECT 5.330 1217.145 7.090 1219.975 ;
        RECT 8.550 1217.145 10.310 1218.750 ;
        RECT 2912.530 1217.145 2914.290 1219.975 ;
      LAYER pwell ;
        RECT 5.665 1215.755 5.835 1215.925 ;
        RECT 8.885 1215.755 9.055 1215.925 ;
        RECT 2913.785 1215.755 2913.955 1215.925 ;
      LAYER nwell ;
        RECT 5.330 1211.705 7.090 1214.535 ;
        RECT 2912.530 1211.705 2914.290 1214.535 ;
      LAYER pwell ;
        RECT 5.665 1210.315 5.835 1210.485 ;
        RECT 2913.785 1210.315 2913.955 1210.485 ;
      LAYER nwell ;
        RECT 5.330 1206.265 7.090 1209.095 ;
        RECT 2912.530 1206.265 2914.290 1209.095 ;
      LAYER pwell ;
        RECT 5.665 1204.875 5.835 1205.045 ;
        RECT 2913.785 1204.875 2913.955 1205.045 ;
      LAYER nwell ;
        RECT 5.330 1200.825 7.090 1203.655 ;
        RECT 2912.530 1200.825 2914.290 1203.655 ;
      LAYER pwell ;
        RECT 5.665 1199.435 5.835 1199.605 ;
        RECT 2913.785 1199.435 2913.955 1199.605 ;
      LAYER nwell ;
        RECT 5.330 1195.385 7.090 1198.215 ;
        RECT 2912.530 1195.385 2914.290 1198.215 ;
      LAYER pwell ;
        RECT 5.665 1193.995 5.835 1194.165 ;
        RECT 2913.785 1193.995 2913.955 1194.165 ;
      LAYER nwell ;
        RECT 5.330 1189.945 7.090 1192.775 ;
        RECT 2912.530 1189.945 2914.290 1192.775 ;
      LAYER pwell ;
        RECT 5.665 1188.555 5.835 1188.725 ;
        RECT 2913.785 1188.555 2913.955 1188.725 ;
      LAYER nwell ;
        RECT 5.330 1184.505 7.090 1187.335 ;
        RECT 2912.530 1184.505 2914.290 1187.335 ;
      LAYER pwell ;
        RECT 5.665 1183.115 5.835 1183.285 ;
        RECT 2913.785 1183.115 2913.955 1183.285 ;
      LAYER nwell ;
        RECT 5.330 1179.065 7.090 1181.895 ;
        RECT 2912.530 1179.065 2914.290 1181.895 ;
      LAYER pwell ;
        RECT 5.665 1177.675 5.835 1177.845 ;
        RECT 2913.785 1177.675 2913.955 1177.845 ;
      LAYER nwell ;
        RECT 5.330 1173.625 7.090 1176.455 ;
        RECT 2912.530 1173.625 2914.290 1176.455 ;
      LAYER pwell ;
        RECT 5.665 1172.235 5.835 1172.405 ;
        RECT 2913.785 1172.235 2913.955 1172.405 ;
      LAYER nwell ;
        RECT 5.330 1168.185 7.090 1171.015 ;
        RECT 2912.530 1168.185 2914.290 1171.015 ;
      LAYER pwell ;
        RECT 5.665 1166.795 5.835 1166.965 ;
        RECT 2913.785 1166.795 2913.955 1166.965 ;
      LAYER nwell ;
        RECT 5.330 1162.745 7.090 1165.575 ;
        RECT 2912.530 1162.745 2914.290 1165.575 ;
      LAYER pwell ;
        RECT 5.665 1161.355 5.835 1161.525 ;
        RECT 2913.785 1161.355 2913.955 1161.525 ;
      LAYER nwell ;
        RECT 5.330 1157.305 7.090 1160.135 ;
        RECT 2912.530 1157.305 2914.290 1160.135 ;
      LAYER pwell ;
        RECT 5.665 1155.915 5.835 1156.085 ;
        RECT 2913.785 1155.915 2913.955 1156.085 ;
      LAYER nwell ;
        RECT 5.330 1151.865 7.090 1154.695 ;
        RECT 2912.530 1151.865 2914.290 1154.695 ;
      LAYER pwell ;
        RECT 5.665 1150.475 5.835 1150.645 ;
        RECT 2913.785 1150.475 2913.955 1150.645 ;
      LAYER nwell ;
        RECT 5.330 1146.425 7.090 1149.255 ;
        RECT 2912.530 1146.425 2914.290 1149.255 ;
      LAYER pwell ;
        RECT 5.665 1145.035 5.835 1145.205 ;
        RECT 2913.785 1145.035 2913.955 1145.205 ;
      LAYER nwell ;
        RECT 5.330 1140.985 7.090 1143.815 ;
        RECT 2912.530 1140.985 2914.290 1143.815 ;
      LAYER pwell ;
        RECT 5.665 1139.595 5.835 1139.765 ;
        RECT 2913.785 1139.595 2913.955 1139.765 ;
      LAYER nwell ;
        RECT 5.330 1135.545 7.090 1138.375 ;
        RECT 2912.530 1135.545 2914.290 1138.375 ;
      LAYER pwell ;
        RECT 5.665 1134.155 5.835 1134.325 ;
        RECT 2913.785 1134.155 2913.955 1134.325 ;
      LAYER nwell ;
        RECT 5.330 1130.105 7.090 1132.935 ;
        RECT 2912.530 1130.105 2914.290 1132.935 ;
      LAYER pwell ;
        RECT 5.665 1128.715 5.835 1128.885 ;
        RECT 2913.785 1128.715 2913.955 1128.885 ;
      LAYER nwell ;
        RECT 5.330 1124.665 7.090 1127.495 ;
        RECT 2912.530 1124.665 2914.290 1127.495 ;
      LAYER pwell ;
        RECT 5.665 1123.275 5.835 1123.445 ;
        RECT 2913.785 1123.275 2913.955 1123.445 ;
      LAYER nwell ;
        RECT 5.330 1119.225 7.090 1122.055 ;
        RECT 2912.530 1119.225 2914.290 1122.055 ;
      LAYER pwell ;
        RECT 5.665 1117.835 5.835 1118.005 ;
        RECT 2913.785 1117.835 2913.955 1118.005 ;
      LAYER nwell ;
        RECT 5.330 1113.785 7.090 1116.615 ;
        RECT 2912.530 1113.785 2914.290 1116.615 ;
      LAYER pwell ;
        RECT 5.665 1112.395 5.835 1112.565 ;
        RECT 8.885 1112.395 9.055 1112.565 ;
        RECT 2913.785 1112.395 2913.955 1112.565 ;
      LAYER nwell ;
        RECT 5.330 1108.345 7.090 1111.175 ;
        RECT 8.550 1109.570 10.310 1111.175 ;
        RECT 2912.530 1108.345 2914.290 1111.175 ;
      LAYER pwell ;
        RECT 5.665 1106.955 5.835 1107.125 ;
        RECT 2913.785 1106.955 2913.955 1107.125 ;
      LAYER nwell ;
        RECT 5.330 1102.905 7.090 1105.735 ;
        RECT 2912.530 1102.905 2914.290 1105.735 ;
      LAYER pwell ;
        RECT 5.665 1101.515 5.835 1101.685 ;
        RECT 2913.785 1101.515 2913.955 1101.685 ;
      LAYER nwell ;
        RECT 5.330 1097.465 7.090 1100.295 ;
        RECT 2912.530 1097.465 2914.290 1100.295 ;
      LAYER pwell ;
        RECT 5.665 1096.075 5.835 1096.245 ;
        RECT 2913.785 1096.075 2913.955 1096.245 ;
      LAYER nwell ;
        RECT 5.330 1092.025 7.090 1094.855 ;
        RECT 2912.530 1092.025 2914.290 1094.855 ;
      LAYER pwell ;
        RECT 5.665 1090.635 5.835 1090.805 ;
        RECT 2913.785 1090.635 2913.955 1090.805 ;
      LAYER nwell ;
        RECT 5.330 1086.585 7.090 1089.415 ;
        RECT 2912.530 1086.585 2914.290 1089.415 ;
      LAYER pwell ;
        RECT 5.665 1085.195 5.835 1085.365 ;
        RECT 2913.785 1085.195 2913.955 1085.365 ;
      LAYER nwell ;
        RECT 5.330 1081.145 7.090 1083.975 ;
        RECT 2912.530 1081.145 2914.290 1083.975 ;
      LAYER pwell ;
        RECT 5.665 1079.755 5.835 1079.925 ;
        RECT 2913.785 1079.755 2913.955 1079.925 ;
      LAYER nwell ;
        RECT 5.330 1075.705 7.090 1078.535 ;
        RECT 2912.530 1075.705 2914.290 1078.535 ;
      LAYER pwell ;
        RECT 5.665 1074.315 5.835 1074.485 ;
        RECT 2913.785 1074.315 2913.955 1074.485 ;
      LAYER nwell ;
        RECT 5.330 1070.265 7.090 1073.095 ;
        RECT 2912.530 1070.265 2914.290 1073.095 ;
      LAYER pwell ;
        RECT 5.665 1068.875 5.835 1069.045 ;
        RECT 2913.785 1068.875 2913.955 1069.045 ;
      LAYER nwell ;
        RECT 5.330 1064.825 7.090 1067.655 ;
        RECT 2912.530 1064.825 2914.290 1067.655 ;
      LAYER pwell ;
        RECT 5.665 1063.435 5.835 1063.605 ;
        RECT 2913.785 1063.435 2913.955 1063.605 ;
      LAYER nwell ;
        RECT 5.330 1059.385 7.090 1062.215 ;
        RECT 2912.530 1059.385 2914.290 1062.215 ;
      LAYER pwell ;
        RECT 5.665 1057.995 5.835 1058.165 ;
        RECT 2913.785 1057.995 2913.955 1058.165 ;
      LAYER nwell ;
        RECT 5.330 1053.945 7.090 1056.775 ;
        RECT 2912.530 1053.945 2914.290 1056.775 ;
      LAYER pwell ;
        RECT 5.665 1052.555 5.835 1052.725 ;
        RECT 2913.785 1052.555 2913.955 1052.725 ;
      LAYER nwell ;
        RECT 5.330 1048.505 7.090 1051.335 ;
        RECT 2912.530 1048.505 2914.290 1051.335 ;
      LAYER pwell ;
        RECT 5.665 1047.115 5.835 1047.285 ;
        RECT 2913.785 1047.115 2913.955 1047.285 ;
      LAYER nwell ;
        RECT 5.330 1043.065 7.090 1045.895 ;
        RECT 2912.530 1043.065 2914.290 1045.895 ;
      LAYER pwell ;
        RECT 5.665 1041.675 5.835 1041.845 ;
        RECT 2913.785 1041.675 2913.955 1041.845 ;
      LAYER nwell ;
        RECT 5.330 1037.625 7.090 1040.455 ;
        RECT 2912.530 1037.625 2914.290 1040.455 ;
      LAYER pwell ;
        RECT 5.665 1036.235 5.835 1036.405 ;
        RECT 8.885 1036.235 9.055 1036.405 ;
        RECT 2913.785 1036.235 2913.955 1036.405 ;
      LAYER nwell ;
        RECT 5.330 1032.185 7.090 1035.015 ;
        RECT 8.550 1033.410 10.310 1035.015 ;
        RECT 2912.530 1032.185 2914.290 1035.015 ;
      LAYER pwell ;
        RECT 5.665 1030.795 5.835 1030.965 ;
        RECT 2913.785 1030.795 2913.955 1030.965 ;
      LAYER nwell ;
        RECT 5.330 1026.745 7.090 1029.575 ;
        RECT 2912.530 1026.745 2914.290 1029.575 ;
      LAYER pwell ;
        RECT 5.665 1025.355 5.835 1025.525 ;
        RECT 2913.785 1025.355 2913.955 1025.525 ;
      LAYER nwell ;
        RECT 5.330 1021.305 7.090 1024.135 ;
        RECT 2912.530 1021.305 2914.290 1024.135 ;
      LAYER pwell ;
        RECT 5.665 1019.915 5.835 1020.085 ;
        RECT 2913.785 1019.915 2913.955 1020.085 ;
      LAYER nwell ;
        RECT 5.330 1015.865 7.090 1018.695 ;
        RECT 2912.530 1015.865 2914.290 1018.695 ;
      LAYER pwell ;
        RECT 5.665 1014.475 5.835 1014.645 ;
        RECT 2913.785 1014.475 2913.955 1014.645 ;
      LAYER nwell ;
        RECT 5.330 1010.425 7.090 1013.255 ;
        RECT 2912.530 1010.425 2914.290 1013.255 ;
      LAYER pwell ;
        RECT 5.665 1009.035 5.835 1009.205 ;
        RECT 2909.185 1009.035 2909.355 1009.205 ;
        RECT 2913.785 1009.035 2913.955 1009.205 ;
      LAYER nwell ;
        RECT 5.330 1004.985 7.090 1007.815 ;
        RECT 2912.530 1004.985 2914.290 1007.815 ;
      LAYER pwell ;
        RECT 5.665 1003.595 5.835 1003.765 ;
        RECT 2913.785 1003.595 2913.955 1003.765 ;
      LAYER nwell ;
        RECT 5.330 999.545 7.090 1002.375 ;
        RECT 2912.530 999.545 2914.290 1002.375 ;
      LAYER pwell ;
        RECT 5.665 998.155 5.835 998.325 ;
        RECT 2909.185 998.155 2909.355 998.325 ;
        RECT 2913.785 998.155 2913.955 998.325 ;
      LAYER nwell ;
        RECT 5.330 994.105 7.090 996.935 ;
        RECT 2912.530 994.105 2914.290 996.935 ;
      LAYER pwell ;
        RECT 5.665 992.715 5.835 992.885 ;
        RECT 2913.785 992.715 2913.955 992.885 ;
      LAYER nwell ;
        RECT 5.330 988.665 7.090 991.495 ;
        RECT 2912.530 988.665 2914.290 991.495 ;
      LAYER pwell ;
        RECT 5.665 987.275 5.835 987.445 ;
        RECT 2913.785 987.275 2913.955 987.445 ;
      LAYER nwell ;
        RECT 5.330 983.225 7.090 986.055 ;
        RECT 2912.530 983.225 2914.290 986.055 ;
      LAYER pwell ;
        RECT 5.665 981.835 5.835 982.005 ;
        RECT 2913.785 981.835 2913.955 982.005 ;
      LAYER nwell ;
        RECT 5.330 977.785 7.090 980.615 ;
        RECT 2912.530 977.785 2914.290 980.615 ;
      LAYER pwell ;
        RECT 5.665 976.395 5.835 976.565 ;
        RECT 2913.785 976.395 2913.955 976.565 ;
      LAYER nwell ;
        RECT 5.330 972.345 7.090 975.175 ;
        RECT 2912.530 972.345 2914.290 975.175 ;
      LAYER pwell ;
        RECT 5.665 970.955 5.835 971.125 ;
        RECT 2913.785 970.955 2913.955 971.125 ;
      LAYER nwell ;
        RECT 5.330 966.905 7.090 969.735 ;
        RECT 2912.530 966.905 2914.290 969.735 ;
      LAYER pwell ;
        RECT 5.665 965.515 5.835 965.685 ;
        RECT 2913.785 965.515 2913.955 965.685 ;
      LAYER nwell ;
        RECT 5.330 961.465 7.090 964.295 ;
        RECT 2912.530 961.465 2914.290 964.295 ;
      LAYER pwell ;
        RECT 5.665 960.075 5.835 960.245 ;
        RECT 2913.785 960.075 2913.955 960.245 ;
      LAYER nwell ;
        RECT 5.330 956.025 7.090 958.855 ;
        RECT 2912.530 956.025 2914.290 958.855 ;
      LAYER pwell ;
        RECT 5.665 954.635 5.835 954.805 ;
        RECT 2913.785 954.635 2913.955 954.805 ;
      LAYER nwell ;
        RECT 5.330 950.585 7.090 953.415 ;
        RECT 2912.530 950.585 2914.290 953.415 ;
      LAYER pwell ;
        RECT 5.665 949.195 5.835 949.365 ;
        RECT 2913.785 949.195 2913.955 949.365 ;
      LAYER nwell ;
        RECT 5.330 945.145 7.090 947.975 ;
        RECT 2912.530 945.145 2914.290 947.975 ;
      LAYER pwell ;
        RECT 5.665 943.755 5.835 943.925 ;
        RECT 2913.785 943.755 2913.955 943.925 ;
      LAYER nwell ;
        RECT 5.330 939.705 7.090 942.535 ;
        RECT 2912.530 939.705 2914.290 942.535 ;
      LAYER pwell ;
        RECT 5.665 938.315 5.835 938.485 ;
        RECT 2913.785 938.315 2913.955 938.485 ;
      LAYER nwell ;
        RECT 5.330 934.265 7.090 937.095 ;
        RECT 2912.530 934.265 2914.290 937.095 ;
      LAYER pwell ;
        RECT 5.665 932.875 5.835 933.045 ;
        RECT 2913.785 932.875 2913.955 933.045 ;
      LAYER nwell ;
        RECT 5.330 928.825 7.090 931.655 ;
        RECT 2912.530 928.825 2914.290 931.655 ;
      LAYER pwell ;
        RECT 5.665 927.435 5.835 927.605 ;
        RECT 2913.785 927.435 2913.955 927.605 ;
      LAYER nwell ;
        RECT 5.330 923.385 7.090 926.215 ;
        RECT 2912.530 923.385 2914.290 926.215 ;
      LAYER pwell ;
        RECT 5.665 921.995 5.835 922.165 ;
        RECT 2913.785 921.995 2913.955 922.165 ;
      LAYER nwell ;
        RECT 5.330 917.945 7.090 920.775 ;
        RECT 2912.530 917.945 2914.290 920.775 ;
      LAYER pwell ;
        RECT 5.665 916.555 5.835 916.725 ;
        RECT 2913.785 916.555 2913.955 916.725 ;
      LAYER nwell ;
        RECT 5.330 912.505 7.090 915.335 ;
        RECT 2912.530 912.505 2914.290 915.335 ;
      LAYER pwell ;
        RECT 5.665 911.115 5.835 911.285 ;
        RECT 2913.785 911.115 2913.955 911.285 ;
      LAYER nwell ;
        RECT 5.330 907.065 7.090 909.895 ;
        RECT 2912.530 907.065 2914.290 909.895 ;
      LAYER pwell ;
        RECT 5.665 905.675 5.835 905.845 ;
        RECT 2913.785 905.675 2913.955 905.845 ;
      LAYER nwell ;
        RECT 5.330 901.625 7.090 904.455 ;
        RECT 2912.530 901.625 2914.290 904.455 ;
      LAYER pwell ;
        RECT 5.665 900.235 5.835 900.405 ;
        RECT 2913.785 900.235 2913.955 900.405 ;
      LAYER nwell ;
        RECT 5.330 896.185 7.090 899.015 ;
        RECT 2912.530 896.185 2914.290 899.015 ;
      LAYER pwell ;
        RECT 5.665 894.795 5.835 894.965 ;
        RECT 2913.785 894.795 2913.955 894.965 ;
      LAYER nwell ;
        RECT 5.330 890.745 7.090 893.575 ;
        RECT 2912.530 890.745 2914.290 893.575 ;
      LAYER pwell ;
        RECT 5.665 889.355 5.835 889.525 ;
        RECT 2913.785 889.355 2913.955 889.525 ;
      LAYER nwell ;
        RECT 5.330 885.305 7.090 888.135 ;
        RECT 2912.530 885.305 2914.290 888.135 ;
      LAYER pwell ;
        RECT 5.665 883.915 5.835 884.085 ;
        RECT 2913.785 883.915 2913.955 884.085 ;
      LAYER nwell ;
        RECT 5.330 879.865 7.090 882.695 ;
        RECT 2912.530 879.865 2914.290 882.695 ;
      LAYER pwell ;
        RECT 5.665 878.475 5.835 878.645 ;
        RECT 2913.785 878.475 2913.955 878.645 ;
      LAYER nwell ;
        RECT 5.330 874.425 7.090 877.255 ;
        RECT 2912.530 874.425 2914.290 877.255 ;
      LAYER pwell ;
        RECT 5.665 873.035 5.835 873.205 ;
        RECT 2913.785 873.035 2913.955 873.205 ;
      LAYER nwell ;
        RECT 5.330 868.985 7.090 871.815 ;
        RECT 2912.530 868.985 2914.290 871.815 ;
      LAYER pwell ;
        RECT 5.665 867.595 5.835 867.765 ;
        RECT 2913.785 867.595 2913.955 867.765 ;
      LAYER nwell ;
        RECT 5.330 863.545 7.090 866.375 ;
        RECT 2912.530 863.545 2914.290 866.375 ;
      LAYER pwell ;
        RECT 5.665 862.155 5.835 862.325 ;
        RECT 2913.785 862.155 2913.955 862.325 ;
      LAYER nwell ;
        RECT 5.330 858.105 7.090 860.935 ;
        RECT 2912.530 858.105 2914.290 860.935 ;
      LAYER pwell ;
        RECT 5.665 856.715 5.835 856.885 ;
        RECT 2913.785 856.715 2913.955 856.885 ;
      LAYER nwell ;
        RECT 5.330 852.665 7.090 855.495 ;
        RECT 2912.530 852.665 2914.290 855.495 ;
      LAYER pwell ;
        RECT 5.665 851.275 5.835 851.445 ;
        RECT 2913.785 851.275 2913.955 851.445 ;
      LAYER nwell ;
        RECT 5.330 847.225 7.090 850.055 ;
        RECT 2912.530 847.225 2914.290 850.055 ;
      LAYER pwell ;
        RECT 5.665 845.835 5.835 846.005 ;
        RECT 2913.785 845.835 2913.955 846.005 ;
      LAYER nwell ;
        RECT 5.330 841.785 7.090 844.615 ;
        RECT 2912.530 841.785 2914.290 844.615 ;
      LAYER pwell ;
        RECT 5.665 840.395 5.835 840.565 ;
        RECT 2913.785 840.395 2913.955 840.565 ;
      LAYER nwell ;
        RECT 5.330 836.345 7.090 839.175 ;
        RECT 2912.530 836.345 2914.290 839.175 ;
      LAYER pwell ;
        RECT 5.665 834.955 5.835 835.125 ;
        RECT 2913.785 834.955 2913.955 835.125 ;
      LAYER nwell ;
        RECT 5.330 830.905 7.090 833.735 ;
        RECT 2912.530 830.905 2914.290 833.735 ;
      LAYER pwell ;
        RECT 5.665 829.515 5.835 829.685 ;
        RECT 2913.785 829.515 2913.955 829.685 ;
      LAYER nwell ;
        RECT 5.330 825.465 7.090 828.295 ;
        RECT 2912.530 825.465 2914.290 828.295 ;
      LAYER pwell ;
        RECT 5.665 824.075 5.835 824.245 ;
        RECT 2913.785 824.075 2913.955 824.245 ;
      LAYER nwell ;
        RECT 5.330 820.025 7.090 822.855 ;
        RECT 2912.530 820.025 2914.290 822.855 ;
      LAYER pwell ;
        RECT 5.665 818.635 5.835 818.805 ;
        RECT 2913.785 818.635 2913.955 818.805 ;
      LAYER nwell ;
        RECT 5.330 814.585 7.090 817.415 ;
        RECT 2912.530 814.585 2914.290 817.415 ;
      LAYER pwell ;
        RECT 5.665 813.195 5.835 813.365 ;
        RECT 2909.185 813.195 2909.355 813.365 ;
        RECT 2913.785 813.195 2913.955 813.365 ;
      LAYER nwell ;
        RECT 5.330 809.145 7.090 811.975 ;
        RECT 2912.530 809.145 2914.290 811.975 ;
      LAYER pwell ;
        RECT 5.665 807.755 5.835 807.925 ;
        RECT 2913.785 807.755 2913.955 807.925 ;
      LAYER nwell ;
        RECT 5.330 803.705 7.090 806.535 ;
        RECT 2912.530 803.705 2914.290 806.535 ;
      LAYER pwell ;
        RECT 5.665 802.315 5.835 802.485 ;
        RECT 2913.785 802.315 2913.955 802.485 ;
      LAYER nwell ;
        RECT 5.330 798.265 7.090 801.095 ;
        RECT 2912.530 798.265 2914.290 801.095 ;
      LAYER pwell ;
        RECT 5.665 796.875 5.835 797.045 ;
        RECT 2913.785 796.875 2913.955 797.045 ;
      LAYER nwell ;
        RECT 5.330 792.825 7.090 795.655 ;
        RECT 2912.530 792.825 2914.290 795.655 ;
      LAYER pwell ;
        RECT 5.665 791.435 5.835 791.605 ;
        RECT 2913.785 791.435 2913.955 791.605 ;
      LAYER nwell ;
        RECT 5.330 787.385 7.090 790.215 ;
        RECT 2912.530 787.385 2914.290 790.215 ;
      LAYER pwell ;
        RECT 5.665 785.995 5.835 786.165 ;
        RECT 2913.785 785.995 2913.955 786.165 ;
      LAYER nwell ;
        RECT 5.330 781.945 7.090 784.775 ;
        RECT 2912.530 781.945 2914.290 784.775 ;
      LAYER pwell ;
        RECT 5.665 780.555 5.835 780.725 ;
        RECT 2913.785 780.555 2913.955 780.725 ;
      LAYER nwell ;
        RECT 5.330 776.505 7.090 779.335 ;
        RECT 2912.530 776.505 2914.290 779.335 ;
      LAYER pwell ;
        RECT 5.665 775.115 5.835 775.285 ;
        RECT 2913.785 775.115 2913.955 775.285 ;
      LAYER nwell ;
        RECT 5.330 771.065 7.090 773.895 ;
        RECT 2912.530 771.065 2914.290 773.895 ;
      LAYER pwell ;
        RECT 5.665 769.675 5.835 769.845 ;
        RECT 2913.785 769.675 2913.955 769.845 ;
      LAYER nwell ;
        RECT 5.330 765.625 7.090 768.455 ;
        RECT 2912.530 765.625 2914.290 768.455 ;
      LAYER pwell ;
        RECT 5.665 764.235 5.835 764.405 ;
        RECT 2913.785 764.235 2913.955 764.405 ;
      LAYER nwell ;
        RECT 5.330 760.185 7.090 763.015 ;
        RECT 2912.530 760.185 2914.290 763.015 ;
      LAYER pwell ;
        RECT 5.665 758.795 5.835 758.965 ;
        RECT 2913.785 758.795 2913.955 758.965 ;
      LAYER nwell ;
        RECT 5.330 754.745 7.090 757.575 ;
        RECT 2912.530 754.745 2914.290 757.575 ;
      LAYER pwell ;
        RECT 5.665 753.355 5.835 753.525 ;
        RECT 2913.785 753.355 2913.955 753.525 ;
      LAYER nwell ;
        RECT 5.330 749.305 7.090 752.135 ;
        RECT 2912.530 749.305 2914.290 752.135 ;
      LAYER pwell ;
        RECT 5.665 747.915 5.835 748.085 ;
        RECT 2913.785 747.915 2913.955 748.085 ;
      LAYER nwell ;
        RECT 5.330 743.865 7.090 746.695 ;
        RECT 2912.530 743.865 2914.290 746.695 ;
      LAYER pwell ;
        RECT 5.665 742.475 5.835 742.645 ;
        RECT 2913.785 742.475 2913.955 742.645 ;
      LAYER nwell ;
        RECT 5.330 738.425 7.090 741.255 ;
        RECT 2912.530 738.425 2914.290 741.255 ;
      LAYER pwell ;
        RECT 5.665 737.035 5.835 737.205 ;
        RECT 2909.185 737.035 2909.355 737.205 ;
        RECT 2913.785 737.035 2913.955 737.205 ;
      LAYER nwell ;
        RECT 5.330 732.985 7.090 735.815 ;
        RECT 2912.530 732.985 2914.290 735.815 ;
      LAYER pwell ;
        RECT 5.665 731.595 5.835 731.765 ;
        RECT 2913.785 731.595 2913.955 731.765 ;
      LAYER nwell ;
        RECT 5.330 727.545 7.090 730.375 ;
        RECT 2912.530 727.545 2914.290 730.375 ;
      LAYER pwell ;
        RECT 5.665 726.155 5.835 726.325 ;
        RECT 2913.785 726.155 2913.955 726.325 ;
      LAYER nwell ;
        RECT 5.330 722.105 7.090 724.935 ;
        RECT 8.550 722.105 10.310 723.710 ;
        RECT 2912.530 722.105 2914.290 724.935 ;
      LAYER pwell ;
        RECT 5.665 720.715 5.835 720.885 ;
        RECT 8.885 720.715 9.055 720.885 ;
        RECT 2913.785 720.715 2913.955 720.885 ;
      LAYER nwell ;
        RECT 5.330 716.665 7.090 719.495 ;
        RECT 2912.530 716.665 2914.290 719.495 ;
      LAYER pwell ;
        RECT 5.665 715.275 5.835 715.445 ;
        RECT 2913.785 715.275 2913.955 715.445 ;
      LAYER nwell ;
        RECT 5.330 711.225 7.090 714.055 ;
        RECT 2912.530 711.225 2914.290 714.055 ;
      LAYER pwell ;
        RECT 5.665 709.835 5.835 710.005 ;
        RECT 2913.785 709.835 2913.955 710.005 ;
      LAYER nwell ;
        RECT 5.330 705.785 7.090 708.615 ;
        RECT 2912.530 705.785 2914.290 708.615 ;
      LAYER pwell ;
        RECT 5.665 704.395 5.835 704.565 ;
        RECT 2913.785 704.395 2913.955 704.565 ;
      LAYER nwell ;
        RECT 5.330 700.345 7.090 703.175 ;
        RECT 2912.530 700.345 2914.290 703.175 ;
      LAYER pwell ;
        RECT 5.665 698.955 5.835 699.125 ;
        RECT 2913.785 698.955 2913.955 699.125 ;
      LAYER nwell ;
        RECT 5.330 694.905 7.090 697.735 ;
        RECT 2912.530 694.905 2914.290 697.735 ;
      LAYER pwell ;
        RECT 5.665 693.515 5.835 693.685 ;
        RECT 2913.785 693.515 2913.955 693.685 ;
      LAYER nwell ;
        RECT 5.330 689.465 7.090 692.295 ;
        RECT 2912.530 689.465 2914.290 692.295 ;
      LAYER pwell ;
        RECT 5.665 688.075 5.835 688.245 ;
        RECT 2913.785 688.075 2913.955 688.245 ;
      LAYER nwell ;
        RECT 5.330 684.025 7.090 686.855 ;
        RECT 2912.530 684.025 2914.290 686.855 ;
      LAYER pwell ;
        RECT 5.665 682.635 5.835 682.805 ;
        RECT 2913.785 682.635 2913.955 682.805 ;
      LAYER nwell ;
        RECT 5.330 678.585 7.090 681.415 ;
        RECT 2912.530 678.585 2914.290 681.415 ;
      LAYER pwell ;
        RECT 5.665 677.195 5.835 677.365 ;
        RECT 2913.785 677.195 2913.955 677.365 ;
      LAYER nwell ;
        RECT 5.330 673.145 7.090 675.975 ;
        RECT 2912.530 673.145 2914.290 675.975 ;
      LAYER pwell ;
        RECT 5.665 671.755 5.835 671.925 ;
        RECT 2913.785 671.755 2913.955 671.925 ;
      LAYER nwell ;
        RECT 5.330 667.705 7.090 670.535 ;
        RECT 2912.530 667.705 2914.290 670.535 ;
      LAYER pwell ;
        RECT 5.665 666.315 5.835 666.485 ;
        RECT 2913.785 666.315 2913.955 666.485 ;
      LAYER nwell ;
        RECT 5.330 662.265 7.090 665.095 ;
        RECT 2912.530 662.265 2914.290 665.095 ;
      LAYER pwell ;
        RECT 5.665 660.875 5.835 661.045 ;
        RECT 2913.785 660.875 2913.955 661.045 ;
      LAYER nwell ;
        RECT 5.330 656.825 7.090 659.655 ;
        RECT 2912.530 656.825 2914.290 659.655 ;
      LAYER pwell ;
        RECT 5.665 655.435 5.835 655.605 ;
        RECT 2913.785 655.435 2913.955 655.605 ;
      LAYER nwell ;
        RECT 5.330 651.385 7.090 654.215 ;
        RECT 2912.530 651.385 2914.290 654.215 ;
      LAYER pwell ;
        RECT 5.665 649.995 5.835 650.165 ;
        RECT 2913.785 649.995 2913.955 650.165 ;
      LAYER nwell ;
        RECT 5.330 645.945 7.090 648.775 ;
        RECT 2912.530 645.945 2914.290 648.775 ;
      LAYER pwell ;
        RECT 5.665 644.555 5.835 644.725 ;
        RECT 2913.785 644.555 2913.955 644.725 ;
      LAYER nwell ;
        RECT 5.330 640.505 7.090 643.335 ;
        RECT 2912.530 640.505 2914.290 643.335 ;
      LAYER pwell ;
        RECT 5.665 639.115 5.835 639.285 ;
        RECT 2913.785 639.115 2913.955 639.285 ;
      LAYER nwell ;
        RECT 5.330 635.065 7.090 637.895 ;
        RECT 2912.530 635.065 2914.290 637.895 ;
      LAYER pwell ;
        RECT 5.665 633.675 5.835 633.845 ;
        RECT 2913.785 633.675 2913.955 633.845 ;
      LAYER nwell ;
        RECT 5.330 629.625 7.090 632.455 ;
        RECT 8.550 629.625 10.310 631.230 ;
        RECT 2912.530 629.625 2914.290 632.455 ;
      LAYER pwell ;
        RECT 5.665 628.235 5.835 628.405 ;
        RECT 8.885 628.235 9.055 628.405 ;
        RECT 2913.785 628.235 2913.955 628.405 ;
      LAYER nwell ;
        RECT 5.330 624.185 7.090 627.015 ;
        RECT 2912.530 624.185 2914.290 627.015 ;
      LAYER pwell ;
        RECT 5.665 622.795 5.835 622.965 ;
        RECT 2913.785 622.795 2913.955 622.965 ;
      LAYER nwell ;
        RECT 5.330 618.745 7.090 621.575 ;
        RECT 2912.530 618.745 2914.290 621.575 ;
      LAYER pwell ;
        RECT 5.665 617.355 5.835 617.525 ;
        RECT 2913.785 617.355 2913.955 617.525 ;
      LAYER nwell ;
        RECT 5.330 613.305 7.090 616.135 ;
        RECT 2912.530 613.305 2914.290 616.135 ;
      LAYER pwell ;
        RECT 5.665 611.915 5.835 612.085 ;
        RECT 2913.785 611.915 2913.955 612.085 ;
      LAYER nwell ;
        RECT 5.330 607.865 7.090 610.695 ;
        RECT 2912.530 607.865 2914.290 610.695 ;
      LAYER pwell ;
        RECT 5.665 606.475 5.835 606.645 ;
        RECT 2913.785 606.475 2913.955 606.645 ;
      LAYER nwell ;
        RECT 5.330 602.425 7.090 605.255 ;
        RECT 8.550 602.425 10.310 604.030 ;
        RECT 2912.530 602.425 2914.290 605.255 ;
      LAYER pwell ;
        RECT 5.665 601.035 5.835 601.205 ;
        RECT 8.885 601.035 9.055 601.205 ;
        RECT 2913.785 601.035 2913.955 601.205 ;
      LAYER nwell ;
        RECT 5.330 596.985 7.090 599.815 ;
        RECT 2912.530 596.985 2914.290 599.815 ;
      LAYER pwell ;
        RECT 5.665 595.595 5.835 595.765 ;
        RECT 2913.785 595.595 2913.955 595.765 ;
      LAYER nwell ;
        RECT 5.330 591.545 7.090 594.375 ;
        RECT 2912.530 591.545 2914.290 594.375 ;
      LAYER pwell ;
        RECT 5.665 590.155 5.835 590.325 ;
        RECT 2913.785 590.155 2913.955 590.325 ;
      LAYER nwell ;
        RECT 5.330 586.105 7.090 588.935 ;
        RECT 2912.530 586.105 2914.290 588.935 ;
      LAYER pwell ;
        RECT 5.665 584.715 5.835 584.885 ;
        RECT 2913.785 584.715 2913.955 584.885 ;
      LAYER nwell ;
        RECT 5.330 580.665 7.090 583.495 ;
        RECT 2912.530 580.665 2914.290 583.495 ;
      LAYER pwell ;
        RECT 5.665 579.275 5.835 579.445 ;
        RECT 2913.785 579.275 2913.955 579.445 ;
      LAYER nwell ;
        RECT 5.330 575.225 7.090 578.055 ;
        RECT 2912.530 575.225 2914.290 578.055 ;
      LAYER pwell ;
        RECT 5.665 573.835 5.835 574.005 ;
        RECT 2913.785 573.835 2913.955 574.005 ;
      LAYER nwell ;
        RECT 5.330 569.785 7.090 572.615 ;
        RECT 2912.530 569.785 2914.290 572.615 ;
      LAYER pwell ;
        RECT 5.665 568.395 5.835 568.565 ;
        RECT 2913.785 568.395 2913.955 568.565 ;
      LAYER nwell ;
        RECT 5.330 564.345 7.090 567.175 ;
        RECT 2912.530 564.345 2914.290 567.175 ;
      LAYER pwell ;
        RECT 5.665 562.955 5.835 563.125 ;
        RECT 2913.785 562.955 2913.955 563.125 ;
      LAYER nwell ;
        RECT 5.330 558.905 7.090 561.735 ;
        RECT 2912.530 558.905 2914.290 561.735 ;
      LAYER pwell ;
        RECT 5.665 557.515 5.835 557.685 ;
        RECT 2913.785 557.515 2913.955 557.685 ;
      LAYER nwell ;
        RECT 5.330 553.465 7.090 556.295 ;
        RECT 2912.530 553.465 2914.290 556.295 ;
      LAYER pwell ;
        RECT 5.665 552.075 5.835 552.245 ;
        RECT 2913.785 552.075 2913.955 552.245 ;
      LAYER nwell ;
        RECT 5.330 548.025 7.090 550.855 ;
        RECT 2912.530 548.025 2914.290 550.855 ;
      LAYER pwell ;
        RECT 5.665 546.635 5.835 546.805 ;
        RECT 2913.785 546.635 2913.955 546.805 ;
      LAYER nwell ;
        RECT 5.330 542.585 7.090 545.415 ;
        RECT 2912.530 542.585 2914.290 545.415 ;
      LAYER pwell ;
        RECT 5.665 541.195 5.835 541.365 ;
        RECT 2913.785 541.195 2913.955 541.365 ;
      LAYER nwell ;
        RECT 5.330 537.145 7.090 539.975 ;
        RECT 2912.530 537.145 2914.290 539.975 ;
      LAYER pwell ;
        RECT 5.665 535.755 5.835 535.925 ;
        RECT 2913.785 535.755 2913.955 535.925 ;
      LAYER nwell ;
        RECT 5.330 531.705 7.090 534.535 ;
        RECT 2912.530 531.705 2914.290 534.535 ;
      LAYER pwell ;
        RECT 5.665 530.315 5.835 530.485 ;
        RECT 2913.785 530.315 2913.955 530.485 ;
      LAYER nwell ;
        RECT 5.330 526.265 7.090 529.095 ;
        RECT 2912.530 526.265 2914.290 529.095 ;
      LAYER pwell ;
        RECT 5.665 524.875 5.835 525.045 ;
        RECT 2913.785 524.875 2913.955 525.045 ;
      LAYER nwell ;
        RECT 5.330 520.825 7.090 523.655 ;
        RECT 2912.530 520.825 2914.290 523.655 ;
      LAYER pwell ;
        RECT 5.665 519.435 5.835 519.605 ;
        RECT 2913.785 519.435 2913.955 519.605 ;
      LAYER nwell ;
        RECT 5.330 515.385 7.090 518.215 ;
        RECT 2912.530 515.385 2914.290 518.215 ;
      LAYER pwell ;
        RECT 5.665 513.995 5.835 514.165 ;
        RECT 2913.785 513.995 2913.955 514.165 ;
      LAYER nwell ;
        RECT 5.330 509.945 7.090 512.775 ;
        RECT 2912.530 509.945 2914.290 512.775 ;
      LAYER pwell ;
        RECT 5.665 508.555 5.835 508.725 ;
        RECT 2913.785 508.555 2913.955 508.725 ;
      LAYER nwell ;
        RECT 5.330 504.505 7.090 507.335 ;
        RECT 2912.530 504.505 2914.290 507.335 ;
      LAYER pwell ;
        RECT 5.665 503.115 5.835 503.285 ;
        RECT 2913.785 503.115 2913.955 503.285 ;
      LAYER nwell ;
        RECT 5.330 499.065 7.090 501.895 ;
        RECT 2912.530 499.065 2914.290 501.895 ;
      LAYER pwell ;
        RECT 5.665 497.675 5.835 497.845 ;
        RECT 2913.785 497.675 2913.955 497.845 ;
      LAYER nwell ;
        RECT 5.330 493.625 7.090 496.455 ;
        RECT 2912.530 493.625 2914.290 496.455 ;
      LAYER pwell ;
        RECT 5.665 492.235 5.835 492.405 ;
        RECT 2913.785 492.235 2913.955 492.405 ;
      LAYER nwell ;
        RECT 5.330 488.185 7.090 491.015 ;
        RECT 2912.530 488.185 2914.290 491.015 ;
      LAYER pwell ;
        RECT 5.665 486.795 5.835 486.965 ;
        RECT 2913.785 486.795 2913.955 486.965 ;
      LAYER nwell ;
        RECT 5.330 482.745 7.090 485.575 ;
        RECT 2912.530 482.745 2914.290 485.575 ;
      LAYER pwell ;
        RECT 5.665 481.355 5.835 481.525 ;
        RECT 2913.785 481.355 2913.955 481.525 ;
      LAYER nwell ;
        RECT 5.330 477.305 7.090 480.135 ;
        RECT 2912.530 477.305 2914.290 480.135 ;
      LAYER pwell ;
        RECT 5.665 475.915 5.835 476.085 ;
        RECT 2913.785 475.915 2913.955 476.085 ;
      LAYER nwell ;
        RECT 5.330 471.865 7.090 474.695 ;
        RECT 2912.530 471.865 2914.290 474.695 ;
      LAYER pwell ;
        RECT 5.665 470.475 5.835 470.645 ;
        RECT 2909.185 470.475 2909.355 470.645 ;
        RECT 2913.785 470.475 2913.955 470.645 ;
      LAYER nwell ;
        RECT 5.330 466.425 7.090 469.255 ;
        RECT 2912.530 466.425 2914.290 469.255 ;
      LAYER pwell ;
        RECT 5.665 465.035 5.835 465.205 ;
        RECT 2913.785 465.035 2913.955 465.205 ;
      LAYER nwell ;
        RECT 5.330 460.985 7.090 463.815 ;
        RECT 2912.530 460.985 2914.290 463.815 ;
      LAYER pwell ;
        RECT 5.665 459.595 5.835 459.765 ;
        RECT 2913.785 459.595 2913.955 459.765 ;
      LAYER nwell ;
        RECT 5.330 455.545 7.090 458.375 ;
        RECT 2912.530 455.545 2914.290 458.375 ;
      LAYER pwell ;
        RECT 5.665 454.155 5.835 454.325 ;
        RECT 2913.785 454.155 2913.955 454.325 ;
      LAYER nwell ;
        RECT 5.330 450.105 7.090 452.935 ;
        RECT 2912.530 450.105 2914.290 452.935 ;
      LAYER pwell ;
        RECT 5.665 448.715 5.835 448.885 ;
        RECT 2910.565 448.715 2910.735 448.885 ;
        RECT 2913.785 448.715 2913.955 448.885 ;
      LAYER nwell ;
        RECT 5.330 444.665 7.090 447.495 ;
        RECT 2912.530 444.665 2914.290 447.495 ;
      LAYER pwell ;
        RECT 5.665 443.275 5.835 443.445 ;
        RECT 8.885 443.275 9.055 443.445 ;
        RECT 2913.785 443.275 2913.955 443.445 ;
      LAYER nwell ;
        RECT 5.330 439.225 7.090 442.055 ;
        RECT 8.550 439.225 10.310 442.055 ;
        RECT 2912.530 439.225 2914.290 442.055 ;
      LAYER pwell ;
        RECT 5.665 437.835 5.835 438.005 ;
        RECT 8.885 437.835 9.055 438.005 ;
        RECT 2913.785 437.835 2913.955 438.005 ;
      LAYER nwell ;
        RECT 5.330 433.785 7.090 436.615 ;
        RECT 2912.530 433.785 2914.290 436.615 ;
      LAYER pwell ;
        RECT 5.665 432.395 5.835 432.565 ;
        RECT 2913.785 432.395 2913.955 432.565 ;
      LAYER nwell ;
        RECT 5.330 428.345 7.090 431.175 ;
        RECT 2912.530 428.345 2914.290 431.175 ;
      LAYER pwell ;
        RECT 5.665 426.955 5.835 427.125 ;
        RECT 2913.785 426.955 2913.955 427.125 ;
      LAYER nwell ;
        RECT 5.330 422.905 7.090 425.735 ;
        RECT 2912.530 422.905 2914.290 425.735 ;
      LAYER pwell ;
        RECT 5.665 421.515 5.835 421.685 ;
        RECT 2913.785 421.515 2913.955 421.685 ;
      LAYER nwell ;
        RECT 5.330 417.465 7.090 420.295 ;
        RECT 2912.530 417.465 2914.290 420.295 ;
      LAYER pwell ;
        RECT 5.665 416.075 5.835 416.245 ;
        RECT 2913.785 416.075 2913.955 416.245 ;
      LAYER nwell ;
        RECT 5.330 412.025 7.090 414.855 ;
        RECT 2912.530 412.025 2914.290 414.855 ;
      LAYER pwell ;
        RECT 5.665 410.635 5.835 410.805 ;
        RECT 2913.785 410.635 2913.955 410.805 ;
      LAYER nwell ;
        RECT 5.330 406.585 7.090 409.415 ;
        RECT 2912.530 406.585 2914.290 409.415 ;
      LAYER pwell ;
        RECT 5.665 405.195 5.835 405.365 ;
        RECT 2913.785 405.195 2913.955 405.365 ;
      LAYER nwell ;
        RECT 5.330 401.145 7.090 403.975 ;
        RECT 8.550 401.145 10.310 402.750 ;
        RECT 2912.530 401.145 2914.290 403.975 ;
      LAYER pwell ;
        RECT 5.665 399.755 5.835 399.925 ;
        RECT 8.885 399.755 9.055 399.925 ;
        RECT 2913.785 399.755 2913.955 399.925 ;
      LAYER nwell ;
        RECT 5.330 395.705 7.090 398.535 ;
        RECT 2912.530 395.705 2914.290 398.535 ;
      LAYER pwell ;
        RECT 5.665 394.315 5.835 394.485 ;
        RECT 8.885 394.315 9.055 394.485 ;
        RECT 2913.785 394.315 2913.955 394.485 ;
      LAYER nwell ;
        RECT 5.330 390.265 7.090 393.095 ;
        RECT 8.550 391.490 10.310 393.095 ;
        RECT 2912.530 390.265 2914.290 393.095 ;
      LAYER pwell ;
        RECT 5.665 388.875 5.835 389.045 ;
        RECT 2913.785 388.875 2913.955 389.045 ;
      LAYER nwell ;
        RECT 5.330 384.825 7.090 387.655 ;
        RECT 2912.530 384.825 2914.290 387.655 ;
      LAYER pwell ;
        RECT 5.665 383.435 5.835 383.605 ;
        RECT 2913.785 383.435 2913.955 383.605 ;
      LAYER nwell ;
        RECT 5.330 379.385 7.090 382.215 ;
        RECT 2912.530 379.385 2914.290 382.215 ;
      LAYER pwell ;
        RECT 5.665 377.995 5.835 378.165 ;
        RECT 2913.785 377.995 2913.955 378.165 ;
      LAYER nwell ;
        RECT 5.330 373.945 7.090 376.775 ;
        RECT 2912.530 373.945 2914.290 376.775 ;
      LAYER pwell ;
        RECT 5.665 372.555 5.835 372.725 ;
        RECT 2913.785 372.555 2913.955 372.725 ;
      LAYER nwell ;
        RECT 5.330 368.505 7.090 371.335 ;
        RECT 2912.530 368.505 2914.290 371.335 ;
      LAYER pwell ;
        RECT 5.665 367.115 5.835 367.285 ;
        RECT 2913.785 367.115 2913.955 367.285 ;
      LAYER nwell ;
        RECT 5.330 363.065 7.090 365.895 ;
        RECT 2912.530 363.065 2914.290 365.895 ;
      LAYER pwell ;
        RECT 5.665 361.675 5.835 361.845 ;
        RECT 2913.785 361.675 2913.955 361.845 ;
      LAYER nwell ;
        RECT 5.330 357.625 7.090 360.455 ;
        RECT 2912.530 357.625 2914.290 360.455 ;
      LAYER pwell ;
        RECT 5.665 356.235 5.835 356.405 ;
        RECT 2913.785 356.235 2913.955 356.405 ;
      LAYER nwell ;
        RECT 5.330 352.185 7.090 355.015 ;
        RECT 2912.530 352.185 2914.290 355.015 ;
      LAYER pwell ;
        RECT 5.665 350.795 5.835 350.965 ;
        RECT 2913.785 350.795 2913.955 350.965 ;
      LAYER nwell ;
        RECT 5.330 346.745 7.090 349.575 ;
        RECT 2912.530 346.745 2914.290 349.575 ;
      LAYER pwell ;
        RECT 5.665 345.355 5.835 345.525 ;
        RECT 2913.785 345.355 2913.955 345.525 ;
      LAYER nwell ;
        RECT 5.330 341.305 7.090 344.135 ;
        RECT 2912.530 341.305 2914.290 344.135 ;
      LAYER pwell ;
        RECT 5.665 339.915 5.835 340.085 ;
        RECT 2913.785 339.915 2913.955 340.085 ;
      LAYER nwell ;
        RECT 5.330 335.865 7.090 338.695 ;
        RECT 2912.530 335.865 2914.290 338.695 ;
      LAYER pwell ;
        RECT 5.665 334.475 5.835 334.645 ;
        RECT 2913.785 334.475 2913.955 334.645 ;
      LAYER nwell ;
        RECT 5.330 330.425 7.090 333.255 ;
        RECT 2912.530 330.425 2914.290 333.255 ;
      LAYER pwell ;
        RECT 5.665 329.035 5.835 329.205 ;
        RECT 2913.785 329.035 2913.955 329.205 ;
      LAYER nwell ;
        RECT 5.330 324.985 7.090 327.815 ;
        RECT 2912.530 324.985 2914.290 327.815 ;
      LAYER pwell ;
        RECT 5.665 323.595 5.835 323.765 ;
        RECT 2913.785 323.595 2913.955 323.765 ;
      LAYER nwell ;
        RECT 5.330 319.545 7.090 322.375 ;
        RECT 2912.530 319.545 2914.290 322.375 ;
      LAYER pwell ;
        RECT 5.665 318.155 5.835 318.325 ;
        RECT 2913.785 318.155 2913.955 318.325 ;
      LAYER nwell ;
        RECT 5.330 314.105 7.090 316.935 ;
        RECT 8.550 314.105 10.310 315.710 ;
        RECT 2912.530 314.105 2914.290 316.935 ;
      LAYER pwell ;
        RECT 5.665 312.715 5.835 312.885 ;
        RECT 8.885 312.715 9.055 312.885 ;
        RECT 2913.785 312.715 2913.955 312.885 ;
      LAYER nwell ;
        RECT 5.330 308.665 7.090 311.495 ;
        RECT 2912.530 308.665 2914.290 311.495 ;
      LAYER pwell ;
        RECT 5.665 307.275 5.835 307.445 ;
        RECT 2913.785 307.275 2913.955 307.445 ;
      LAYER nwell ;
        RECT 5.330 303.225 7.090 306.055 ;
        RECT 2912.530 303.225 2914.290 306.055 ;
      LAYER pwell ;
        RECT 5.665 301.835 5.835 302.005 ;
        RECT 2913.785 301.835 2913.955 302.005 ;
      LAYER nwell ;
        RECT 5.330 297.785 7.090 300.615 ;
        RECT 2912.530 297.785 2914.290 300.615 ;
      LAYER pwell ;
        RECT 5.665 296.395 5.835 296.565 ;
        RECT 2913.785 296.395 2913.955 296.565 ;
      LAYER nwell ;
        RECT 5.330 292.345 7.090 295.175 ;
        RECT 2912.530 292.345 2914.290 295.175 ;
      LAYER pwell ;
        RECT 5.665 290.955 5.835 291.125 ;
        RECT 2909.185 290.955 2909.355 291.125 ;
        RECT 2913.785 290.955 2913.955 291.125 ;
      LAYER nwell ;
        RECT 5.330 286.905 7.090 289.735 ;
        RECT 2912.530 286.905 2914.290 289.735 ;
      LAYER pwell ;
        RECT 5.665 285.515 5.835 285.685 ;
        RECT 2913.785 285.515 2913.955 285.685 ;
      LAYER nwell ;
        RECT 5.330 281.465 7.090 284.295 ;
        RECT 2912.530 281.465 2914.290 284.295 ;
      LAYER pwell ;
        RECT 5.665 280.075 5.835 280.245 ;
        RECT 2913.785 280.075 2913.955 280.245 ;
      LAYER nwell ;
        RECT 5.330 276.025 7.090 278.855 ;
        RECT 2912.530 276.025 2914.290 278.855 ;
      LAYER pwell ;
        RECT 5.665 274.635 5.835 274.805 ;
        RECT 2913.785 274.635 2913.955 274.805 ;
      LAYER nwell ;
        RECT 5.330 270.585 7.090 273.415 ;
        RECT 2912.530 270.585 2914.290 273.415 ;
      LAYER pwell ;
        RECT 5.665 269.195 5.835 269.365 ;
        RECT 2913.785 269.195 2913.955 269.365 ;
      LAYER nwell ;
        RECT 5.330 265.145 7.090 267.975 ;
        RECT 2912.530 265.145 2914.290 267.975 ;
      LAYER pwell ;
        RECT 5.665 263.755 5.835 263.925 ;
        RECT 2913.785 263.755 2913.955 263.925 ;
      LAYER nwell ;
        RECT 5.330 259.705 7.090 262.535 ;
        RECT 2912.530 259.705 2914.290 262.535 ;
      LAYER pwell ;
        RECT 5.665 258.315 5.835 258.485 ;
        RECT 2913.785 258.315 2913.955 258.485 ;
      LAYER nwell ;
        RECT 5.330 254.265 7.090 257.095 ;
        RECT 2912.530 254.265 2914.290 257.095 ;
      LAYER pwell ;
        RECT 5.665 252.875 5.835 253.045 ;
        RECT 2913.785 252.875 2913.955 253.045 ;
      LAYER nwell ;
        RECT 5.330 248.825 7.090 251.655 ;
        RECT 2912.530 248.825 2914.290 251.655 ;
      LAYER pwell ;
        RECT 5.665 247.435 5.835 247.605 ;
        RECT 2913.785 247.435 2913.955 247.605 ;
      LAYER nwell ;
        RECT 5.330 243.385 7.090 246.215 ;
        RECT 2912.530 243.385 2914.290 246.215 ;
      LAYER pwell ;
        RECT 5.665 241.995 5.835 242.165 ;
        RECT 2913.785 241.995 2913.955 242.165 ;
      LAYER nwell ;
        RECT 5.330 237.945 7.090 240.775 ;
        RECT 2912.530 237.945 2914.290 240.775 ;
      LAYER pwell ;
        RECT 5.665 236.555 5.835 236.725 ;
        RECT 2913.785 236.555 2913.955 236.725 ;
      LAYER nwell ;
        RECT 5.330 232.505 7.090 235.335 ;
        RECT 2912.530 232.505 2914.290 235.335 ;
      LAYER pwell ;
        RECT 5.665 231.115 5.835 231.285 ;
        RECT 2910.565 231.115 2910.735 231.285 ;
        RECT 2913.785 231.115 2913.955 231.285 ;
      LAYER nwell ;
        RECT 5.330 227.065 7.090 229.895 ;
        RECT 2912.530 227.065 2914.290 229.895 ;
      LAYER pwell ;
        RECT 5.665 225.675 5.835 225.845 ;
        RECT 2913.785 225.675 2913.955 225.845 ;
      LAYER nwell ;
        RECT 5.330 221.625 7.090 224.455 ;
        RECT 2912.530 221.625 2914.290 224.455 ;
      LAYER pwell ;
        RECT 5.665 220.235 5.835 220.405 ;
        RECT 2913.785 220.235 2913.955 220.405 ;
      LAYER nwell ;
        RECT 5.330 216.185 7.090 219.015 ;
        RECT 2912.530 216.185 2914.290 219.015 ;
      LAYER pwell ;
        RECT 5.665 214.795 5.835 214.965 ;
        RECT 2913.785 214.795 2913.955 214.965 ;
      LAYER nwell ;
        RECT 5.330 210.745 7.090 213.575 ;
        RECT 2912.530 210.745 2914.290 213.575 ;
      LAYER pwell ;
        RECT 5.665 209.355 5.835 209.525 ;
        RECT 2913.785 209.355 2913.955 209.525 ;
      LAYER nwell ;
        RECT 5.330 205.305 7.090 208.135 ;
        RECT 2912.530 205.305 2914.290 208.135 ;
      LAYER pwell ;
        RECT 5.665 203.915 5.835 204.085 ;
        RECT 2913.785 203.915 2913.955 204.085 ;
      LAYER nwell ;
        RECT 5.330 199.865 7.090 202.695 ;
        RECT 2912.530 199.865 2914.290 202.695 ;
      LAYER pwell ;
        RECT 5.665 198.475 5.835 198.645 ;
        RECT 2913.785 198.475 2913.955 198.645 ;
      LAYER nwell ;
        RECT 5.330 194.425 7.090 197.255 ;
        RECT 2912.530 194.425 2914.290 197.255 ;
      LAYER pwell ;
        RECT 5.665 193.035 5.835 193.205 ;
        RECT 2913.785 193.035 2913.955 193.205 ;
      LAYER nwell ;
        RECT 5.330 188.985 7.090 191.815 ;
        RECT 2912.530 188.985 2914.290 191.815 ;
      LAYER pwell ;
        RECT 5.665 187.595 5.835 187.765 ;
        RECT 2913.785 187.595 2913.955 187.765 ;
      LAYER nwell ;
        RECT 5.330 183.545 7.090 186.375 ;
        RECT 2912.530 183.545 2914.290 186.375 ;
      LAYER pwell ;
        RECT 5.665 182.155 5.835 182.325 ;
        RECT 2913.785 182.155 2913.955 182.325 ;
      LAYER nwell ;
        RECT 5.330 178.105 7.090 180.935 ;
        RECT 2912.530 178.105 2914.290 180.935 ;
      LAYER pwell ;
        RECT 5.665 176.715 5.835 176.885 ;
        RECT 2913.785 176.715 2913.955 176.885 ;
      LAYER nwell ;
        RECT 5.330 172.665 7.090 175.495 ;
        RECT 2912.530 172.665 2914.290 175.495 ;
      LAYER pwell ;
        RECT 5.665 171.275 5.835 171.445 ;
        RECT 2913.785 171.275 2913.955 171.445 ;
      LAYER nwell ;
        RECT 5.330 167.225 7.090 170.055 ;
        RECT 2912.530 167.225 2914.290 170.055 ;
      LAYER pwell ;
        RECT 5.665 165.835 5.835 166.005 ;
        RECT 2913.785 165.835 2913.955 166.005 ;
      LAYER nwell ;
        RECT 5.330 161.785 7.090 164.615 ;
        RECT 2912.530 161.785 2914.290 164.615 ;
      LAYER pwell ;
        RECT 5.665 160.395 5.835 160.565 ;
        RECT 2913.785 160.395 2913.955 160.565 ;
      LAYER nwell ;
        RECT 5.330 156.345 7.090 159.175 ;
        RECT 2912.530 156.345 2914.290 159.175 ;
      LAYER pwell ;
        RECT 5.665 154.955 5.835 155.125 ;
        RECT 2913.785 154.955 2913.955 155.125 ;
      LAYER nwell ;
        RECT 5.330 150.905 7.090 153.735 ;
        RECT 2912.530 150.905 2914.290 153.735 ;
      LAYER pwell ;
        RECT 5.665 149.515 5.835 149.685 ;
        RECT 2913.785 149.515 2913.955 149.685 ;
      LAYER nwell ;
        RECT 5.330 145.465 7.090 148.295 ;
        RECT 2912.530 145.465 2914.290 148.295 ;
      LAYER pwell ;
        RECT 5.665 144.075 5.835 144.245 ;
        RECT 2913.785 144.075 2913.955 144.245 ;
      LAYER nwell ;
        RECT 5.330 140.025 7.090 142.855 ;
        RECT 2912.530 140.025 2914.290 142.855 ;
      LAYER pwell ;
        RECT 5.665 138.635 5.835 138.805 ;
        RECT 2913.785 138.635 2913.955 138.805 ;
      LAYER nwell ;
        RECT 5.330 134.585 7.090 137.415 ;
        RECT 2912.530 134.585 2914.290 137.415 ;
      LAYER pwell ;
        RECT 5.665 133.195 5.835 133.365 ;
        RECT 2913.785 133.195 2913.955 133.365 ;
      LAYER nwell ;
        RECT 5.330 129.145 7.090 131.975 ;
        RECT 2912.530 129.145 2914.290 131.975 ;
      LAYER pwell ;
        RECT 5.665 127.755 5.835 127.925 ;
        RECT 7.045 127.755 7.215 127.925 ;
        RECT 2913.785 127.755 2913.955 127.925 ;
      LAYER nwell ;
        RECT 5.330 124.930 15.830 126.535 ;
        RECT 5.330 123.705 7.090 124.930 ;
        RECT 2912.530 123.705 2914.290 126.535 ;
      LAYER pwell ;
        RECT 5.665 122.315 5.835 122.485 ;
        RECT 2913.785 122.315 2913.955 122.485 ;
      LAYER nwell ;
        RECT 5.330 118.265 7.090 121.095 ;
        RECT 2912.530 118.265 2914.290 121.095 ;
      LAYER pwell ;
        RECT 5.665 116.875 5.835 117.045 ;
        RECT 2913.785 116.875 2913.955 117.045 ;
      LAYER nwell ;
        RECT 5.330 112.825 7.090 115.655 ;
        RECT 2912.530 112.825 2914.290 115.655 ;
      LAYER pwell ;
        RECT 5.665 111.435 5.835 111.605 ;
        RECT 2913.785 111.435 2913.955 111.605 ;
      LAYER nwell ;
        RECT 5.330 107.385 7.090 110.215 ;
        RECT 2912.530 107.385 2914.290 110.215 ;
      LAYER pwell ;
        RECT 5.665 105.995 5.835 106.165 ;
        RECT 8.885 105.995 9.055 106.165 ;
        RECT 2913.785 105.995 2913.955 106.165 ;
      LAYER nwell ;
        RECT 5.330 101.945 7.090 104.775 ;
        RECT 8.550 103.170 10.310 104.775 ;
        RECT 2912.530 101.945 2914.290 104.775 ;
      LAYER pwell ;
        RECT 5.665 100.555 5.835 100.725 ;
        RECT 2913.785 100.555 2913.955 100.725 ;
      LAYER nwell ;
        RECT 5.330 96.505 7.090 99.335 ;
        RECT 2912.530 96.505 2914.290 99.335 ;
      LAYER pwell ;
        RECT 5.665 95.115 5.835 95.285 ;
        RECT 2913.785 95.115 2913.955 95.285 ;
      LAYER nwell ;
        RECT 5.330 91.065 7.090 93.895 ;
        RECT 2912.530 91.065 2914.290 93.895 ;
      LAYER pwell ;
        RECT 5.665 89.675 5.835 89.845 ;
        RECT 2913.785 89.675 2913.955 89.845 ;
      LAYER nwell ;
        RECT 5.330 85.625 7.090 88.455 ;
        RECT 2912.530 85.625 2914.290 88.455 ;
      LAYER pwell ;
        RECT 5.665 84.235 5.835 84.405 ;
        RECT 2913.785 84.235 2913.955 84.405 ;
      LAYER nwell ;
        RECT 5.330 80.185 7.090 83.015 ;
        RECT 2912.530 80.185 2914.290 83.015 ;
      LAYER pwell ;
        RECT 5.665 78.795 5.835 78.965 ;
        RECT 2913.785 78.795 2913.955 78.965 ;
      LAYER nwell ;
        RECT 5.330 74.745 7.090 77.575 ;
        RECT 2912.530 74.745 2914.290 77.575 ;
      LAYER pwell ;
        RECT 5.665 73.355 5.835 73.525 ;
        RECT 2913.785 73.355 2913.955 73.525 ;
      LAYER nwell ;
        RECT 5.330 69.305 7.090 72.135 ;
        RECT 2912.530 69.305 2914.290 72.135 ;
      LAYER pwell ;
        RECT 5.665 67.915 5.835 68.085 ;
        RECT 2913.785 67.915 2913.955 68.085 ;
      LAYER nwell ;
        RECT 5.330 63.865 7.090 66.695 ;
        RECT 2912.530 63.865 2914.290 66.695 ;
      LAYER pwell ;
        RECT 5.665 62.475 5.835 62.645 ;
        RECT 2909.185 62.475 2909.355 62.645 ;
        RECT 2913.785 62.475 2913.955 62.645 ;
      LAYER nwell ;
        RECT 5.330 58.425 7.090 61.255 ;
        RECT 2912.530 58.425 2914.290 61.255 ;
      LAYER pwell ;
        RECT 5.665 57.035 5.835 57.205 ;
        RECT 2913.785 57.035 2913.955 57.205 ;
      LAYER nwell ;
        RECT 5.330 52.985 7.090 55.815 ;
        RECT 2912.530 52.985 2914.290 55.815 ;
      LAYER pwell ;
        RECT 5.665 51.595 5.835 51.765 ;
        RECT 2913.785 51.595 2913.955 51.765 ;
      LAYER nwell ;
        RECT 5.330 47.545 7.090 50.375 ;
        RECT 2912.530 47.545 2914.290 50.375 ;
      LAYER pwell ;
        RECT 5.665 46.155 5.835 46.325 ;
        RECT 2913.785 46.155 2913.955 46.325 ;
      LAYER nwell ;
        RECT 5.330 43.710 7.090 44.935 ;
        RECT 5.330 42.105 15.830 43.710 ;
        RECT 2912.530 42.105 2914.290 44.935 ;
      LAYER pwell ;
        RECT 5.665 40.715 5.835 40.885 ;
        RECT 7.045 40.715 7.215 40.885 ;
        RECT 2913.785 40.715 2913.955 40.885 ;
      LAYER nwell ;
        RECT 5.330 36.665 7.090 39.495 ;
        RECT 2912.530 36.665 2914.290 39.495 ;
      LAYER pwell ;
        RECT 5.665 35.275 5.835 35.445 ;
        RECT 2913.785 35.275 2913.955 35.445 ;
      LAYER nwell ;
        RECT 5.330 31.225 7.090 34.055 ;
        RECT 2912.530 31.225 2914.290 34.055 ;
      LAYER pwell ;
        RECT 5.665 29.835 5.835 30.005 ;
        RECT 2913.785 29.835 2913.955 30.005 ;
      LAYER nwell ;
        RECT 5.330 25.785 7.090 28.615 ;
        RECT 2912.530 25.785 2914.290 28.615 ;
      LAYER pwell ;
        RECT 5.665 24.395 5.835 24.565 ;
        RECT 2913.785 24.395 2913.955 24.565 ;
      LAYER nwell ;
        RECT 5.330 21.950 7.090 23.175 ;
        RECT 5.330 20.345 14.450 21.950 ;
        RECT 2912.530 20.345 2914.290 23.175 ;
      LAYER pwell ;
        RECT 5.665 18.955 5.835 19.125 ;
        RECT 7.045 18.955 7.220 19.125 ;
        RECT 2909.185 18.955 2909.355 19.125 ;
        RECT 2910.565 18.955 2910.735 19.125 ;
        RECT 2913.785 18.955 2913.955 19.125 ;
      LAYER nwell ;
        RECT 5.330 14.905 15.830 17.735 ;
        RECT 2912.530 14.905 2914.290 17.735 ;
      LAYER pwell ;
        RECT 5.665 13.515 5.835 13.685 ;
        RECT 7.045 13.515 7.215 13.685 ;
        RECT 8.885 13.515 9.055 13.685 ;
        RECT 10.265 13.515 10.435 13.685 ;
        RECT 16.705 13.515 16.875 13.685 ;
        RECT 58.105 13.515 58.275 13.685 ;
        RECT 59.485 13.515 59.655 13.685 ;
        RECT 77.425 13.515 77.595 13.685 ;
        RECT 82.025 13.515 82.195 13.685 ;
        RECT 82.945 13.515 83.115 13.685 ;
        RECT 101.345 13.515 101.515 13.685 ;
        RECT 104.570 13.515 104.740 13.685 ;
        RECT 120.205 13.515 120.375 13.685 ;
        RECT 134.465 13.515 134.635 13.685 ;
        RECT 142.290 13.515 142.460 13.685 ;
        RECT 146.425 13.515 146.595 13.685 ;
        RECT 152.870 13.515 153.040 13.685 ;
        RECT 160.685 13.515 160.855 13.685 ;
        RECT 162.525 13.515 162.695 13.685 ;
        RECT 181.385 13.515 181.555 13.685 ;
        RECT 194.265 13.515 194.435 13.685 ;
        RECT 198.405 13.515 198.575 13.685 ;
        RECT 205.770 13.515 205.940 13.685 ;
        RECT 208.530 13.515 208.700 13.685 ;
        RECT 218.185 13.515 218.355 13.685 ;
        RECT 225.545 13.515 225.715 13.685 ;
        RECT 227.845 13.515 228.015 13.685 ;
        RECT 237.050 13.515 237.220 13.685 ;
        RECT 240.265 13.515 240.435 13.685 ;
        RECT 259.125 13.515 259.295 13.685 ;
        RECT 262.805 13.515 262.975 13.685 ;
        RECT 267.865 13.515 268.035 13.685 ;
        RECT 277.525 13.515 277.695 13.685 ;
        RECT 283.045 13.515 283.215 13.685 ;
        RECT 289.025 13.515 289.195 13.685 ;
        RECT 292.705 13.515 292.875 13.685 ;
        RECT 304.665 13.515 304.835 13.685 ;
        RECT 306.045 13.515 306.215 13.685 ;
        RECT 307.885 13.515 308.055 13.685 ;
        RECT 309.725 13.515 309.895 13.685 ;
        RECT 314.325 13.515 314.495 13.685 ;
        RECT 317.545 13.515 317.715 13.685 ;
        RECT 329.045 13.515 329.215 13.685 ;
        RECT 339.165 13.515 339.335 13.685 ;
        RECT 347.905 13.515 348.075 13.685 ;
        RECT 352.505 13.515 352.675 13.685 ;
        RECT 357.105 13.515 357.275 13.685 ;
        RECT 359.870 13.515 360.040 13.685 ;
        RECT 368.150 13.515 368.320 13.685 ;
        RECT 385.170 13.515 385.340 13.685 ;
        RECT 391.145 13.515 391.315 13.685 ;
        RECT 393.905 13.515 394.075 13.685 ;
        RECT 395.745 13.515 395.915 13.685 ;
        RECT 399.885 13.515 400.055 13.685 ;
        RECT 413.690 13.515 413.860 13.685 ;
        RECT 425.645 13.515 425.815 13.685 ;
        RECT 445.425 13.515 445.595 13.685 ;
        RECT 450.945 13.515 451.115 13.685 ;
        RECT 457.845 13.515 458.015 13.685 ;
        RECT 467.045 13.515 467.215 13.685 ;
        RECT 480.845 13.515 481.015 13.685 ;
        RECT 494.645 13.515 494.815 13.685 ;
        RECT 527.765 13.515 527.935 13.685 ;
        RECT 536.045 13.515 536.215 13.685 ;
        RECT 538.805 13.515 538.975 13.685 ;
        RECT 564.105 13.515 564.275 13.685 ;
        RECT 571.005 13.515 571.175 13.685 ;
        RECT 571.925 13.515 572.095 13.685 ;
        RECT 1382.445 13.515 1382.615 13.685 ;
        RECT 1400.845 13.515 1401.015 13.685 ;
        RECT 1503.885 13.515 1504.055 13.685 ;
        RECT 1525.965 13.515 1526.135 13.685 ;
        RECT 1535.625 13.515 1535.795 13.685 ;
        RECT 1539.305 13.515 1539.475 13.685 ;
        RECT 1542.525 13.515 1542.695 13.685 ;
        RECT 1559.085 13.515 1559.255 13.685 ;
        RECT 1575.645 13.515 1575.815 13.685 ;
        RECT 1588.525 13.515 1588.695 13.685 ;
        RECT 1625.785 13.515 1625.955 13.685 ;
        RECT 1648.785 13.515 1648.955 13.685 ;
        RECT 1760.105 13.515 1760.275 13.685 ;
        RECT 1773.905 13.515 1774.075 13.685 ;
        RECT 1830.025 13.515 1830.195 13.685 ;
        RECT 1913.285 13.515 1913.455 13.685 ;
        RECT 1925.705 13.515 1925.875 13.685 ;
        RECT 1931.685 13.515 1931.855 13.685 ;
        RECT 1947.785 13.515 1947.955 13.685 ;
        RECT 1973.085 13.515 1973.255 13.685 ;
        RECT 1982.745 13.515 1982.915 13.685 ;
        RECT 1991.945 13.515 1992.115 13.685 ;
        RECT 1995.165 13.515 1995.335 13.685 ;
        RECT 1999.765 13.515 1999.935 13.685 ;
        RECT 2018.165 13.515 2018.335 13.685 ;
        RECT 2024.605 13.515 2024.775 13.685 ;
        RECT 2037.485 13.515 2037.655 13.685 ;
        RECT 2059.105 13.515 2059.275 13.685 ;
        RECT 2060.485 13.515 2060.655 13.685 ;
        RECT 2073.825 13.515 2073.995 13.685 ;
        RECT 2089.925 13.515 2090.095 13.685 ;
        RECT 2105.105 13.515 2105.275 13.685 ;
        RECT 2124.885 13.515 2125.055 13.685 ;
        RECT 2135.465 13.515 2135.635 13.685 ;
        RECT 2136.845 13.515 2137.015 13.685 ;
        RECT 2140.985 13.515 2141.155 13.685 ;
        RECT 2174.105 13.515 2174.275 13.685 ;
        RECT 2179.165 13.515 2179.335 13.685 ;
        RECT 2189.745 13.515 2189.915 13.685 ;
        RECT 2192.045 13.515 2192.215 13.685 ;
        RECT 2233.905 13.515 2234.075 13.685 ;
        RECT 2238.505 13.515 2238.675 13.685 ;
        RECT 2240.805 13.515 2240.975 13.685 ;
        RECT 2271.625 13.515 2271.795 13.685 ;
        RECT 2276.685 13.515 2276.855 13.685 ;
        RECT 2296.465 13.515 2296.635 13.685 ;
        RECT 2321.305 13.515 2321.475 13.685 ;
        RECT 2427.565 13.515 2427.735 13.685 ;
        RECT 2439.525 13.515 2439.695 13.685 ;
        RECT 2490.125 13.515 2490.295 13.685 ;
        RECT 2496.105 13.515 2496.275 13.685 ;
        RECT 2497.485 13.515 2497.655 13.685 ;
        RECT 2500.245 13.515 2500.415 13.685 ;
        RECT 2501.625 13.515 2501.795 13.685 ;
        RECT 2509.445 13.515 2509.615 13.685 ;
        RECT 2525.085 13.515 2525.255 13.685 ;
        RECT 2530.145 13.515 2530.315 13.685 ;
        RECT 2533.825 13.515 2533.995 13.685 ;
        RECT 2547.625 13.515 2547.795 13.685 ;
        RECT 2551.305 13.515 2551.475 13.685 ;
        RECT 2554.065 13.515 2554.235 13.685 ;
        RECT 2569.245 13.515 2569.415 13.685 ;
        RECT 2580.745 13.515 2580.915 13.685 ;
        RECT 2585.805 13.515 2585.975 13.685 ;
        RECT 2592.705 13.515 2592.875 13.685 ;
        RECT 2597.765 13.515 2597.935 13.685 ;
        RECT 2609.265 13.515 2609.435 13.685 ;
        RECT 2655.265 13.515 2655.435 13.685 ;
        RECT 2686.085 13.515 2686.255 13.685 ;
        RECT 2688.385 13.515 2688.555 13.685 ;
        RECT 2725.645 13.515 2725.815 13.685 ;
        RECT 2727.025 13.515 2727.195 13.685 ;
        RECT 2730.245 13.515 2730.415 13.685 ;
        RECT 2855.365 13.515 2855.535 13.685 ;
        RECT 2907.345 13.515 2907.515 13.685 ;
        RECT 2908.725 13.515 2908.895 13.685 ;
        RECT 2909.185 13.515 2909.355 13.685 ;
        RECT 2910.565 13.515 2910.735 13.685 ;
        RECT 2913.785 13.515 2913.955 13.685 ;
      LAYER nwell ;
        RECT 5.330 10.690 7.090 12.295 ;
        RECT 8.550 10.690 11.690 12.295 ;
        RECT 81.690 10.690 90.810 12.295 ;
        RECT 225.210 10.690 232.030 12.295 ;
        RECT 239.930 10.690 244.450 12.295 ;
        RECT 352.170 10.690 353.930 12.295 ;
        RECT 450.610 10.690 457.430 12.295 ;
        RECT 2908.850 10.690 2910.610 12.295 ;
        RECT 2912.530 10.690 2914.290 12.295 ;
      LAYER li1 ;
        RECT 9.745 3504.340 10.265 3505.825 ;
        RECT 11.125 3504.340 11.645 3505.825 ;
        RECT 8.825 3223.455 9.345 3224.940 ;
        RECT 8.825 3011.295 9.345 3012.780 ;
        RECT 8.825 2971.220 9.345 2972.705 ;
        RECT 8.825 2954.900 9.345 2956.385 ;
        RECT 8.825 2884.180 9.345 2885.665 ;
        RECT 8.825 2869.855 9.345 2871.340 ;
        RECT 8.825 2499.935 9.345 2501.420 ;
        RECT 8.825 2380.255 9.345 2381.740 ;
        RECT 8.825 1983.135 9.345 1984.620 ;
        RECT 8.825 1953.940 9.345 1955.425 ;
        RECT 8.825 1776.415 9.345 1777.900 ;
        RECT 8.825 1705.695 9.345 1707.180 ;
        RECT 8.825 1580.575 9.345 1582.060 ;
        RECT 8.825 1328.340 9.345 1329.825 ;
        RECT 8.825 1284.820 9.345 1286.305 ;
        RECT 8.825 1273.940 9.345 1275.425 ;
        RECT 8.825 1216.095 9.345 1217.580 ;
        RECT 8.825 1110.740 9.345 1112.225 ;
        RECT 8.825 1034.580 9.345 1036.065 ;
        RECT 8.825 721.055 9.345 722.540 ;
        RECT 8.825 628.575 9.345 630.060 ;
        RECT 8.825 601.375 9.345 602.860 ;
        RECT 8.825 441.620 9.345 443.105 ;
        RECT 8.825 438.175 9.345 439.660 ;
        RECT 8.825 400.095 9.345 401.580 ;
        RECT 8.825 392.660 9.345 394.145 ;
        RECT 8.825 313.055 9.345 314.540 ;
        RECT 7.075 127.205 7.245 127.495 ;
        RECT 7.075 127.035 7.740 127.205 ;
        RECT 7.510 126.045 7.740 127.035 ;
        RECT 7.075 125.875 7.740 126.045 ;
        RECT 7.075 125.375 7.245 125.875 ;
        RECT 7.915 125.375 8.140 127.495 ;
        RECT 8.790 127.305 9.120 127.475 ;
        RECT 9.300 127.305 10.050 127.475 ;
        RECT 8.340 126.175 8.620 126.775 ;
        RECT 8.790 125.775 8.960 127.305 ;
        RECT 9.130 126.805 9.710 127.135 ;
        RECT 9.130 125.935 9.370 126.805 ;
        RECT 9.880 126.525 10.050 127.305 ;
        RECT 10.850 127.305 11.310 127.475 ;
        RECT 11.540 127.305 12.210 127.475 ;
        RECT 10.850 127.075 11.020 127.305 ;
        RECT 10.220 126.775 11.020 127.075 ;
        RECT 11.190 126.805 11.740 127.135 ;
        RECT 10.220 126.745 10.390 126.775 ;
        RECT 10.510 126.525 10.680 126.595 ;
        RECT 9.880 126.355 10.680 126.525 ;
        RECT 10.170 126.265 10.680 126.355 ;
        RECT 9.560 125.830 10.000 126.185 ;
        RECT 8.790 125.400 9.025 125.775 ;
        RECT 10.170 125.650 10.340 126.265 ;
        RECT 9.270 125.480 10.340 125.650 ;
        RECT 10.850 125.705 11.020 126.775 ;
        RECT 11.190 125.875 11.380 126.595 ;
        RECT 11.550 126.265 11.740 126.805 ;
        RECT 12.040 126.765 12.210 127.305 ;
        RECT 12.990 127.105 13.350 127.545 ;
        RECT 12.990 126.935 13.490 127.105 ;
        RECT 13.320 126.765 13.490 126.935 ;
        RECT 13.700 126.765 2906.300 3506.300 ;
        RECT 2909.125 3504.340 2909.645 3505.825 ;
        RECT 2910.505 3504.340 2911.025 3505.825 ;
        RECT 2909.125 3400.980 2909.645 3402.465 ;
        RECT 2910.505 3364.895 2911.025 3366.380 ;
        RECT 2910.505 3201.695 2911.025 3203.180 ;
        RECT 2909.125 3096.340 2909.645 3097.825 ;
        RECT 2910.505 2913.375 2911.025 2914.860 ;
        RECT 2909.125 2775.380 2909.645 2776.865 ;
        RECT 2909.125 2628.500 2909.645 2629.985 ;
        RECT 2909.125 2601.300 2909.645 2602.785 ;
        RECT 2909.125 2461.855 2909.645 2463.340 ;
        RECT 2909.125 2432.660 2909.645 2434.145 ;
        RECT 2909.125 2385.695 2909.645 2387.180 ;
        RECT 2909.125 2264.020 2909.645 2265.505 ;
        RECT 2909.125 2117.140 2909.645 2118.625 ;
        RECT 2909.125 1934.175 2909.645 1935.660 ;
        RECT 2909.125 1671.060 2909.645 1672.545 ;
        RECT 2909.125 1526.175 2909.645 1527.660 ;
        RECT 2909.125 1515.295 2909.645 1516.780 ;
        RECT 2909.125 1471.775 2909.645 1473.260 ;
        RECT 2909.125 1301.140 2909.645 1302.625 ;
        RECT 2909.125 1265.055 2909.645 1266.540 ;
        RECT 2909.125 1007.380 2909.645 1008.865 ;
        RECT 2909.125 996.500 2909.645 997.985 ;
        RECT 2909.125 811.540 2909.645 813.025 ;
        RECT 2909.125 735.380 2909.645 736.865 ;
        RECT 2909.125 468.820 2909.645 470.305 ;
        RECT 2910.505 449.055 2911.025 450.540 ;
        RECT 2909.125 289.300 2909.645 290.785 ;
        RECT 2910.505 231.455 2911.025 232.940 ;
        RECT 12.040 126.595 13.130 126.765 ;
        RECT 13.320 126.595 2906.300 126.765 ;
        RECT 11.550 125.935 11.870 126.265 ;
        RECT 10.850 125.375 11.100 125.705 ;
        RECT 12.040 125.675 12.210 126.595 ;
        RECT 13.320 126.340 13.490 126.595 ;
        RECT 12.380 126.170 13.490 126.340 ;
        RECT 12.380 126.010 13.240 126.170 ;
        RECT 11.325 125.505 12.210 125.675 ;
        RECT 13.070 125.385 13.240 126.010 ;
        RECT 9.265 105.195 9.595 105.825 ;
        RECT 10.725 105.485 10.895 109.735 ;
        RECT 8.845 104.755 9.175 105.005 ;
        RECT 9.345 104.595 9.595 105.195 ;
        RECT 9.265 103.615 9.595 104.595 ;
        RECT 7.075 42.765 7.245 43.265 ;
        RECT 7.075 42.595 7.740 42.765 ;
        RECT 7.510 41.605 7.740 42.595 ;
        RECT 7.075 41.435 7.740 41.605 ;
        RECT 7.075 41.145 7.245 41.435 ;
        RECT 7.915 41.145 8.140 43.265 ;
        RECT 8.790 42.865 9.025 43.240 ;
        RECT 9.270 42.990 10.340 43.160 ;
        RECT 8.340 41.865 8.620 42.465 ;
        RECT 8.790 41.335 8.960 42.865 ;
        RECT 9.130 41.835 9.370 42.705 ;
        RECT 9.560 42.455 10.000 42.810 ;
        RECT 10.170 42.375 10.340 42.990 ;
        RECT 10.850 42.935 11.100 43.265 ;
        RECT 11.325 42.965 12.210 43.135 ;
        RECT 10.170 42.285 10.680 42.375 ;
        RECT 9.880 42.115 10.680 42.285 ;
        RECT 9.130 41.505 9.710 41.835 ;
        RECT 9.880 41.335 10.050 42.115 ;
        RECT 10.510 42.045 10.680 42.115 ;
        RECT 10.220 41.865 10.390 41.895 ;
        RECT 10.850 41.865 11.020 42.935 ;
        RECT 11.190 42.045 11.380 42.765 ;
        RECT 11.550 42.375 11.870 42.705 ;
        RECT 10.220 41.565 11.020 41.865 ;
        RECT 11.550 41.835 11.740 42.375 ;
        RECT 8.790 41.165 9.120 41.335 ;
        RECT 9.300 41.165 10.050 41.335 ;
        RECT 10.850 41.335 11.020 41.565 ;
        RECT 11.190 41.505 11.740 41.835 ;
        RECT 12.040 42.045 12.210 42.965 ;
        RECT 13.070 42.630 13.240 43.255 ;
        RECT 12.380 42.470 13.240 42.630 ;
        RECT 12.380 42.300 13.490 42.470 ;
        RECT 13.320 42.045 13.490 42.300 ;
        RECT 13.700 42.045 2906.300 126.595 ;
        RECT 2909.125 60.820 2909.645 62.305 ;
        RECT 12.040 41.875 13.130 42.045 ;
        RECT 13.320 41.875 2906.300 42.045 ;
        RECT 12.040 41.335 12.210 41.875 ;
        RECT 13.320 41.705 13.490 41.875 ;
        RECT 10.850 41.165 11.310 41.335 ;
        RECT 11.540 41.165 12.210 41.335 ;
        RECT 12.990 41.535 13.490 41.705 ;
        RECT 12.990 41.095 13.350 41.535 ;
        RECT 7.035 20.995 7.285 21.505 ;
        RECT 7.875 20.995 8.125 21.505 ;
        RECT 8.715 21.335 9.805 21.505 ;
        RECT 8.715 20.995 8.965 21.335 ;
        RECT 9.555 21.175 9.805 21.335 ;
        RECT 10.495 21.335 11.585 21.505 ;
        RECT 10.495 21.175 10.745 21.335 ;
        RECT 7.035 20.825 8.965 20.995 ;
        RECT 8.755 20.495 8.965 20.825 ;
        RECT 9.135 21.005 9.385 21.165 ;
        RECT 10.915 21.005 11.165 21.165 ;
        RECT 9.135 20.455 9.520 21.005 ;
        RECT 10.035 20.825 11.165 21.005 ;
        RECT 11.335 20.825 11.585 21.335 ;
        RECT 12.175 20.995 12.425 21.505 ;
        RECT 13.015 20.995 13.265 21.505 ;
        RECT 12.175 20.825 13.265 20.995 ;
        RECT 10.035 20.705 10.205 20.825 ;
        RECT 9.855 20.535 10.205 20.705 ;
        RECT 13.015 20.695 13.265 20.825 ;
        RECT 13.700 20.695 2906.300 41.875 ;
        RECT 7.705 20.115 8.245 20.315 ;
        RECT 9.135 19.945 9.345 20.455 ;
        RECT 9.855 20.285 10.045 20.535 ;
        RECT 10.375 20.485 11.865 20.655 ;
        RECT 10.375 20.365 10.545 20.485 ;
        RECT 9.515 20.115 10.045 20.285 ;
        RECT 10.215 20.115 10.545 20.365 ;
        RECT 10.715 20.115 11.335 20.315 ;
        RECT 11.505 20.115 11.865 20.485 ;
        RECT 12.035 20.285 12.360 20.655 ;
        RECT 13.015 20.455 2906.300 20.695 ;
        RECT 12.035 20.115 13.340 20.285 ;
        RECT 9.855 19.945 10.045 20.115 ;
        RECT 13.510 19.945 2906.300 20.455 ;
        RECT 7.415 19.515 7.665 19.945 ;
        RECT 7.835 19.775 9.425 19.945 ;
        RECT 7.835 19.685 8.170 19.775 ;
        RECT 7.415 19.295 8.585 19.515 ;
        RECT 9.095 19.295 9.425 19.775 ;
        RECT 9.855 19.765 11.625 19.945 ;
        RECT 10.455 19.295 10.785 19.765 ;
        RECT 11.295 19.295 11.625 19.765 ;
        RECT 12.135 19.765 2906.300 19.945 ;
        RECT 12.135 19.315 12.465 19.765 ;
        RECT 12.975 19.315 13.305 19.765 ;
        RECT 7.075 18.405 7.245 18.695 ;
        RECT 7.075 18.235 7.740 18.405 ;
        RECT 7.510 17.245 7.740 18.235 ;
        RECT 7.075 17.075 7.740 17.245 ;
        RECT 7.075 16.575 7.245 17.075 ;
        RECT 7.915 16.575 8.140 18.695 ;
        RECT 8.790 18.505 9.120 18.675 ;
        RECT 9.300 18.505 10.050 18.675 ;
        RECT 8.340 17.375 8.620 17.975 ;
        RECT 8.790 16.975 8.960 18.505 ;
        RECT 9.130 18.005 9.710 18.335 ;
        RECT 9.130 17.135 9.370 18.005 ;
        RECT 9.880 17.725 10.050 18.505 ;
        RECT 10.850 18.505 11.310 18.675 ;
        RECT 11.540 18.505 12.210 18.675 ;
        RECT 10.850 18.275 11.020 18.505 ;
        RECT 10.220 17.975 11.020 18.275 ;
        RECT 11.190 18.005 11.740 18.335 ;
        RECT 10.220 17.945 10.390 17.975 ;
        RECT 10.510 17.725 10.680 17.795 ;
        RECT 9.880 17.555 10.680 17.725 ;
        RECT 10.170 17.465 10.680 17.555 ;
        RECT 9.560 17.030 10.000 17.385 ;
        RECT 8.790 16.600 9.025 16.975 ;
        RECT 10.170 16.850 10.340 17.465 ;
        RECT 9.270 16.680 10.340 16.850 ;
        RECT 10.850 16.905 11.020 17.975 ;
        RECT 11.190 17.075 11.380 17.795 ;
        RECT 11.550 17.465 11.740 18.005 ;
        RECT 12.040 17.965 12.210 18.505 ;
        RECT 12.990 18.305 13.350 18.745 ;
        RECT 12.990 18.135 13.490 18.305 ;
        RECT 13.320 17.965 13.490 18.135 ;
        RECT 13.700 17.965 2906.300 19.765 ;
        RECT 12.040 17.795 13.130 17.965 ;
        RECT 13.320 17.795 2906.300 17.965 ;
        RECT 11.550 17.135 11.870 17.465 ;
        RECT 10.850 16.575 11.100 16.905 ;
        RECT 12.040 16.875 12.210 17.795 ;
        RECT 13.320 17.540 13.490 17.795 ;
        RECT 12.380 17.370 13.490 17.540 ;
        RECT 12.380 17.210 13.240 17.370 ;
        RECT 11.325 16.705 12.210 16.875 ;
        RECT 13.070 16.585 13.240 17.210 ;
        RECT 7.075 15.565 7.245 16.065 ;
        RECT 7.075 15.395 7.740 15.565 ;
        RECT 7.510 14.405 7.740 15.395 ;
        RECT 7.075 14.235 7.740 14.405 ;
        RECT 7.075 13.945 7.245 14.235 ;
        RECT 7.915 13.945 8.140 16.065 ;
        RECT 8.790 15.665 9.025 16.040 ;
        RECT 9.270 15.790 10.340 15.960 ;
        RECT 8.340 14.665 8.620 15.265 ;
        RECT 8.790 14.135 8.960 15.665 ;
        RECT 9.130 14.635 9.370 15.505 ;
        RECT 9.560 15.255 10.000 15.610 ;
        RECT 10.170 15.175 10.340 15.790 ;
        RECT 10.850 15.735 11.100 16.065 ;
        RECT 11.325 15.765 12.210 15.935 ;
        RECT 10.170 15.085 10.680 15.175 ;
        RECT 9.880 14.915 10.680 15.085 ;
        RECT 9.130 14.305 9.710 14.635 ;
        RECT 9.880 14.135 10.050 14.915 ;
        RECT 10.510 14.845 10.680 14.915 ;
        RECT 10.220 14.665 10.390 14.695 ;
        RECT 10.850 14.665 11.020 15.735 ;
        RECT 11.190 14.845 11.380 15.565 ;
        RECT 11.550 15.175 11.870 15.505 ;
        RECT 10.220 14.365 11.020 14.665 ;
        RECT 11.550 14.635 11.740 15.175 ;
        RECT 8.790 13.965 9.120 14.135 ;
        RECT 9.300 13.965 10.050 14.135 ;
        RECT 10.850 14.135 11.020 14.365 ;
        RECT 11.190 14.305 11.740 14.635 ;
        RECT 12.040 14.845 12.210 15.765 ;
        RECT 13.070 15.430 13.240 16.055 ;
        RECT 12.380 15.270 13.240 15.430 ;
        RECT 12.380 15.100 13.490 15.270 ;
        RECT 13.320 14.845 13.490 15.100 ;
        RECT 13.700 14.845 2906.300 17.795 ;
        RECT 2909.125 17.300 2909.645 18.785 ;
        RECT 2910.505 17.300 2911.025 18.785 ;
        RECT 12.040 14.675 13.130 14.845 ;
        RECT 13.320 14.675 2906.300 14.845 ;
        RECT 12.040 14.135 12.210 14.675 ;
        RECT 13.320 14.505 13.490 14.675 ;
        RECT 10.850 13.965 11.310 14.135 ;
        RECT 11.540 13.965 12.210 14.135 ;
        RECT 12.990 14.335 13.490 14.505 ;
        RECT 12.990 13.895 13.350 14.335 ;
        RECT 13.700 13.700 2906.300 14.675 ;
        RECT 2907.285 13.855 2907.805 15.340 ;
        RECT 2908.665 13.855 2909.185 15.340 ;
        RECT 2910.505 13.855 2911.025 15.340 ;
        RECT 9.265 12.715 9.595 13.345 ;
        RECT 9.345 12.115 9.595 12.715 ;
        RECT 9.265 11.135 9.595 12.115 ;
        RECT 10.205 11.860 10.725 13.345 ;
        RECT 82.055 12.965 82.225 13.255 ;
        RECT 82.055 12.795 82.720 12.965 ;
        RECT 82.490 11.805 82.720 12.795 ;
        RECT 82.055 11.635 82.720 11.805 ;
        RECT 82.055 11.135 82.225 11.635 ;
        RECT 82.895 11.135 83.120 13.255 ;
        RECT 83.770 13.065 84.100 13.235 ;
        RECT 84.280 13.065 85.030 13.235 ;
        RECT 83.320 11.935 83.600 12.535 ;
        RECT 83.770 11.535 83.940 13.065 ;
        RECT 84.110 12.565 84.690 12.895 ;
        RECT 84.110 11.695 84.350 12.565 ;
        RECT 84.860 12.285 85.030 13.065 ;
        RECT 85.830 13.065 86.290 13.235 ;
        RECT 86.520 13.065 87.190 13.235 ;
        RECT 85.830 12.835 86.000 13.065 ;
        RECT 85.200 12.535 86.000 12.835 ;
        RECT 86.170 12.565 86.720 12.895 ;
        RECT 85.200 12.505 85.370 12.535 ;
        RECT 85.490 12.285 85.660 12.355 ;
        RECT 84.860 12.115 85.660 12.285 ;
        RECT 85.150 12.025 85.660 12.115 ;
        RECT 84.540 11.590 84.980 11.945 ;
        RECT 83.770 11.160 84.005 11.535 ;
        RECT 85.150 11.410 85.320 12.025 ;
        RECT 84.250 11.240 85.320 11.410 ;
        RECT 85.830 11.465 86.000 12.535 ;
        RECT 86.170 11.635 86.360 12.355 ;
        RECT 86.530 12.025 86.720 12.565 ;
        RECT 87.020 12.525 87.190 13.065 ;
        RECT 87.970 12.865 88.330 13.305 ;
        RECT 180.005 13.005 180.175 13.700 ;
        RECT 189.205 13.005 189.375 13.700 ;
        RECT 87.970 12.695 88.470 12.865 ;
        RECT 88.300 12.525 88.470 12.695 ;
        RECT 193.345 12.835 193.515 13.700 ;
        RECT 206.135 13.125 207.305 13.345 ;
        RECT 193.345 12.665 193.975 12.835 ;
        RECT 206.135 12.695 206.385 13.125 ;
        RECT 206.555 12.865 206.890 12.955 ;
        RECT 207.815 12.865 208.145 13.345 ;
        RECT 209.175 12.875 209.505 13.345 ;
        RECT 210.015 12.875 210.345 13.345 ;
        RECT 206.555 12.695 208.145 12.865 ;
        RECT 208.575 12.695 210.345 12.875 ;
        RECT 210.855 12.875 211.185 13.325 ;
        RECT 211.695 12.875 212.025 13.325 ;
        RECT 226.000 12.875 226.330 13.335 ;
        RECT 226.840 12.875 227.170 13.345 ;
        RECT 227.780 13.125 229.870 13.345 ;
        RECT 210.855 12.695 212.540 12.875 ;
        RECT 87.020 12.355 88.110 12.525 ;
        RECT 88.300 12.355 90.120 12.525 ;
        RECT 86.530 11.695 86.850 12.025 ;
        RECT 85.830 11.135 86.080 11.465 ;
        RECT 87.020 11.435 87.190 12.355 ;
        RECT 88.300 12.100 88.470 12.355 ;
        RECT 206.425 12.325 206.965 12.525 ;
        RECT 207.855 12.185 208.065 12.695 ;
        RECT 208.575 12.525 208.765 12.695 ;
        RECT 208.235 12.355 208.765 12.525 ;
        RECT 87.360 11.930 88.470 12.100 ;
        RECT 87.360 11.770 88.220 11.930 ;
        RECT 207.475 11.815 207.685 12.145 ;
        RECT 86.305 11.265 87.190 11.435 ;
        RECT 88.050 11.145 88.220 11.770 ;
        RECT 205.755 11.645 207.685 11.815 ;
        RECT 205.755 11.135 206.005 11.645 ;
        RECT 206.595 11.135 206.845 11.645 ;
        RECT 207.435 11.305 207.685 11.645 ;
        RECT 207.855 11.635 208.240 12.185 ;
        RECT 208.575 12.105 208.765 12.355 ;
        RECT 208.935 12.275 209.265 12.525 ;
        RECT 209.435 12.325 210.055 12.525 ;
        RECT 209.095 12.155 209.265 12.275 ;
        RECT 210.225 12.155 210.585 12.525 ;
        RECT 208.575 11.935 208.925 12.105 ;
        RECT 209.095 11.985 210.585 12.155 ;
        RECT 210.755 12.355 212.060 12.525 ;
        RECT 210.755 11.985 211.080 12.355 ;
        RECT 212.230 12.185 212.540 12.695 ;
        RECT 208.755 11.815 208.925 11.935 ;
        RECT 211.735 11.945 212.540 12.185 ;
        RECT 225.485 12.695 227.170 12.875 ;
        RECT 227.815 12.865 229.370 12.955 ;
        RECT 227.340 12.695 229.370 12.865 ;
        RECT 229.540 12.865 229.870 13.125 ;
        RECT 230.380 12.875 230.710 13.345 ;
        RECT 231.220 12.875 231.550 13.345 ;
        RECT 230.380 12.865 231.550 12.875 ;
        RECT 229.540 12.695 231.550 12.865 ;
        RECT 240.585 13.225 240.920 13.345 ;
        RECT 240.585 13.035 241.845 13.225 ;
        RECT 240.585 12.795 240.920 13.035 ;
        RECT 241.655 12.985 241.845 13.035 ;
        RECT 242.570 12.985 242.760 13.085 ;
        RECT 243.430 12.985 243.620 13.345 ;
        RECT 255.445 13.005 256.075 13.175 ;
        RECT 241.655 12.795 242.400 12.985 ;
        RECT 225.485 12.155 225.770 12.695 ;
        RECT 227.340 12.525 227.630 12.695 ;
        RECT 225.940 12.325 227.630 12.525 ;
        RECT 225.485 11.985 227.130 12.155 ;
        RECT 211.735 11.815 211.985 11.945 ;
        RECT 208.755 11.635 209.885 11.815 ;
        RECT 207.855 11.475 208.105 11.635 ;
        RECT 209.635 11.475 209.885 11.635 ;
        RECT 208.275 11.305 208.525 11.465 ;
        RECT 207.435 11.135 208.525 11.305 ;
        RECT 209.215 11.305 209.465 11.465 ;
        RECT 210.055 11.305 210.305 11.815 ;
        RECT 209.215 11.135 210.305 11.305 ;
        RECT 210.895 11.645 211.985 11.815 ;
        RECT 210.895 11.135 211.145 11.645 ;
        RECT 211.735 11.135 211.985 11.645 ;
        RECT 213.585 7.905 213.755 11.475 ;
        RECT 226.040 11.135 226.290 11.985 ;
        RECT 226.880 11.135 227.130 11.985 ;
        RECT 227.300 11.815 227.630 12.325 ;
        RECT 227.820 12.155 228.355 12.525 ;
        RECT 228.525 12.325 229.080 12.525 ;
        RECT 229.250 12.155 229.580 12.525 ;
        RECT 227.820 11.985 229.580 12.155 ;
        RECT 229.750 12.155 230.080 12.525 ;
        RECT 230.965 12.325 231.755 12.525 ;
        RECT 230.965 12.155 231.135 12.325 ;
        RECT 229.750 11.985 231.135 12.155 ;
        RECT 240.235 12.260 240.995 12.605 ;
        RECT 242.190 12.580 242.400 12.795 ;
        RECT 242.570 12.755 244.175 12.985 ;
        RECT 227.300 11.645 230.670 11.815 ;
        RECT 228.660 11.475 228.910 11.645 ;
        RECT 230.420 11.475 230.670 11.645 ;
        RECT 228.240 11.305 228.490 11.475 ;
        RECT 229.080 11.305 229.330 11.475 ;
        RECT 228.240 11.135 229.330 11.305 ;
        RECT 230.000 11.305 230.250 11.475 ;
        RECT 230.840 11.305 231.090 11.815 ;
        RECT 230.000 11.135 231.090 11.305 ;
        RECT 240.235 11.265 240.485 12.260 ;
        RECT 242.190 12.245 243.725 12.580 ;
        RECT 242.190 12.020 242.400 12.245 ;
        RECT 243.895 12.065 244.175 12.755 ;
        RECT 255.905 12.665 256.075 13.005 ;
        RECT 263.260 12.875 263.590 13.335 ;
        RECT 264.100 12.875 264.430 13.345 ;
        RECT 265.040 13.125 267.130 13.345 ;
        RECT 262.745 12.695 264.430 12.875 ;
        RECT 265.075 12.865 266.630 12.955 ;
        RECT 264.600 12.695 266.630 12.865 ;
        RECT 266.800 12.865 267.130 13.125 ;
        RECT 267.640 12.875 267.970 13.345 ;
        RECT 268.480 12.875 268.810 13.345 ;
        RECT 267.640 12.865 268.810 12.875 ;
        RECT 266.800 12.695 268.810 12.865 ;
        RECT 240.665 11.850 242.400 12.020 ;
        RECT 240.665 11.135 240.845 11.850 ;
        RECT 241.640 11.135 241.820 11.850 ;
        RECT 242.570 11.840 244.175 12.065 ;
        RECT 242.570 11.135 242.760 11.840 ;
        RECT 243.430 11.835 244.175 11.840 ;
        RECT 243.430 11.135 243.620 11.835 ;
        RECT 255.445 7.565 255.615 12.495 ;
        RECT 262.745 12.155 263.030 12.695 ;
        RECT 264.600 12.525 264.890 12.695 ;
        RECT 263.200 12.325 264.890 12.525 ;
        RECT 262.745 11.985 264.390 12.155 ;
        RECT 263.300 11.135 263.550 11.985 ;
        RECT 264.140 11.135 264.390 11.985 ;
        RECT 264.560 11.815 264.890 12.325 ;
        RECT 265.080 12.155 265.615 12.525 ;
        RECT 265.785 12.325 266.340 12.525 ;
        RECT 266.510 12.155 266.840 12.525 ;
        RECT 265.080 11.985 266.840 12.155 ;
        RECT 267.010 12.155 267.340 12.525 ;
        RECT 268.225 12.325 269.015 12.525 ;
        RECT 268.225 12.155 268.395 12.325 ;
        RECT 267.010 11.985 268.395 12.155 ;
        RECT 264.560 11.645 267.930 11.815 ;
        RECT 265.920 11.475 266.170 11.645 ;
        RECT 267.680 11.475 267.930 11.645 ;
        RECT 265.500 11.305 265.750 11.475 ;
        RECT 266.340 11.305 266.590 11.475 ;
        RECT 265.500 11.135 266.590 11.305 ;
        RECT 267.260 11.305 267.510 11.475 ;
        RECT 268.100 11.305 268.350 11.815 ;
        RECT 267.260 11.135 268.350 11.305 ;
        RECT 269.245 7.225 269.415 8.755 ;
        RECT 269.705 7.565 269.875 12.155 ;
        RECT 270.165 11.985 270.335 13.700 ;
        RECT 279.365 11.645 279.535 12.835 ;
        RECT 285.345 11.985 285.515 13.700 ;
        RECT 291.785 12.325 291.955 13.700 ;
        RECT 306.505 9.265 306.675 12.155 ;
        RECT 327.665 11.645 327.835 12.835 ;
        RECT 352.885 12.715 353.215 13.345 ;
        RECT 352.465 12.275 352.795 12.525 ;
        RECT 352.965 12.115 353.215 12.715 ;
        RECT 352.885 11.135 353.215 12.115 ;
        RECT 375.505 9.945 375.675 13.175 ;
        RECT 391.175 12.965 391.345 13.255 ;
        RECT 391.175 12.795 391.840 12.965 ;
        RECT 391.610 11.805 391.840 12.795 ;
        RECT 391.175 11.635 391.840 11.805 ;
        RECT 391.175 11.135 391.345 11.635 ;
        RECT 392.015 11.135 392.240 13.255 ;
        RECT 392.890 13.065 393.220 13.235 ;
        RECT 393.400 13.065 394.150 13.235 ;
        RECT 392.440 11.935 392.720 12.535 ;
        RECT 392.890 11.535 393.060 13.065 ;
        RECT 393.230 12.565 393.810 12.895 ;
        RECT 393.230 11.695 393.470 12.565 ;
        RECT 393.980 12.285 394.150 13.065 ;
        RECT 394.950 13.065 395.410 13.235 ;
        RECT 395.640 13.065 396.310 13.235 ;
        RECT 394.950 12.835 395.120 13.065 ;
        RECT 394.320 12.535 395.120 12.835 ;
        RECT 395.290 12.565 395.840 12.895 ;
        RECT 394.320 12.505 394.490 12.535 ;
        RECT 394.610 12.285 394.780 12.355 ;
        RECT 393.980 12.115 394.780 12.285 ;
        RECT 394.270 12.025 394.780 12.115 ;
        RECT 393.660 11.590 394.100 11.945 ;
        RECT 392.890 11.160 393.125 11.535 ;
        RECT 394.270 11.410 394.440 12.025 ;
        RECT 393.370 11.240 394.440 11.410 ;
        RECT 394.950 11.465 395.120 12.535 ;
        RECT 395.290 11.635 395.480 12.355 ;
        RECT 395.650 12.025 395.840 12.565 ;
        RECT 396.140 12.525 396.310 13.065 ;
        RECT 397.090 12.865 397.450 13.305 ;
        RECT 397.090 12.695 397.590 12.865 ;
        RECT 400.265 12.715 400.595 13.345 ;
        RECT 451.400 12.875 451.730 13.335 ;
        RECT 452.240 12.875 452.570 13.345 ;
        RECT 453.180 13.125 455.270 13.345 ;
        RECT 397.420 12.525 397.590 12.695 ;
        RECT 396.140 12.355 397.230 12.525 ;
        RECT 397.420 12.355 399.240 12.525 ;
        RECT 395.650 11.695 395.970 12.025 ;
        RECT 394.950 11.135 395.200 11.465 ;
        RECT 396.140 11.435 396.310 12.355 ;
        RECT 397.420 12.100 397.590 12.355 ;
        RECT 399.845 12.275 400.175 12.525 ;
        RECT 400.345 12.115 400.595 12.715 ;
        RECT 450.885 12.695 452.570 12.875 ;
        RECT 453.215 12.865 454.770 12.955 ;
        RECT 452.740 12.695 454.770 12.865 ;
        RECT 454.940 12.865 455.270 13.125 ;
        RECT 455.780 12.875 456.110 13.345 ;
        RECT 456.620 12.875 456.950 13.345 ;
        RECT 455.780 12.865 456.950 12.875 ;
        RECT 454.940 12.695 456.950 12.865 ;
        RECT 396.480 11.930 397.590 12.100 ;
        RECT 396.480 11.770 397.340 11.930 ;
        RECT 395.425 11.265 396.310 11.435 ;
        RECT 397.170 11.145 397.340 11.770 ;
        RECT 400.265 11.135 400.595 12.115 ;
        RECT 450.025 9.265 450.195 12.495 ;
        RECT 450.885 12.155 451.170 12.695 ;
        RECT 452.740 12.525 453.030 12.695 ;
        RECT 451.340 12.325 453.030 12.525 ;
        RECT 450.885 11.985 452.530 12.155 ;
        RECT 451.440 11.135 451.690 11.985 ;
        RECT 452.280 11.135 452.530 11.985 ;
        RECT 452.700 11.815 453.030 12.325 ;
        RECT 453.220 12.155 453.755 12.525 ;
        RECT 453.925 12.325 454.480 12.525 ;
        RECT 454.650 12.155 454.980 12.525 ;
        RECT 453.220 11.985 454.980 12.155 ;
        RECT 455.150 12.155 455.480 12.525 ;
        RECT 456.365 12.325 457.155 12.525 ;
        RECT 456.365 12.155 456.535 12.325 ;
        RECT 455.150 11.985 456.535 12.155 ;
        RECT 2909.125 11.860 2909.645 13.345 ;
        RECT 452.700 11.645 456.070 11.815 ;
        RECT 454.060 11.475 454.310 11.645 ;
        RECT 455.820 11.475 456.070 11.645 ;
        RECT 453.640 11.305 453.890 11.475 ;
        RECT 454.480 11.305 454.730 11.475 ;
        RECT 453.640 11.135 454.730 11.305 ;
        RECT 455.400 11.305 455.650 11.475 ;
        RECT 456.240 11.305 456.490 11.815 ;
        RECT 455.400 11.135 456.490 11.305 ;
      LAYER mcon ;
        RECT 9.345 13.005 9.515 13.175 ;
        RECT 82.490 11.645 82.660 11.815 ;
        RECT 82.950 12.665 83.120 12.835 ;
        RECT 83.405 11.985 83.575 12.155 ;
        RECT 84.350 12.665 84.520 12.835 ;
        RECT 86.190 12.665 86.360 12.835 ;
        RECT 84.810 11.645 84.980 11.815 ;
        RECT 86.190 11.645 86.360 11.815 ;
        RECT 193.805 12.665 193.975 12.835 ;
        RECT 226.005 13.005 226.175 13.175 ;
        RECT 206.685 12.325 206.855 12.495 ;
        RECT 208.070 11.985 208.240 12.155 ;
        RECT 209.445 12.325 209.615 12.495 ;
        RECT 210.365 12.325 210.535 12.495 ;
        RECT 210.850 11.985 211.020 12.155 ;
        RECT 211.745 11.305 211.915 11.475 ;
        RECT 213.585 11.305 213.755 11.475 ;
        RECT 228.765 12.325 228.935 12.495 ;
        RECT 228.305 11.985 228.475 12.155 ;
        RECT 231.525 12.325 231.695 12.495 ;
        RECT 240.265 12.325 240.435 12.495 ;
        RECT 263.265 13.005 263.435 13.175 ;
        RECT 243.945 11.985 244.115 12.155 ;
        RECT 255.445 12.325 255.615 12.495 ;
        RECT 266.025 12.325 266.195 12.495 ;
        RECT 266.485 11.985 266.655 12.155 ;
        RECT 267.405 11.985 267.575 12.155 ;
        RECT 269.705 11.985 269.875 12.155 ;
        RECT 279.365 12.665 279.535 12.835 ;
        RECT 327.665 12.665 327.835 12.835 ;
        RECT 306.505 11.985 306.675 12.155 ;
        RECT 352.965 12.665 353.135 12.835 ;
        RECT 352.505 12.325 352.675 12.495 ;
        RECT 375.505 13.005 375.675 13.175 ;
        RECT 391.610 11.645 391.780 11.815 ;
        RECT 392.070 12.665 392.240 12.835 ;
        RECT 392.525 12.325 392.695 12.495 ;
        RECT 393.470 12.665 393.640 12.835 ;
        RECT 395.310 12.665 395.480 12.835 ;
        RECT 393.930 11.645 394.100 11.815 ;
        RECT 395.310 11.645 395.480 11.815 ;
        RECT 451.405 13.005 451.575 13.175 ;
        RECT 399.885 12.325 400.055 12.495 ;
        RECT 400.345 11.645 400.515 11.815 ;
        RECT 450.025 12.325 450.195 12.495 ;
        RECT 454.165 12.325 454.335 12.495 ;
        RECT 454.625 11.985 454.795 12.155 ;
        RECT 456.925 12.325 457.095 12.495 ;
        RECT 269.245 8.585 269.415 8.755 ;
        RECT 269.705 8.585 269.875 8.755 ;
        RECT 7.510 125.885 7.680 126.055 ;
        RECT 7.970 126.905 8.140 127.075 ;
        RECT 8.425 126.225 8.595 126.395 ;
        RECT 9.370 126.905 9.540 127.075 ;
        RECT 11.210 126.905 11.380 127.075 ;
        RECT 9.830 125.885 10.000 126.055 ;
        RECT 11.210 125.885 11.380 126.055 ;
        RECT 10.725 109.565 10.895 109.735 ;
        RECT 9.345 105.485 9.515 105.655 ;
        RECT 8.845 104.805 9.015 104.975 ;
        RECT 7.510 42.585 7.680 42.755 ;
        RECT 8.425 42.245 8.595 42.415 ;
        RECT 7.970 41.565 8.140 41.735 ;
        RECT 9.830 42.585 10.000 42.755 ;
        RECT 9.370 41.565 9.540 41.735 ;
        RECT 11.210 42.585 11.380 42.755 ;
        RECT 11.210 41.565 11.380 41.735 ;
        RECT 9.350 20.485 9.520 20.655 ;
        RECT 7.965 20.145 8.135 20.315 ;
        RECT 10.725 20.145 10.895 20.315 ;
        RECT 11.645 20.145 11.815 20.315 ;
        RECT 12.130 20.485 12.300 20.655 ;
        RECT 13.485 20.485 13.655 20.655 ;
        RECT 7.510 17.085 7.680 17.255 ;
        RECT 7.970 18.105 8.140 18.275 ;
        RECT 8.425 17.765 8.595 17.935 ;
        RECT 9.370 18.105 9.540 18.275 ;
        RECT 11.210 18.105 11.380 18.275 ;
        RECT 9.830 17.085 10.000 17.255 ;
        RECT 11.210 17.085 11.380 17.255 ;
        RECT 7.510 15.385 7.680 15.555 ;
        RECT 8.425 14.705 8.595 14.875 ;
        RECT 7.970 14.365 8.140 14.535 ;
        RECT 9.830 15.385 10.000 15.555 ;
        RECT 9.370 14.365 9.540 14.535 ;
        RECT 11.210 15.385 11.380 15.555 ;
        RECT 11.210 14.365 11.380 14.535 ;
      LAYER met1 ;
        RECT 9.730 155.960 10.050 156.020 ;
        RECT 13.700 155.960 2906.300 3506.300 ;
        RECT 9.730 155.820 2906.300 155.960 ;
        RECT 9.730 155.760 10.050 155.820 ;
        RECT 8.810 152.900 9.130 152.960 ;
        RECT 13.700 152.900 2906.300 155.820 ;
        RECT 8.810 152.760 2906.300 152.900 ;
        RECT 8.810 152.700 9.130 152.760 ;
        RECT 7.910 127.060 8.200 127.105 ;
        RECT 9.310 127.060 9.600 127.105 ;
        RECT 11.150 127.060 11.440 127.105 ;
        RECT 7.910 126.920 11.440 127.060 ;
        RECT 7.910 126.875 8.200 126.920 ;
        RECT 9.310 126.875 9.600 126.920 ;
        RECT 11.150 126.875 11.440 126.920 ;
        RECT 8.350 126.380 8.670 126.440 ;
        RECT 8.155 126.240 8.670 126.380 ;
        RECT 8.350 126.180 8.670 126.240 ;
        RECT 7.450 126.040 7.740 126.085 ;
        RECT 9.770 126.040 10.060 126.085 ;
        RECT 11.150 126.040 11.440 126.085 ;
        RECT 7.450 125.900 11.440 126.040 ;
        RECT 7.450 125.855 7.740 125.900 ;
        RECT 9.770 125.855 10.060 125.900 ;
        RECT 11.150 125.855 11.440 125.900 ;
        RECT 10.665 109.720 10.955 109.765 ;
        RECT 13.700 109.720 2906.300 152.760 ;
        RECT 10.665 109.580 2906.300 109.720 ;
        RECT 10.665 109.535 10.955 109.580 ;
        RECT 9.285 105.640 9.575 105.685 ;
        RECT 10.665 105.640 10.955 105.685 ;
        RECT 9.285 105.500 10.955 105.640 ;
        RECT 9.285 105.455 9.575 105.500 ;
        RECT 10.665 105.455 10.955 105.500 ;
        RECT 8.785 104.775 9.075 105.005 ;
        RECT 8.900 104.620 9.040 104.775 ;
        RECT 13.700 104.620 2906.300 109.580 ;
        RECT 8.900 104.480 2906.300 104.620 ;
        RECT 8.350 90.340 8.670 90.400 ;
        RECT 13.700 90.340 2906.300 104.480 ;
        RECT 8.350 90.200 2906.300 90.340 ;
        RECT 8.350 90.140 8.670 90.200 ;
        RECT 7.450 42.740 7.740 42.785 ;
        RECT 9.770 42.740 10.060 42.785 ;
        RECT 11.150 42.740 11.440 42.785 ;
        RECT 7.450 42.600 11.440 42.740 ;
        RECT 7.450 42.555 7.740 42.600 ;
        RECT 9.770 42.555 10.060 42.600 ;
        RECT 11.150 42.555 11.440 42.600 ;
        RECT 8.365 42.400 8.655 42.445 ;
        RECT 13.700 42.400 2906.300 90.200 ;
        RECT 8.365 42.260 2906.300 42.400 ;
        RECT 8.365 42.215 8.655 42.260 ;
        RECT 7.910 41.720 8.200 41.765 ;
        RECT 9.310 41.720 9.600 41.765 ;
        RECT 11.150 41.720 11.440 41.765 ;
        RECT 7.910 41.580 11.440 41.720 ;
        RECT 7.910 41.535 8.200 41.580 ;
        RECT 9.310 41.535 9.600 41.580 ;
        RECT 11.150 41.535 11.440 41.580 ;
        RECT 13.700 24.100 2906.300 42.260 ;
        RECT 13.410 23.840 2906.300 24.100 ;
        RECT 13.700 20.700 2906.300 23.840 ;
        RECT 9.290 20.640 9.580 20.685 ;
        RECT 12.070 20.640 12.360 20.685 ;
        RECT 13.410 20.640 2906.300 20.700 ;
        RECT 7.980 20.500 9.040 20.640 ;
        RECT 7.980 20.345 8.120 20.500 ;
        RECT 7.905 20.115 8.195 20.345 ;
        RECT 8.900 20.300 9.040 20.500 ;
        RECT 9.290 20.500 12.360 20.640 ;
        RECT 13.215 20.500 2906.300 20.640 ;
        RECT 9.290 20.455 9.580 20.500 ;
        RECT 12.070 20.455 12.360 20.500 ;
        RECT 13.410 20.440 2906.300 20.500 ;
        RECT 10.650 20.300 10.970 20.360 ;
        RECT 11.570 20.300 11.890 20.360 ;
        RECT 8.900 20.160 10.970 20.300 ;
        RECT 11.375 20.160 11.890 20.300 ;
        RECT 10.650 20.100 10.970 20.160 ;
        RECT 11.570 20.100 11.890 20.160 ;
        RECT 10.190 18.600 10.510 18.660 ;
        RECT 13.700 18.600 2906.300 20.440 ;
        RECT 10.190 18.460 2906.300 18.600 ;
        RECT 10.190 18.400 10.510 18.460 ;
        RECT 7.910 18.260 8.200 18.305 ;
        RECT 9.310 18.260 9.600 18.305 ;
        RECT 11.150 18.260 11.440 18.305 ;
        RECT 7.910 18.120 11.440 18.260 ;
        RECT 7.910 18.075 8.200 18.120 ;
        RECT 9.310 18.075 9.600 18.120 ;
        RECT 11.150 18.075 11.440 18.120 ;
        RECT 8.365 17.920 8.655 17.965 ;
        RECT 8.810 17.920 9.130 17.980 ;
        RECT 8.365 17.780 9.130 17.920 ;
        RECT 8.365 17.735 8.655 17.780 ;
        RECT 8.810 17.720 9.130 17.780 ;
        RECT 10.650 17.580 10.970 17.640 ;
        RECT 13.700 17.580 2906.300 18.460 ;
        RECT 10.650 17.440 2906.300 17.580 ;
        RECT 10.650 17.380 10.970 17.440 ;
        RECT 7.450 17.240 7.740 17.285 ;
        RECT 9.770 17.240 10.060 17.285 ;
        RECT 11.150 17.240 11.440 17.285 ;
        RECT 7.450 17.100 11.440 17.240 ;
        RECT 7.450 17.055 7.740 17.100 ;
        RECT 9.770 17.055 10.060 17.100 ;
        RECT 11.150 17.055 11.440 17.100 ;
        RECT 7.450 15.540 7.740 15.585 ;
        RECT 9.770 15.540 10.060 15.585 ;
        RECT 11.150 15.540 11.440 15.585 ;
        RECT 7.450 15.400 11.440 15.540 ;
        RECT 7.450 15.355 7.740 15.400 ;
        RECT 9.770 15.355 10.060 15.400 ;
        RECT 11.150 15.355 11.440 15.400 ;
        RECT 8.365 14.860 8.655 14.905 ;
        RECT 9.730 14.860 10.050 14.920 ;
        RECT 8.365 14.720 10.050 14.860 ;
        RECT 8.365 14.675 8.655 14.720 ;
        RECT 9.730 14.660 10.050 14.720 ;
        RECT 7.910 14.520 8.200 14.565 ;
        RECT 9.310 14.520 9.600 14.565 ;
        RECT 11.150 14.520 11.440 14.565 ;
        RECT 7.910 14.380 11.440 14.520 ;
        RECT 7.910 14.335 8.200 14.380 ;
        RECT 9.310 14.335 9.600 14.380 ;
        RECT 11.150 14.335 11.440 14.380 ;
        RECT 13.700 13.700 2906.300 17.440 ;
        RECT 9.285 13.160 9.575 13.205 ;
        RECT 10.190 13.160 10.510 13.220 ;
        RECT 9.285 13.020 10.510 13.160 ;
        RECT 9.285 12.975 9.575 13.020 ;
        RECT 10.190 12.960 10.510 13.020 ;
        RECT 179.945 13.160 180.235 13.205 ;
        RECT 189.145 13.160 189.435 13.205 ;
        RECT 225.930 13.160 226.250 13.220 ;
        RECT 255.385 13.160 255.675 13.205 ;
        RECT 263.190 13.160 263.510 13.220 ;
        RECT 268.250 13.160 268.570 13.220 ;
        RECT 375.445 13.160 375.735 13.205 ;
        RECT 179.945 13.020 189.435 13.160 ;
        RECT 225.735 13.020 226.250 13.160 ;
        RECT 179.945 12.975 180.235 13.020 ;
        RECT 189.145 12.975 189.435 13.020 ;
        RECT 225.930 12.960 226.250 13.020 ;
        RECT 226.480 13.020 255.675 13.160 ;
        RECT 262.995 13.020 263.510 13.160 ;
        RECT 82.890 12.820 83.180 12.865 ;
        RECT 84.290 12.820 84.580 12.865 ;
        RECT 86.130 12.820 86.420 12.865 ;
        RECT 82.890 12.680 86.420 12.820 ;
        RECT 82.890 12.635 83.180 12.680 ;
        RECT 84.290 12.635 84.580 12.680 ;
        RECT 86.130 12.635 86.420 12.680 ;
        RECT 193.745 12.820 194.035 12.865 ;
        RECT 197.870 12.820 198.190 12.880 ;
        RECT 193.745 12.680 198.190 12.820 ;
        RECT 193.745 12.635 194.035 12.680 ;
        RECT 197.870 12.620 198.190 12.680 ;
        RECT 210.750 12.620 211.070 12.880 ;
        RECT 156.010 12.480 156.330 12.540 ;
        RECT 167.510 12.480 167.830 12.540 ;
        RECT 156.010 12.340 167.830 12.480 ;
        RECT 156.010 12.280 156.330 12.340 ;
        RECT 167.510 12.280 167.830 12.340 ;
        RECT 184.530 12.480 184.850 12.540 ;
        RECT 193.270 12.480 193.590 12.540 ;
        RECT 199.250 12.480 199.570 12.540 ;
        RECT 184.530 12.340 199.570 12.480 ;
        RECT 184.530 12.280 184.850 12.340 ;
        RECT 193.270 12.280 193.590 12.340 ;
        RECT 199.250 12.280 199.570 12.340 ;
        RECT 206.625 12.480 206.915 12.525 ;
        RECT 207.070 12.480 207.390 12.540 ;
        RECT 209.385 12.480 209.675 12.525 ;
        RECT 210.290 12.480 210.610 12.540 ;
        RECT 206.625 12.340 209.675 12.480 ;
        RECT 210.095 12.340 210.610 12.480 ;
        RECT 210.840 12.480 210.980 12.620 ;
        RECT 226.480 12.480 226.620 13.020 ;
        RECT 255.385 12.975 255.675 13.020 ;
        RECT 263.190 12.960 263.510 13.020 ;
        RECT 263.740 13.020 268.020 13.160 ;
        RECT 255.845 12.820 256.135 12.865 ;
        RECT 263.740 12.820 263.880 13.020 ;
        RECT 231.540 12.680 255.600 12.820 ;
        RECT 228.690 12.480 229.010 12.540 ;
        RECT 231.540 12.525 231.680 12.680 ;
        RECT 210.840 12.340 226.620 12.480 ;
        RECT 228.495 12.340 229.010 12.480 ;
        RECT 206.625 12.295 206.915 12.340 ;
        RECT 207.070 12.280 207.390 12.340 ;
        RECT 209.385 12.295 209.675 12.340 ;
        RECT 210.290 12.280 210.610 12.340 ;
        RECT 228.690 12.280 229.010 12.340 ;
        RECT 231.465 12.295 231.755 12.525 ;
        RECT 238.810 12.480 239.130 12.540 ;
        RECT 255.460 12.525 255.600 12.680 ;
        RECT 255.845 12.680 263.880 12.820 ;
        RECT 267.880 12.820 268.020 13.020 ;
        RECT 268.250 13.020 375.735 13.160 ;
        RECT 268.250 12.960 268.570 13.020 ;
        RECT 375.445 12.975 375.735 13.020 ;
        RECT 396.130 13.160 396.450 13.220 ;
        RECT 400.270 13.160 400.590 13.220 ;
        RECT 451.330 13.160 451.650 13.220 ;
        RECT 396.130 13.020 400.590 13.160 ;
        RECT 451.135 13.020 451.650 13.160 ;
        RECT 396.130 12.960 396.450 13.020 ;
        RECT 400.270 12.960 400.590 13.020 ;
        RECT 451.330 12.960 451.650 13.020 ;
        RECT 279.305 12.820 279.595 12.865 ;
        RECT 267.880 12.680 279.595 12.820 ;
        RECT 255.845 12.635 256.135 12.680 ;
        RECT 279.305 12.635 279.595 12.680 ;
        RECT 298.610 12.820 298.930 12.880 ;
        RECT 309.650 12.820 309.970 12.880 ;
        RECT 298.610 12.680 309.970 12.820 ;
        RECT 298.610 12.620 298.930 12.680 ;
        RECT 309.650 12.620 309.970 12.680 ;
        RECT 327.605 12.820 327.895 12.865 ;
        RECT 352.905 12.820 353.195 12.865 ;
        RECT 327.605 12.680 353.195 12.820 ;
        RECT 327.605 12.635 327.895 12.680 ;
        RECT 352.905 12.635 353.195 12.680 ;
        RECT 392.010 12.820 392.300 12.865 ;
        RECT 393.410 12.820 393.700 12.865 ;
        RECT 395.250 12.820 395.540 12.865 ;
        RECT 529.990 12.820 530.310 12.880 ;
        RECT 392.010 12.680 395.540 12.820 ;
        RECT 392.010 12.635 392.300 12.680 ;
        RECT 393.410 12.635 393.700 12.680 ;
        RECT 395.250 12.635 395.540 12.680 ;
        RECT 454.640 12.680 530.310 12.820 ;
        RECT 240.205 12.480 240.495 12.525 ;
        RECT 238.810 12.340 240.495 12.480 ;
        RECT 238.810 12.280 239.130 12.340 ;
        RECT 240.205 12.295 240.495 12.340 ;
        RECT 255.385 12.295 255.675 12.525 ;
        RECT 265.490 12.480 265.810 12.540 ;
        RECT 265.965 12.480 266.255 12.525 ;
        RECT 265.490 12.340 266.255 12.480 ;
        RECT 265.490 12.280 265.810 12.340 ;
        RECT 265.965 12.295 266.255 12.340 ;
        RECT 291.725 12.480 292.015 12.525 ;
        RECT 326.670 12.480 326.990 12.540 ;
        RECT 291.725 12.340 326.990 12.480 ;
        RECT 291.725 12.295 292.015 12.340 ;
        RECT 326.670 12.280 326.990 12.340 ;
        RECT 352.445 12.480 352.735 12.525 ;
        RECT 353.810 12.480 354.130 12.540 ;
        RECT 392.450 12.480 392.770 12.540 ;
        RECT 399.810 12.480 400.130 12.540 ;
        RECT 352.445 12.340 354.130 12.480 ;
        RECT 392.255 12.340 392.770 12.480 ;
        RECT 399.615 12.340 400.130 12.480 ;
        RECT 352.445 12.295 352.735 12.340 ;
        RECT 353.810 12.280 354.130 12.340 ;
        RECT 392.450 12.280 392.770 12.340 ;
        RECT 399.810 12.280 400.130 12.340 ;
        RECT 400.270 12.480 400.590 12.540 ;
        RECT 449.965 12.480 450.255 12.525 ;
        RECT 454.105 12.480 454.395 12.525 ;
        RECT 400.270 12.340 401.420 12.480 ;
        RECT 400.270 12.280 400.590 12.340 ;
        RECT 83.345 12.140 83.635 12.185 ;
        RECT 145.890 12.140 146.210 12.200 ;
        RECT 83.345 12.000 146.210 12.140 ;
        RECT 83.345 11.955 83.635 12.000 ;
        RECT 145.890 11.940 146.210 12.000 ;
        RECT 208.010 12.140 208.300 12.185 ;
        RECT 210.790 12.140 211.080 12.185 ;
        RECT 228.230 12.140 228.550 12.200 ;
        RECT 208.010 12.000 211.080 12.140 ;
        RECT 228.035 12.000 228.550 12.140 ;
        RECT 208.010 11.955 208.300 12.000 ;
        RECT 210.790 11.955 211.080 12.000 ;
        RECT 228.230 11.940 228.550 12.000 ;
        RECT 242.490 12.140 242.810 12.200 ;
        RECT 243.885 12.140 244.175 12.185 ;
        RECT 242.490 12.000 244.175 12.140 ;
        RECT 242.490 11.940 242.810 12.000 ;
        RECT 243.885 11.955 244.175 12.000 ;
        RECT 266.425 12.140 266.715 12.185 ;
        RECT 266.870 12.140 267.190 12.200 ;
        RECT 266.425 12.000 267.190 12.140 ;
        RECT 266.425 11.955 266.715 12.000 ;
        RECT 266.870 11.940 267.190 12.000 ;
        RECT 267.345 12.140 267.635 12.185 ;
        RECT 269.645 12.140 269.935 12.185 ;
        RECT 267.345 12.000 269.935 12.140 ;
        RECT 267.345 11.955 267.635 12.000 ;
        RECT 269.645 11.955 269.935 12.000 ;
        RECT 270.105 12.140 270.395 12.185 ;
        RECT 285.285 12.140 285.575 12.185 ;
        RECT 270.105 12.000 285.575 12.140 ;
        RECT 270.105 11.955 270.395 12.000 ;
        RECT 285.285 11.955 285.575 12.000 ;
        RECT 304.590 12.140 304.910 12.200 ;
        RECT 306.445 12.140 306.735 12.185 ;
        RECT 304.590 12.000 306.735 12.140 ;
        RECT 401.280 12.140 401.420 12.340 ;
        RECT 449.965 12.340 454.395 12.480 ;
        RECT 449.965 12.295 450.255 12.340 ;
        RECT 454.105 12.295 454.395 12.340 ;
        RECT 454.640 12.185 454.780 12.680 ;
        RECT 529.990 12.620 530.310 12.680 ;
        RECT 456.865 12.480 457.155 12.525 ;
        RECT 457.770 12.480 458.090 12.540 ;
        RECT 456.865 12.340 458.090 12.480 ;
        RECT 456.865 12.295 457.155 12.340 ;
        RECT 457.770 12.280 458.090 12.340 ;
        RECT 454.565 12.140 454.855 12.185 ;
        RECT 401.280 12.000 454.855 12.140 ;
        RECT 304.590 11.940 304.910 12.000 ;
        RECT 306.445 11.955 306.735 12.000 ;
        RECT 454.565 11.955 454.855 12.000 ;
        RECT 82.430 11.800 82.720 11.845 ;
        RECT 84.750 11.800 85.040 11.845 ;
        RECT 86.130 11.800 86.420 11.845 ;
        RECT 82.430 11.660 86.420 11.800 ;
        RECT 82.430 11.615 82.720 11.660 ;
        RECT 84.750 11.615 85.040 11.660 ;
        RECT 86.130 11.615 86.420 11.660 ;
        RECT 160.610 11.800 160.930 11.860 ;
        RECT 279.305 11.800 279.595 11.845 ;
        RECT 327.605 11.800 327.895 11.845 ;
        RECT 160.610 11.660 230.300 11.800 ;
        RECT 160.610 11.600 160.930 11.660 ;
        RECT 211.685 11.460 211.975 11.505 ;
        RECT 213.525 11.460 213.815 11.505 ;
        RECT 211.685 11.320 213.815 11.460 ;
        RECT 230.160 11.460 230.300 11.660 ;
        RECT 279.305 11.660 327.895 11.800 ;
        RECT 279.305 11.615 279.595 11.660 ;
        RECT 327.605 11.615 327.895 11.660 ;
        RECT 391.550 11.800 391.840 11.845 ;
        RECT 393.870 11.800 394.160 11.845 ;
        RECT 395.250 11.800 395.540 11.845 ;
        RECT 400.285 11.800 400.575 11.845 ;
        RECT 391.550 11.660 395.540 11.800 ;
        RECT 391.550 11.615 391.840 11.660 ;
        RECT 393.870 11.615 394.160 11.660 ;
        RECT 395.250 11.615 395.540 11.660 ;
        RECT 395.760 11.660 400.575 11.800 ;
        RECT 395.760 11.460 395.900 11.660 ;
        RECT 400.285 11.615 400.575 11.660 ;
        RECT 230.160 11.320 395.900 11.460 ;
        RECT 211.685 11.275 211.975 11.320 ;
        RECT 213.525 11.275 213.815 11.320 ;
        RECT 228.230 10.100 228.550 10.160 ;
        RECT 266.870 10.100 267.190 10.160 ;
        RECT 228.230 9.960 267.190 10.100 ;
        RECT 228.230 9.900 228.550 9.960 ;
        RECT 266.870 9.900 267.190 9.960 ;
        RECT 273.310 10.100 273.630 10.160 ;
        RECT 279.750 10.100 280.070 10.160 ;
        RECT 273.310 9.960 280.070 10.100 ;
        RECT 273.310 9.900 273.630 9.960 ;
        RECT 279.750 9.900 280.070 9.960 ;
        RECT 375.445 10.100 375.735 10.145 ;
        RECT 396.130 10.100 396.450 10.160 ;
        RECT 375.445 9.960 396.450 10.100 ;
        RECT 375.445 9.915 375.735 9.960 ;
        RECT 396.130 9.900 396.450 9.960 ;
        RECT 306.445 9.420 306.735 9.465 ;
        RECT 318.390 9.420 318.710 9.480 ;
        RECT 449.965 9.420 450.255 9.465 ;
        RECT 306.445 9.280 450.255 9.420 ;
        RECT 306.445 9.235 306.735 9.280 ;
        RECT 318.390 9.220 318.710 9.280 ;
        RECT 449.965 9.235 450.255 9.280 ;
        RECT 179.470 8.740 179.790 8.800 ;
        RECT 269.185 8.740 269.475 8.785 ;
        RECT 179.470 8.600 269.475 8.740 ;
        RECT 179.470 8.540 179.790 8.600 ;
        RECT 269.185 8.555 269.475 8.600 ;
        RECT 269.645 8.740 269.935 8.785 ;
        RECT 330.810 8.740 331.130 8.800 ;
        RECT 269.645 8.600 331.130 8.740 ;
        RECT 269.645 8.555 269.935 8.600 ;
        RECT 330.810 8.540 331.130 8.600 ;
        RECT 54.810 8.400 55.130 8.460 ;
        RECT 282.970 8.400 283.290 8.460 ;
        RECT 54.810 8.260 283.290 8.400 ;
        RECT 54.810 8.200 55.130 8.260 ;
        RECT 282.970 8.200 283.290 8.260 ;
        RECT 213.525 8.060 213.815 8.105 ;
        RECT 426.490 8.060 426.810 8.120 ;
        RECT 213.525 7.920 426.810 8.060 ;
        RECT 213.525 7.875 213.815 7.920 ;
        RECT 426.490 7.860 426.810 7.920 ;
        RECT 255.385 7.720 255.675 7.765 ;
        RECT 269.645 7.720 269.935 7.765 ;
        RECT 255.385 7.580 269.935 7.720 ;
        RECT 255.385 7.535 255.675 7.580 ;
        RECT 269.645 7.535 269.935 7.580 ;
        RECT 279.750 7.720 280.070 7.780 ;
        RECT 399.810 7.720 400.130 7.780 ;
        RECT 279.750 7.580 400.130 7.720 ;
        RECT 279.750 7.520 280.070 7.580 ;
        RECT 399.810 7.520 400.130 7.580 ;
        RECT 269.185 7.380 269.475 7.425 ;
        RECT 298.610 7.380 298.930 7.440 ;
        RECT 269.185 7.240 298.930 7.380 ;
        RECT 269.185 7.195 269.475 7.240 ;
        RECT 298.610 7.180 298.930 7.240 ;
      LAYER via ;
        RECT 10.220 12.960 10.480 13.220 ;
        RECT 225.960 12.960 226.220 13.220 ;
        RECT 197.900 12.620 198.160 12.880 ;
        RECT 210.780 12.620 211.040 12.880 ;
        RECT 156.040 12.280 156.300 12.540 ;
        RECT 167.540 12.280 167.800 12.540 ;
        RECT 184.560 12.280 184.820 12.540 ;
        RECT 193.300 12.280 193.560 12.540 ;
        RECT 199.280 12.280 199.540 12.540 ;
        RECT 207.100 12.280 207.360 12.540 ;
        RECT 210.320 12.280 210.580 12.540 ;
        RECT 263.220 12.960 263.480 13.220 ;
        RECT 228.720 12.280 228.980 12.540 ;
        RECT 238.840 12.280 239.100 12.540 ;
        RECT 268.280 12.960 268.540 13.220 ;
        RECT 396.160 12.960 396.420 13.220 ;
        RECT 400.300 12.960 400.560 13.220 ;
        RECT 451.360 12.960 451.620 13.220 ;
        RECT 298.640 12.620 298.900 12.880 ;
        RECT 309.680 12.620 309.940 12.880 ;
        RECT 265.520 12.280 265.780 12.540 ;
        RECT 326.700 12.280 326.960 12.540 ;
        RECT 353.840 12.280 354.100 12.540 ;
        RECT 392.480 12.280 392.740 12.540 ;
        RECT 399.840 12.280 400.100 12.540 ;
        RECT 400.300 12.280 400.560 12.540 ;
        RECT 145.920 11.940 146.180 12.200 ;
        RECT 228.260 11.940 228.520 12.200 ;
        RECT 242.520 11.940 242.780 12.200 ;
        RECT 266.900 11.940 267.160 12.200 ;
        RECT 304.620 11.940 304.880 12.200 ;
        RECT 530.020 12.620 530.280 12.880 ;
        RECT 457.800 12.280 458.060 12.540 ;
        RECT 160.640 11.600 160.900 11.860 ;
        RECT 228.260 9.900 228.520 10.160 ;
        RECT 266.900 9.900 267.160 10.160 ;
        RECT 273.340 9.900 273.600 10.160 ;
        RECT 279.780 9.900 280.040 10.160 ;
        RECT 396.160 9.900 396.420 10.160 ;
        RECT 318.420 9.220 318.680 9.480 ;
        RECT 179.500 8.540 179.760 8.800 ;
        RECT 330.840 8.540 331.100 8.800 ;
        RECT 54.840 8.200 55.100 8.460 ;
        RECT 283.000 8.200 283.260 8.460 ;
        RECT 426.520 7.860 426.780 8.120 ;
        RECT 279.780 7.520 280.040 7.780 ;
        RECT 399.840 7.520 400.100 7.780 ;
        RECT 298.640 7.180 298.900 7.440 ;
        RECT 9.760 155.760 10.020 156.020 ;
        RECT 8.840 152.700 9.100 152.960 ;
        RECT 8.380 126.180 8.640 126.440 ;
        RECT 8.380 90.140 8.640 90.400 ;
        RECT 13.440 23.840 13.700 24.100 ;
        RECT 13.440 20.440 13.700 20.700 ;
        RECT 10.680 20.100 10.940 20.360 ;
        RECT 11.600 20.100 11.860 20.360 ;
        RECT 10.220 18.400 10.480 18.660 ;
        RECT 8.840 17.720 9.100 17.980 ;
        RECT 10.680 17.380 10.940 17.640 ;
        RECT 9.760 14.660 10.020 14.920 ;
      LAYER met2 ;
        RECT 9.760 155.730 10.020 156.050 ;
        RECT 8.840 152.670 9.100 152.990 ;
        RECT 8.380 126.150 8.640 126.470 ;
        RECT 8.440 90.430 8.580 126.150 ;
        RECT 8.380 90.110 8.640 90.430 ;
        RECT 8.900 18.010 9.040 152.670 ;
        RECT 8.840 17.690 9.100 18.010 ;
        RECT 9.820 14.950 9.960 155.730 ;
        RECT 13.700 24.130 2905.260 3506.300 ;
        RECT 13.440 23.810 2905.260 24.130 ;
        RECT 13.500 20.730 13.640 23.810 ;
        RECT 13.700 20.730 2905.260 23.810 ;
        RECT 13.440 20.410 2905.260 20.730 ;
        RECT 10.680 20.070 10.940 20.390 ;
        RECT 11.600 20.245 11.860 20.390 ;
        RECT 10.220 18.370 10.480 18.690 ;
        RECT 9.760 14.630 10.020 14.950 ;
        RECT 10.280 13.250 10.420 18.370 ;
        RECT 10.740 17.670 10.880 20.070 ;
        RECT 11.590 19.875 11.870 20.245 ;
        RECT 10.680 17.350 10.940 17.670 ;
        RECT 13.700 13.700 2905.260 20.410 ;
        RECT 10.220 12.930 10.480 13.250 ;
        RECT 54.900 8.490 55.040 13.700 ;
        RECT 145.060 13.445 145.200 13.700 ;
        RECT 144.990 13.075 145.270 13.445 ;
        RECT 145.980 12.230 146.120 13.700 ;
        RECT 156.100 12.570 156.240 13.700 ;
        RECT 156.040 12.250 156.300 12.570 ;
        RECT 145.920 11.910 146.180 12.230 ;
        RECT 160.700 11.890 160.840 13.700 ;
        RECT 167.600 12.570 167.740 13.700 ;
        RECT 167.540 12.250 167.800 12.570 ;
        RECT 160.640 11.570 160.900 11.890 ;
        RECT 179.560 8.830 179.700 13.700 ;
        RECT 183.700 13.445 183.840 13.700 ;
        RECT 183.630 13.075 183.910 13.445 ;
        RECT 184.620 12.570 184.760 13.700 ;
        RECT 193.360 12.570 193.500 13.700 ;
        RECT 184.560 12.250 184.820 12.570 ;
        RECT 193.300 12.250 193.560 12.570 ;
        RECT 194.280 11.405 194.420 13.700 ;
        RECT 194.740 13.445 194.880 13.700 ;
        RECT 194.670 13.075 194.950 13.445 ;
        RECT 197.960 12.910 198.100 13.700 ;
        RECT 198.420 13.445 198.560 13.700 ;
        RECT 198.350 13.075 198.630 13.445 ;
        RECT 197.900 12.590 198.160 12.910 ;
        RECT 199.340 12.570 199.480 13.700 ;
        RECT 207.160 12.570 207.300 13.700 ;
        RECT 210.380 12.570 210.520 13.700 ;
        RECT 210.840 12.910 210.980 13.700 ;
        RECT 226.020 13.250 226.160 13.700 ;
        RECT 225.960 12.930 226.220 13.250 ;
        RECT 210.780 12.590 211.040 12.910 ;
        RECT 199.280 12.250 199.540 12.570 ;
        RECT 207.100 12.250 207.360 12.570 ;
        RECT 210.320 12.250 210.580 12.570 ;
        RECT 228.320 12.230 228.460 13.700 ;
        RECT 228.710 12.395 228.990 12.765 ;
        RECT 238.900 12.570 239.040 13.700 ;
        RECT 239.820 13.445 239.960 13.700 ;
        RECT 239.750 13.075 240.030 13.445 ;
        RECT 228.720 12.250 228.980 12.395 ;
        RECT 238.840 12.250 239.100 12.570 ;
        RECT 228.260 11.910 228.520 12.230 ;
        RECT 194.210 11.035 194.490 11.405 ;
        RECT 228.320 10.190 228.460 11.910 ;
        RECT 241.200 11.405 241.340 13.700 ;
        RECT 242.580 12.230 242.720 13.700 ;
        RECT 263.280 13.250 263.420 13.700 ;
        RECT 263.220 12.930 263.480 13.250 ;
        RECT 265.580 12.570 265.720 13.700 ;
        RECT 268.800 13.330 268.940 13.700 ;
        RECT 269.720 13.330 269.860 13.700 ;
        RECT 268.280 12.930 268.540 13.250 ;
        RECT 268.800 13.190 269.860 13.330 ;
        RECT 268.340 12.650 268.480 12.930 ;
        RECT 265.520 12.250 265.780 12.570 ;
        RECT 266.960 12.510 268.480 12.650 ;
        RECT 266.960 12.230 267.100 12.510 ;
        RECT 242.520 11.910 242.780 12.230 ;
        RECT 266.900 11.910 267.160 12.230 ;
        RECT 241.130 11.035 241.410 11.405 ;
        RECT 266.960 10.190 267.100 11.910 ;
        RECT 273.400 10.190 273.540 13.700 ;
        RECT 279.840 10.190 279.980 13.700 ;
        RECT 228.260 9.870 228.520 10.190 ;
        RECT 266.900 9.870 267.160 10.190 ;
        RECT 273.340 9.870 273.600 10.190 ;
        RECT 279.780 9.870 280.040 10.190 ;
        RECT 179.500 8.510 179.760 8.830 ;
        RECT 54.840 8.170 55.100 8.490 ;
        RECT 279.840 7.810 279.980 9.870 ;
        RECT 283.060 8.490 283.200 13.700 ;
        RECT 287.660 13.445 287.800 13.700 ;
        RECT 287.590 13.075 287.870 13.445 ;
        RECT 298.700 12.910 298.840 13.700 ;
        RECT 298.640 12.590 298.900 12.910 ;
        RECT 283.000 8.170 283.260 8.490 ;
        RECT 279.780 7.490 280.040 7.810 ;
        RECT 298.700 7.470 298.840 12.590 ;
        RECT 304.680 12.230 304.820 13.700 ;
        RECT 309.740 12.910 309.880 13.700 ;
        RECT 313.810 13.075 314.090 13.445 ;
        RECT 309.680 12.590 309.940 12.910 ;
        RECT 304.620 11.910 304.880 12.230 ;
        RECT 313.880 11.405 314.020 13.075 ;
        RECT 313.810 11.035 314.090 11.405 ;
        RECT 318.480 9.510 318.620 13.700 ;
        RECT 326.760 12.570 326.900 13.700 ;
        RECT 326.700 12.250 326.960 12.570 ;
        RECT 318.420 9.190 318.680 9.510 ;
        RECT 330.900 8.830 331.040 13.700 ;
        RECT 335.960 11.405 336.100 13.700 ;
        RECT 353.900 12.570 354.040 13.700 ;
        RECT 392.540 12.570 392.680 13.700 ;
        RECT 396.220 13.250 396.360 13.700 ;
        RECT 396.160 12.930 396.420 13.250 ;
        RECT 400.300 12.930 400.560 13.250 ;
        RECT 353.840 12.250 354.100 12.570 ;
        RECT 392.480 12.250 392.740 12.570 ;
        RECT 335.890 11.035 336.170 11.405 ;
        RECT 396.220 10.190 396.360 12.930 ;
        RECT 400.360 12.570 400.500 12.930 ;
        RECT 399.840 12.250 400.100 12.570 ;
        RECT 400.300 12.250 400.560 12.570 ;
        RECT 396.160 9.870 396.420 10.190 ;
        RECT 330.840 8.510 331.100 8.830 ;
        RECT 399.900 7.810 400.040 12.250 ;
        RECT 426.580 8.150 426.720 13.700 ;
        RECT 451.420 13.250 451.560 13.700 ;
        RECT 451.360 12.930 451.620 13.250 ;
        RECT 457.860 12.570 458.000 13.700 ;
        RECT 490.980 12.765 491.120 13.700 ;
        RECT 530.080 12.910 530.220 13.700 ;
        RECT 457.800 12.250 458.060 12.570 ;
        RECT 490.910 12.395 491.190 12.765 ;
        RECT 530.020 12.590 530.280 12.910 ;
        RECT 426.520 7.830 426.780 8.150 ;
        RECT 399.840 7.490 400.100 7.810 ;
        RECT 298.640 7.150 298.900 7.470 ;
      LAYER via2 ;
        RECT 144.990 13.120 145.270 13.400 ;
        RECT 183.630 13.120 183.910 13.400 ;
        RECT 194.670 13.120 194.950 13.400 ;
        RECT 198.350 13.120 198.630 13.400 ;
        RECT 228.710 12.440 228.990 12.720 ;
        RECT 239.750 13.120 240.030 13.400 ;
        RECT 194.210 11.080 194.490 11.360 ;
        RECT 241.130 11.080 241.410 11.360 ;
        RECT 287.590 13.120 287.870 13.400 ;
        RECT 313.810 13.120 314.090 13.400 ;
        RECT 313.810 11.080 314.090 11.360 ;
        RECT 335.890 11.080 336.170 11.360 ;
        RECT 490.910 12.440 491.190 12.720 ;
        RECT 11.590 19.920 11.870 20.200 ;
      LAYER met3 ;
        RECT 11.565 20.210 11.895 20.225 ;
        RECT 13.700 20.210 2906.300 3506.245 ;
        RECT 11.565 19.910 2906.300 20.210 ;
        RECT 11.565 19.895 11.895 19.910 ;
        RECT 13.700 13.700 2906.300 19.910 ;
        RECT 144.965 13.410 145.295 13.425 ;
        RECT 183.605 13.410 183.935 13.425 ;
        RECT 144.965 13.110 183.935 13.410 ;
        RECT 144.965 13.095 145.295 13.110 ;
        RECT 183.605 13.095 183.935 13.110 ;
        RECT 194.645 13.410 194.975 13.425 ;
        RECT 198.325 13.410 198.655 13.425 ;
        RECT 194.645 13.110 198.655 13.410 ;
        RECT 194.645 13.095 194.975 13.110 ;
        RECT 198.325 13.095 198.655 13.110 ;
        RECT 239.725 13.410 240.055 13.425 ;
        RECT 287.565 13.410 287.895 13.425 ;
        RECT 313.785 13.410 314.115 13.425 ;
        RECT 239.725 13.110 314.115 13.410 ;
        RECT 239.725 13.095 240.055 13.110 ;
        RECT 287.565 13.095 287.895 13.110 ;
        RECT 313.785 13.095 314.115 13.110 ;
        RECT 228.685 12.730 229.015 12.745 ;
        RECT 490.885 12.730 491.215 12.745 ;
        RECT 228.685 12.430 491.215 12.730 ;
        RECT 228.685 12.415 229.015 12.430 ;
        RECT 490.885 12.415 491.215 12.430 ;
        RECT 194.185 11.370 194.515 11.385 ;
        RECT 241.105 11.370 241.435 11.385 ;
        RECT 194.185 11.070 241.435 11.370 ;
        RECT 194.185 11.055 194.515 11.070 ;
        RECT 241.105 11.055 241.435 11.070 ;
        RECT 313.785 11.370 314.115 11.385 ;
        RECT 335.865 11.370 336.195 11.385 ;
        RECT 313.785 11.070 336.195 11.370 ;
        RECT 313.785 11.055 314.115 11.070 ;
        RECT 335.865 11.055 336.195 11.070 ;
      LAYER met4 ;
        RECT 49.020 13.700 2887.020 3506.300 ;
      LAYER met5 ;
        RECT 13.700 54.130 2906.300 3477.150 ;
  END
END user_project_wrapper
END LIBRARY

