magic
tech sky130A
magscale 1 2
timestamp 1608218642
<< obsli1 >>
rect 1104 2159 11960 13073
<< obsm1 >>
rect 658 2128 12314 13104
<< metal2 >>
rect 662 14440 718 15240
rect 2042 14440 2098 15240
rect 3514 14440 3570 15240
rect 4986 14440 5042 15240
rect 6458 14440 6514 15240
rect 7838 14440 7894 15240
rect 9310 14440 9366 15240
rect 10782 14440 10838 15240
rect 12254 14440 12310 15240
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4986 0 5042 800
rect 6458 0 6514 800
rect 7838 0 7894 800
rect 9310 0 9366 800
rect 10782 0 10838 800
rect 12254 0 12310 800
<< obsm2 >>
rect 774 14384 1986 14440
rect 2154 14384 3458 14440
rect 3626 14384 4930 14440
rect 5098 14384 6402 14440
rect 6570 14384 7782 14440
rect 7950 14384 9254 14440
rect 9422 14384 10726 14440
rect 10894 14384 12198 14440
rect 664 856 12308 14384
rect 774 800 1986 856
rect 2154 800 3458 856
rect 3626 800 4930 856
rect 5098 800 6402 856
rect 6570 800 7782 856
rect 7950 800 9254 856
rect 9422 800 10726 856
rect 10894 800 12198 856
<< metal3 >>
rect 0 13880 800 14000
rect 12296 13880 13096 14000
rect 0 11296 800 11416
rect 12296 11296 13096 11416
rect 0 8848 800 8968
rect 12296 8848 13096 8968
rect 0 6264 800 6384
rect 12296 6264 13096 6384
rect 0 3680 800 3800
rect 12296 3680 13096 3800
rect 0 1232 800 1352
rect 12296 1232 13096 1352
<< obsm3 >>
rect 880 13800 12216 13973
rect 800 11496 12296 13800
rect 880 11216 12216 11496
rect 800 9048 12296 11216
rect 880 8768 12216 9048
rect 800 6464 12296 8768
rect 880 6184 12216 6464
rect 800 3880 12296 6184
rect 880 3600 12216 3880
rect 800 1432 12296 3600
rect 880 1259 12216 1432
<< metal4 >>
rect 2753 2128 3073 13104
rect 4563 2128 4883 13104
rect 6372 2128 6692 13104
rect 8181 2128 8501 13104
rect 9991 2128 10311 13104
<< obsm4 >>
rect 4963 2128 6292 13104
rect 6772 2128 8101 13104
rect 8581 2128 9911 13104
<< labels >>
rlabel metal2 s 3514 14440 3570 15240 6 cbitin
port 1 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 cbitout
port 2 nsew signal output
rlabel metal2 s 2042 14440 2098 15240 6 confclk
port 3 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 confclko
port 4 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 dempty
port 5 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 din[0]
port 6 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 din[1]
port 7 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 dout[0]
port 8 nsew signal output
rlabel metal2 s 4986 0 5042 800 6 dout[1]
port 9 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 hempty
port 10 nsew signal output
rlabel metal3 s 12296 8848 13096 8968 6 hempty2
port 11 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 lempty
port 12 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 lin[0]
port 13 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 lin[1]
port 14 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 lout[0]
port 15 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 lout[1]
port 16 nsew signal output
rlabel metal3 s 12296 6264 13096 6384 6 rempty
port 17 nsew signal input
rlabel metal2 s 662 14440 718 15240 6 reset
port 18 nsew signal input
rlabel metal2 s 662 0 718 800 6 reseto
port 19 nsew signal output
rlabel metal3 s 12296 3680 13096 3800 6 rin[0]
port 20 nsew signal input
rlabel metal3 s 12296 1232 13096 1352 6 rin[1]
port 21 nsew signal input
rlabel metal3 s 12296 13880 13096 14000 6 rout[0]
port 22 nsew signal output
rlabel metal3 s 12296 11296 13096 11416 6 rout[1]
port 23 nsew signal output
rlabel metal2 s 7838 14440 7894 15240 6 uempty
port 24 nsew signal input
rlabel metal2 s 6458 14440 6514 15240 6 uin[0]
port 25 nsew signal input
rlabel metal2 s 4986 14440 5042 15240 6 uin[1]
port 26 nsew signal input
rlabel metal2 s 12254 14440 12310 15240 6 uout[0]
port 27 nsew signal output
rlabel metal2 s 10782 14440 10838 15240 6 uout[1]
port 28 nsew signal output
rlabel metal2 s 9310 14440 9366 15240 6 vempty
port 29 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 vempty2
port 30 nsew signal output
rlabel metal4 s 9991 2128 10311 13104 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 6372 2128 6692 13104 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 2753 2128 3073 13104 6 vccd1
port 33 nsew power bidirectional
rlabel metal4 s 8181 2128 8501 13104 6 vssd1
port 34 nsew ground bidirectional
rlabel metal4 s 4563 2128 4883 13104 6 vssd1
port 35 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 13096 15240
string LEFview TRUE
<< end >>
