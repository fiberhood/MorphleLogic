*---------------------------------------------------------------------------
* SPDX-FileCopyrightText: 2020 Efabless Corporation
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*---------------------------------------------------------------------------
* NGSPICE file created from sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hvl__decap_8 abstract view
.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__decap_4 abstract view
.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__lsbufhv2lv_1 abstract view
.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_2 abstract view
.subckt sky130_fd_sc_hvl__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_1 abstract view
.subckt sky130_fd_sc_hvl__fill_1 VGND VNB VPB VPWR
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped A X VPWR
XFILLER_1_0 VPWR VPWR FILLER_1_0/VPB FILLER_1_0/VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_48 FILLER_0_8/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_4
XFILLER_0_16 FILLER_0_8/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_40 VPWR VPWR FILLER_1_0/VPB FILLER_1_0/VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_32 VPWR VPWR FILLER_1_0/VPB FILLER_1_0/VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_8 VPWR VPWR FILLER_1_0/VPB FILLER_1_0/VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_24 VPWR VPWR FILLER_1_0/VPB FILLER_1_0/VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_48 VPWR VPWR FILLER_1_0/VPB FILLER_1_0/VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_16 VPWR VPWR FILLER_1_0/VPB FILLER_1_0/VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_40 FILLER_2_0/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_0 FILLER_2_0/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_32 FILLER_2_0/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_0 FILLER_0_8/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_24 FILLER_2_0/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_48 FILLER_2_0/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_4
XFILLER_2_16 FILLER_2_0/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_8 FILLER_2_0/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
Xlvlshiftdown A lvlshiftdown/LVPWR VPWR VPWR VPWR FILLER_0_8/VGND X sky130_fd_sc_hvl__lsbufhv2lv_1
XFILLER_0_8 FILLER_0_8/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_40 FILLER_0_8/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_20 FILLER_0_8/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__fill_2
XFILLER_0_22 FILLER_0_8/VGND VPWR VPWR VPWR sky130_fd_sc_hvl__fill_1
.ends

