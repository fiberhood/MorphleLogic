// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module ycell(cbitin, cbitout, confclk, confclko, dempty, hempty, hempty2, lempty, rempty, reset, reseto, uempty, vempty, vempty2, vccd1, vssd1, din, dout, lin, lout, rin, rout, uin, uout);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  input cbitin;
  output cbitout;
  wire \cfg.cnfg[0] ;
  wire \cfg.cnfg[1] ;
  input confclk;
  output confclko;
  input dempty;
  input [1:0] din;
  output [1:0] dout;
  output hempty;
  output hempty2;
  wire \hfsm.clear ;
  wire \hfsm.lin[0] ;
  wire \hfsm.lin[1] ;
  wire \hfsm.lmatch[0] ;
  wire \hfsm.lmatch[1] ;
  wire \hfsm.nlmempty ;
  input lempty;
  input [1:0] lin;
  output [1:0] lout;
  input rempty;
  input reset;
  output reseto;
  input [1:0] rin;
  output [1:0] rout;
  input uempty;
  input [1:0] uin;
  output [1:0] uout;
  input vccd1;
  output vempty;
  output vempty2;
  wire \vfsm.clear ;
  wire \vfsm.lin[0] ;
  wire \vfsm.lin[1] ;
  wire \vfsm.lmatch[0] ;
  wire \vfsm.lmatch[1] ;
  wire \vfsm.nlmempty ;
  input vssd1;
  sky130_fd_sc_hd__decap_8 FILLER_0_106 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_63 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_67 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_79 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_91 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_94 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_10_11 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_10_112 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_10_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_30 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_10_91 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_11_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_11_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_11_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_11_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_12_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_12_21 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_12_25 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_12_90 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_12_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_13_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_12 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_24 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_13_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_13_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_13_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_13_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_14_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_14_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_14_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_79 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_14_91 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_14_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_15_108 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_15_55 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_15_60 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_72 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_84 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_15_96 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_16_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_16_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_16_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_16_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_110 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_17_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_17_23 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_17_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_17_60 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_17_98 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_18_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_18_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_18_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_18_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_106 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_19_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_19_63 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_74 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_19_86 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_19_92 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_19_94 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_59 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_70 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_75 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_87 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_99 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_13 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_18 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_30 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_68 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_7 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_103 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_51 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_57 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_65 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_91 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_109 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_4_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_4_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_4_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_4_73 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_4_89 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_5_104 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_5_112 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_5_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_80 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_5_92 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_6_108 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_6_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_6_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_6_41 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_6_96 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_101 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_7_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_7_23 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_7_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_8_109 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_8_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_8_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_8_91 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_9_114 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_9_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_10 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_11 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_12 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_13 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_14 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_16 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_17 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_18 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_19 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_20 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_21 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_22 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_23 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_24 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_25 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_26 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_27 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_28 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_29 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_30 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_31 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_33 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_34 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_35 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_36 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_37 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_38 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_39 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_40 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_41 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_42 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_43 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_44 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_45 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_46 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_47 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_48 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_49 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_50 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_51 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_52 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_53 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_54 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_55 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_56 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_57 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_58 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_59 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_6 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_60 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_61 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_62 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_63 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_64 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_65 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_66 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_67 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_68 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_69 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_7 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_70 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_71 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_72 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_8 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_9 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__inv_2 _068_ (
    .A(\hfsm.lmatch[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_029_)
  );
  sky130_fd_sc_hd__inv_2 _069_ (
    .A(\hfsm.lmatch[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_030_)
  );
  sky130_fd_sc_hd__nor2_4 _070_ (
    .A(\hfsm.lin[0] ),
    .B(\hfsm.lin[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_031_)
  );
  sky130_fd_sc_hd__or2_4 _071_ (
    .A(\hfsm.nlmempty ),
    .B(_031_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_032_)
  );
  sky130_fd_sc_hd__inv_2 _072_ (
    .A(uout[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_033_)
  );
  sky130_fd_sc_hd__buf_4 _073_ (
    .A(\cfg.cnfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_034_)
  );
  sky130_fd_sc_hd__inv_2 _074_ (
    .A(_034_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_035_)
  );
  sky130_fd_sc_hd__inv_2 _075_ (
    .A(cbitout),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_036_)
  );
  sky130_fd_sc_hd__buf_2 _076_ (
    .A(_036_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_037_)
  );
  sky130_fd_sc_hd__or3_4 _077_ (
    .A(_035_),
    .B(\cfg.cnfg[1] ),
    .C(_037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_038_)
  );
  sky130_fd_sc_hd__inv_2 _078_ (
    .A(uout[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_039_)
  );
  sky130_fd_sc_hd__or3_4 _079_ (
    .A(_034_),
    .B(\cfg.cnfg[1] ),
    .C(_037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_040_)
  );
  sky130_fd_sc_hd__o22a_4 _080_ (
    .A1(_033_),
    .A2(_038_),
    .B1(_039_),
    .B2(_040_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_041_)
  );
  sky130_fd_sc_hd__o22a_4 _081_ (
    .A1(_033_),
    .A2(_040_),
    .B1(_039_),
    .B2(_038_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_042_)
  );
  sky130_fd_sc_hd__nand2_4 _082_ (
    .A(_041_),
    .B(_042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_043_)
  );
  sky130_fd_sc_hd__a32o_4 _083_ (
    .A1(_029_),
    .A2(_030_),
    .A3(_032_),
    .B1(\hfsm.nlmempty ),
    .B2(_043_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\hfsm.nlmempty )
  );
  sky130_fd_sc_hd__or2_4 _084_ (
    .A(\cfg.cnfg[0] ),
    .B(cbitout),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_044_)
  );
  sky130_fd_sc_hd__inv_2 _085_ (
    .A(_044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(vempty)
  );
  sky130_fd_sc_hd__or2_4 _086_ (
    .A(dempty),
    .B(vempty),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_045_)
  );
  sky130_fd_sc_hd__inv_2 _087_ (
    .A(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_046_)
  );
  sky130_fd_sc_hd__inv_2 _088_ (
    .A(\cfg.cnfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_047_)
  );
  sky130_fd_sc_hd__o21a_4 _089_ (
    .A1(_047_),
    .A2(_036_),
    .B1(_044_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_048_)
  );
  sky130_fd_sc_hd__inv_4 _090_ (
    .A(_048_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_049_)
  );
  sky130_fd_sc_hd__inv_2 _091_ (
    .A(reset),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_050_)
  );
  sky130_fd_sc_hd__inv_2 _092_ (
    .A(uempty),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_051_)
  );
  sky130_fd_sc_hd__or4_4 _093_ (
    .A(_051_),
    .B(dempty),
    .C(uout[1]),
    .D(uout[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_052_)
  );
  sky130_fd_sc_hd__inv_2 _094_ (
    .A(_052_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_053_)
  );
  sky130_fd_sc_hd__a32o_4 _095_ (
    .A1(_050_),
    .A2(_044_),
    .A3(_053_),
    .B1(_051_),
    .B2(uin[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_054_)
  );
  sky130_fd_sc_hd__a32o_4 _096_ (
    .A1(\vfsm.lmatch[1] ),
    .A2(\vfsm.lin[1] ),
    .A3(_049_),
    .B1(_048_),
    .B2(_054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(dout[1])
  );
  sky130_fd_sc_hd__o22a_4 _097_ (
    .A1(_046_),
    .A2(dout[1]),
    .B1(din[1]),
    .B2(_045_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(uout[1])
  );
  sky130_fd_sc_hd__nand2_4 _098_ (
    .A(\vfsm.lmatch[1] ),
    .B(\vfsm.lin[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_055_)
  );
  sky130_fd_sc_hd__inv_2 _099_ (
    .A(\vfsm.lmatch[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_056_)
  );
  sky130_fd_sc_hd__nor2_4 _100_ (
    .A(\vfsm.lin[0] ),
    .B(\vfsm.lin[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_057_)
  );
  sky130_fd_sc_hd__or2_4 _101_ (
    .A(_056_),
    .B(_057_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_058_)
  );
  sky130_fd_sc_hd__and2_4 _102_ (
    .A(uin[0]),
    .B(_051_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_059_)
  );
  sky130_fd_sc_hd__inv_2 _103_ (
    .A(_059_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_060_)
  );
  sky130_fd_sc_hd__a32o_4 _104_ (
    .A1(_049_),
    .A2(_055_),
    .A3(_058_),
    .B1(_048_),
    .B2(_060_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_061_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _105_ (
    .A1_N(_046_),
    .A2_N(_061_),
    .B1(din[0]),
    .B2(_046_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(uout[0])
  );
  sky130_fd_sc_hd__inv_2 _106_ (
    .A(\hfsm.nlmempty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_062_)
  );
  sky130_fd_sc_hd__nor2_4 _107_ (
    .A(_062_),
    .B(_042_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_063_)
  );
  sky130_fd_sc_hd__inv_2 _108_ (
    .A(\hfsm.clear ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_064_)
  );
  sky130_fd_sc_hd__o21a_4 _109_ (
    .A1(\hfsm.lmatch[0] ),
    .A2(_063_),
    .B1(_064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\hfsm.lmatch[0] )
  );
  sky130_fd_sc_hd__nor2_4 _110_ (
    .A(_062_),
    .B(_041_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_065_)
  );
  sky130_fd_sc_hd__o21a_4 _111_ (
    .A1(\hfsm.lmatch[1] ),
    .A2(_065_),
    .B1(_064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\hfsm.lmatch[1] )
  );
  sky130_fd_sc_hd__inv_2 _112_ (
    .A(lempty),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_066_)
  );
  sky130_fd_sc_hd__and2_4 _113_ (
    .A(lin[0]),
    .B(_066_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_067_)
  );
  sky130_fd_sc_hd__o21a_4 _114_ (
    .A1(\hfsm.lin[0] ),
    .A2(_067_),
    .B1(_064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\hfsm.lin[0] )
  );
  sky130_fd_sc_hd__o22a_4 _115_ (
    .A1(_034_),
    .A2(\cfg.cnfg[1] ),
    .B1(_035_),
    .B2(_047_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_000_)
  );
  sky130_fd_sc_hd__nor2_4 _116_ (
    .A(cbitout),
    .B(_000_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(hempty)
  );
  sky130_fd_sc_hd__or2_4 _117_ (
    .A(rempty),
    .B(hempty),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_001_)
  );
  sky130_fd_sc_hd__inv_2 _118_ (
    .A(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_002_)
  );
  sky130_fd_sc_hd__or2_4 _119_ (
    .A(\cfg.cnfg[1] ),
    .B(cbitout),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_003_)
  );
  sky130_fd_sc_hd__a32o_4 _120_ (
    .A1(_034_),
    .A2(_047_),
    .A3(_037_),
    .B1(_049_),
    .B2(_003_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_004_)
  );
  sky130_fd_sc_hd__inv_2 _121_ (
    .A(_004_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_005_)
  );
  sky130_fd_sc_hd__inv_2 _122_ (
    .A(lin[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_006_)
  );
  sky130_fd_sc_hd__a2bb2o_4 _123_ (
    .A1_N(_030_),
    .A2_N(_031_),
    .B1(\hfsm.lmatch[1] ),
    .B2(\hfsm.lin[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_007_)
  );
  sky130_fd_sc_hd__o22a_4 _124_ (
    .A1(_067_),
    .A2(_005_),
    .B1(_004_),
    .B2(_007_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(rout[0])
  );
  sky130_fd_sc_hd__a22oi_4 _125_ (
    .A1(_001_),
    .A2(rout[0]),
    .B1(rin[0]),
    .B2(_002_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_008_)
  );
  sky130_fd_sc_hd__inv_4 _126_ (
    .A(_008_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(lout[0])
  );
  sky130_fd_sc_hd__or2_4 _127_ (
    .A(reset),
    .B(hempty),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_009_)
  );
  sky130_fd_sc_hd__or4_4 _128_ (
    .A(_066_),
    .B(rempty),
    .C(lout[1]),
    .D(_009_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_010_)
  );
  sky130_fd_sc_hd__o22a_4 _129_ (
    .A1(lempty),
    .A2(_006_),
    .B1(lout[0]),
    .B2(_010_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_011_)
  );
  sky130_fd_sc_hd__inv_4 _130_ (
    .A(_011_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_012_)
  );
  sky130_fd_sc_hd__a32o_4 _131_ (
    .A1(\hfsm.lmatch[1] ),
    .A2(\hfsm.lin[1] ),
    .A3(_005_),
    .B1(_004_),
    .B2(_012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(rout[1])
  );
  sky130_fd_sc_hd__o22a_4 _132_ (
    .A1(_002_),
    .A2(rout[1]),
    .B1(rin[1]),
    .B2(_001_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(lout[1])
  );
  sky130_fd_sc_hd__o21a_4 _133_ (
    .A1(\hfsm.lin[1] ),
    .A2(_012_),
    .B1(_064_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\hfsm.lin[1] )
  );
  sky130_fd_sc_hd__or4_4 _134_ (
    .A(\vfsm.nlmempty ),
    .B(_059_),
    .C(_057_),
    .D(_054_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_013_)
  );
  sky130_fd_sc_hd__inv_2 _135_ (
    .A(_013_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_014_)
  );
  sky130_fd_sc_hd__or3_4 _136_ (
    .A(reset),
    .B(vempty),
    .C(_014_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\vfsm.clear )
  );
  sky130_fd_sc_hd__or2_4 _137_ (
    .A(\vfsm.lmatch[1] ),
    .B(\vfsm.lmatch[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_015_)
  );
  sky130_fd_sc_hd__or3_4 _138_ (
    .A(_035_),
    .B(_047_),
    .C(_037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_016_)
  );
  sky130_fd_sc_hd__inv_2 _139_ (
    .A(lout[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_017_)
  );
  sky130_fd_sc_hd__or3_4 _140_ (
    .A(_034_),
    .B(_047_),
    .C(_037_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_018_)
  );
  sky130_fd_sc_hd__o22a_4 _141_ (
    .A1(_008_),
    .A2(_016_),
    .B1(_017_),
    .B2(_018_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_019_)
  );
  sky130_fd_sc_hd__o22a_4 _142_ (
    .A1(_008_),
    .A2(_018_),
    .B1(_017_),
    .B2(_016_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_020_)
  );
  sky130_fd_sc_hd__inv_2 _143_ (
    .A(\vfsm.nlmempty ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_021_)
  );
  sky130_fd_sc_hd__or4_4 _144_ (
    .A(\vfsm.lin[0] ),
    .B(\vfsm.lin[1] ),
    .C(\vfsm.lmatch[1] ),
    .D(\vfsm.lmatch[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_022_)
  );
  sky130_fd_sc_hd__a32o_4 _145_ (
    .A1(_015_),
    .A2(_019_),
    .A3(_020_),
    .B1(_021_),
    .B2(_022_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_023_)
  );
  sky130_fd_sc_hd__inv_2 _146_ (
    .A(_023_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\vfsm.nlmempty )
  );
  sky130_fd_sc_hd__nor2_4 _147_ (
    .A(_021_),
    .B(_020_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_024_)
  );
  sky130_fd_sc_hd__inv_2 _148_ (
    .A(\vfsm.clear ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_025_)
  );
  sky130_fd_sc_hd__o21a_4 _149_ (
    .A1(\vfsm.lmatch[0] ),
    .A2(_024_),
    .B1(_025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\vfsm.lmatch[0] )
  );
  sky130_fd_sc_hd__nor2_4 _150_ (
    .A(_021_),
    .B(_019_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_026_)
  );
  sky130_fd_sc_hd__o21a_4 _151_ (
    .A1(\vfsm.lmatch[1] ),
    .A2(_026_),
    .B1(_025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\vfsm.lmatch[1] )
  );
  sky130_fd_sc_hd__o21a_4 _152_ (
    .A1(\vfsm.lin[0] ),
    .A2(_059_),
    .B1(_025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\vfsm.lin[0] )
  );
  sky130_fd_sc_hd__o21a_4 _153_ (
    .A1(\vfsm.lin[1] ),
    .A2(_054_),
    .B1(_025_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\vfsm.lin[1] )
  );
  sky130_fd_sc_hd__inv_2 _154_ (
    .A(_061_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(dout[0])
  );
  sky130_fd_sc_hd__or4_4 _155_ (
    .A(\hfsm.nlmempty ),
    .B(_031_),
    .C(_067_),
    .D(_012_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(_027_)
  );
  sky130_fd_sc_hd__inv_2 _156_ (
    .A(_027_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(_028_)
  );
  sky130_fd_sc_hd__or2_4 _157_ (
    .A(_009_),
    .B(_028_),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\hfsm.clear )
  );
  sky130_fd_sc_hd__buf_2 _158_ (
    .A(confclk),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(confclko)
  );
  sky130_fd_sc_hd__buf_2 _159_ (
    .A(hempty),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(hempty2)
  );
  sky130_fd_sc_hd__buf_2 _160_ (
    .A(reset),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(reseto)
  );
  sky130_fd_sc_hd__buf_2 _161_ (
    .A(vempty),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(vempty2)
  );
  sky130_fd_sc_hd__dfxtp_4 _162_ (
    .CLK(confclk),
    .D(cbitin),
    .Q(\cfg.cnfg[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _163_ (
    .CLK(confclk),
    .D(\cfg.cnfg[0] ),
    .Q(\cfg.cnfg[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__dfxtp_4 _164_ (
    .CLK(confclk),
    .D(\cfg.cnfg[1] ),
    .Q(cbitout),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
endmodule
