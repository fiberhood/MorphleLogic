VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3519.700 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3519.700 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3519.700 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3519.700 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3519.700 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3519.700 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3519.700 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3519.700 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3519.700 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 0.300 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 0.300 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 0.300 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 0.300 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 0.300 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 0.300 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 0.300 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 87.460 2924.800 88.660 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2433.460 2924.800 2434.660 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2668.740 2924.800 2669.940 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2903.340 2924.800 2904.540 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3137.940 2924.800 3139.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3372.540 2924.800 3373.740 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3519.700 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3519.700 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3519.700 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3519.700 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3519.700 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 322.060 2924.800 323.260 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3519.700 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3519.700 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3519.700 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3519.700 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3410.620 0.300 3411.820 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3123.660 0.300 3124.860 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2836.020 0.300 2837.220 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2549.060 0.300 2550.260 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2261.420 0.300 2262.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1974.460 0.300 1975.660 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 556.660 2924.800 557.860 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1686.820 0.300 1688.020 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1471.260 0.300 1472.460 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1255.700 0.300 1256.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 0.300 1041.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 824.580 0.300 825.780 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 609.700 0.300 610.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 394.140 0.300 395.340 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 178.580 0.300 179.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 791.260 2924.800 792.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1025.860 2924.800 1027.060 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1260.460 2924.800 1261.660 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1495.060 2924.800 1496.260 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1729.660 2924.800 1730.860 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1964.260 2924.800 1965.460 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2198.860 2924.800 2200.060 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 204.420 2924.800 205.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2551.100 2924.800 2552.300 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2785.700 2924.800 2786.900 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3020.300 2924.800 3021.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3254.900 2924.800 3256.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3489.500 2924.800 3490.700 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3519.700 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3519.700 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3519.700 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3519.700 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3519.700 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 439.020 2924.800 440.220 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3519.700 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3519.700 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3519.700 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3519.700 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 0.300 3268.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2979.500 0.300 2980.700 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2692.540 0.300 2693.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2404.900 0.300 2406.100 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.940 0.300 2119.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1830.300 0.300 1831.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 673.620 2924.800 674.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 0.300 1544.540 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1327.780 0.300 1328.980 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1112.220 0.300 1113.420 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 896.660 0.300 897.860 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 681.100 0.300 682.300 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 465.540 0.300 466.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 249.980 0.300 251.180 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 35.100 0.300 36.300 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 908.900 2924.800 910.100 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1143.500 2924.800 1144.700 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1378.100 2924.800 1379.300 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1612.700 2924.800 1613.900 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1847.300 2924.800 1848.500 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2081.900 2924.800 2083.100 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2316.500 2924.800 2317.700 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 145.940 2924.800 147.140 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2492.620 2924.800 2493.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2727.220 2924.800 2728.420 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2961.820 2924.800 2963.020 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3196.420 2924.800 3197.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 3431.020 2924.800 3432.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3519.700 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3519.700 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3519.700 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3519.700 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3519.700 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 380.540 2924.800 381.740 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3519.700 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3519.700 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3519.700 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3519.700 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3339.220 0.300 3340.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3051.580 0.300 3052.780 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2764.620 0.300 2765.820 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2476.980 0.300 2478.180 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2189.340 0.300 2190.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1902.380 0.300 1903.580 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 615.140 2924.800 616.340 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1614.740 0.300 1615.940 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 0.300 1401.060 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1184.300 0.300 1185.500 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 968.740 0.300 969.940 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 753.180 0.300 754.380 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 537.620 0.300 538.820 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 322.060 0.300 323.260 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 106.500 0.300 107.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 849.740 2924.800 850.940 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1084.340 2924.800 1085.540 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1318.940 2924.800 1320.140 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1553.540 2924.800 1554.740 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 1788.820 2924.800 1790.020 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2023.420 2924.800 2024.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2919.700 2258.020 2924.800 2259.220 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.910 -4.800 633.470 0.300 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 0.300 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 0.300 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 0.300 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 0.300 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 0.300 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 0.300 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 0.300 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 0.300 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 0.300 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 0.300 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 0.300 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 0.300 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 0.300 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 0.300 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 0.300 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 0.300 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 0.300 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 0.300 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 0.300 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 0.300 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 0.300 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 0.300 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 0.300 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 0.300 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 0.300 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 0.300 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 0.300 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 0.300 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 0.300 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 0.300 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 0.300 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 0.300 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 0.300 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 0.300 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 0.300 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 0.300 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 0.300 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 0.300 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 0.300 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 0.300 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 0.300 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 0.300 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 0.300 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 0.300 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 0.300 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 0.300 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 0.300 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 0.300 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 0.300 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 0.300 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 0.300 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 0.300 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 0.300 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 0.300 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 0.300 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 0.300 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 0.300 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 0.300 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 0.300 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 0.300 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 0.300 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 0.300 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 0.300 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 0.300 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 0.300 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 0.300 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 0.300 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 0.300 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 0.300 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 0.300 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 0.300 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 0.300 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 0.300 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 0.300 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 0.300 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 0.300 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 0.300 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 0.300 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 0.300 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 0.300 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 0.300 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 0.300 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 0.300 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 0.300 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 0.300 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 0.300 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 0.300 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 0.300 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 0.300 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 0.300 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 0.300 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 0.300 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 0.300 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 0.300 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 0.300 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 0.300 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 0.300 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 0.300 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 0.300 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 0.300 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 0.300 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 0.300 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 0.300 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 0.300 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 0.300 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 0.300 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 0.300 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 0.300 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 0.300 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 0.300 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 0.300 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 0.300 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 0.300 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 0.300 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 0.300 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 0.300 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 0.300 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 0.300 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 0.300 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 0.300 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 0.300 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 0.300 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 0.300 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 0.300 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 0.300 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 0.300 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 0.300 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.890 -4.800 639.450 0.300 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 0.300 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 0.300 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 0.300 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 0.300 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 0.300 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 0.300 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 0.300 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 0.300 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 0.300 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 0.300 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 0.300 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 0.300 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 0.300 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 0.300 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 0.300 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 0.300 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 0.300 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 0.300 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 0.300 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 0.300 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 0.300 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 0.300 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 0.300 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 0.300 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 0.300 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 0.300 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 0.300 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 0.300 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 0.300 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 0.300 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 0.300 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 0.300 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 0.300 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 0.300 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 0.300 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 0.300 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 0.300 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 0.300 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.830 -4.800 657.390 0.300 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 0.300 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 0.300 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 0.300 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 0.300 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 0.300 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 0.300 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 0.300 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 0.300 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 0.300 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 0.300 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.310 -4.800 674.870 0.300 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 0.300 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 0.300 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 0.300 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 0.300 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 0.300 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 0.300 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 0.300 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 0.300 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 0.300 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 0.300 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 0.300 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 0.300 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 0.300 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 0.300 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 0.300 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 0.300 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 0.300 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 0.300 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 0.300 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 0.300 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 0.300 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 0.300 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 0.300 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 0.300 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 0.300 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 0.300 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 0.300 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 0.300 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 0.300 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 0.300 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 0.300 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 0.300 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 0.300 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 0.300 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 0.300 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 0.300 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 0.300 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 0.300 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 0.300 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 0.300 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 0.300 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 0.300 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 0.300 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 0.300 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 0.300 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 0.300 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 0.300 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 0.300 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 0.300 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 0.300 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 0.300 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 0.300 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 0.300 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 0.300 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 0.300 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 0.300 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 0.300 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 0.300 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 0.300 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 0.300 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 0.300 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 0.300 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 0.300 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 0.300 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 0.300 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 0.300 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 0.300 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 0.300 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 0.300 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 0.300 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 0.300 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 0.300 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 0.300 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 0.300 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 0.300 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 0.300 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 0.300 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 0.300 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 0.300 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 0.300 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 0.300 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 0.300 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 0.300 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 0.300 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 0.300 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 0.300 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 0.300 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 0.300 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 0.300 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 0.300 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 0.300 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 0.300 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 0.300 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 0.300 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 0.300 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 0.300 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 0.300 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 0.300 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 0.300 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 0.300 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 0.300 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 0.300 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 0.300 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 0.300 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 0.300 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 0.300 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 0.300 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 0.300 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 0.300 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 0.300 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 0.300 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 0.300 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 0.300 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 0.300 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 0.300 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 0.300 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.810 -4.800 663.370 0.300 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 0.300 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 0.300 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 0.300 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 0.300 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 0.300 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 0.300 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 0.300 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 0.300 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 0.300 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 0.300 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 0.300 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 0.300 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 0.300 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 0.300 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 0.300 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 0.300 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 0.300 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 0.300 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 0.300 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 0.300 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 0.300 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 0.300 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 0.300 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 0.300 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 0.300 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 0.300 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 0.300 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 0.300 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 0.300 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 0.300 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 0.300 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 0.300 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 0.300 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 0.300 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 0.300 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 0.300 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 0.300 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 0.300 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 0.300 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 0.300 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 0.300 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 0.300 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 0.300 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 0.300 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 0.300 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 0.300 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 0.300 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 0.300 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 0.300 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 0.300 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 0.300 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 0.300 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 0.300 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 0.300 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 0.300 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 0.300 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 0.300 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 0.300 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 0.300 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 0.300 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 0.300 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 0.300 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 0.300 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 0.300 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 0.300 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 0.300 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 0.300 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 0.300 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 0.300 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 0.300 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 0.300 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 0.300 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 0.300 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 0.300 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 0.300 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 0.300 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 0.300 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 0.300 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 0.300 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 0.300 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 0.300 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 0.300 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 0.300 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 0.300 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 0.300 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 0.300 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 0.300 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 0.300 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 0.300 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 0.300 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 0.300 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 0.300 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 0.300 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.530 -4.800 241.090 0.300 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.010 -4.800 258.570 0.300 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.950 -4.800 276.510 0.300 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 -4.800 294.450 0.300 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.830 -4.800 312.390 0.300 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.770 -4.800 330.330 0.300 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 0.300 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 -4.800 365.750 0.300 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.130 -4.800 383.690 0.300 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.070 -4.800 401.630 0.300 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 -4.800 62.610 0.300 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 0.300 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.490 -4.800 437.050 0.300 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 0.300 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.370 -4.800 472.930 0.300 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 0.300 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.790 -4.800 508.350 0.300 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.730 -4.800 526.290 0.300 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.670 -4.800 544.230 0.300 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.610 -4.800 562.170 0.300 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.550 -4.800 580.110 0.300 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.970 -4.800 86.530 0.300 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.030 -4.800 597.590 0.300 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.970 -4.800 615.530 0.300 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 0.300 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 -4.800 133.910 0.300 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 0.300 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 -4.800 169.790 0.300 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 0.300 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 -4.800 205.210 0.300 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 0.300 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 0.300 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 -4.800 44.670 0.300 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 -4.800 247.070 0.300 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 0.300 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 -4.800 282.490 0.300 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 0.300 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.810 -4.800 318.370 0.300 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 0.300 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.230 -4.800 353.790 0.300 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.170 -4.800 371.730 0.300 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.110 -4.800 389.670 0.300 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.050 -4.800 407.610 0.300 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.030 -4.800 68.590 0.300 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 0.300 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.470 -4.800 443.030 0.300 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.410 -4.800 460.970 0.300 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.350 -4.800 478.910 0.300 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 0.300 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.770 -4.800 514.330 0.300 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 0.300 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.650 -4.800 550.210 0.300 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 0.300 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.530 -4.800 586.090 0.300 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.490 -4.800 92.050 0.300 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.010 -4.800 603.570 0.300 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.950 -4.800 621.510 0.300 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 0.300 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.330 -4.800 139.890 0.300 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 -4.800 157.830 0.300 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.750 -4.800 175.310 0.300 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 0.300 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 -4.800 211.190 0.300 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.570 -4.800 229.130 0.300 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.090 -4.800 50.650 0.300 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.490 -4.800 253.050 0.300 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 0.300 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 -4.800 288.470 0.300 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 -4.800 306.410 0.300 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.790 -4.800 324.350 0.300 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 0.300 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.210 -4.800 359.770 0.300 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 0.300 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.090 -4.800 395.650 0.300 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 0.300 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 0.300 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.510 -4.800 431.070 0.300 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.450 -4.800 449.010 0.300 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.390 -4.800 466.950 0.300 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.330 -4.800 484.890 0.300 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.270 -4.800 502.830 0.300 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.750 -4.800 520.310 0.300 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.690 -4.800 538.250 0.300 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.630 -4.800 556.190 0.300 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 0.300 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.050 -4.800 591.610 0.300 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 -4.800 98.030 0.300 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 0.300 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.930 -4.800 627.490 0.300 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 -4.800 121.950 0.300 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 0.300 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 -4.800 163.810 0.300 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 -4.800 181.290 0.300 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.670 -4.800 199.230 0.300 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.610 -4.800 217.170 0.300 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.550 -4.800 235.110 0.300 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 -4.800 56.630 0.300 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.990 -4.800 80.550 0.300 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 -4.800 104.010 0.300 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.370 -4.800 127.930 0.300 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 0.300 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 0.300 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 3519.700 7.020 3529.000 ;
        RECT 94.020 3519.700 97.020 3529.000 ;
        RECT 184.020 3519.700 187.020 3529.000 ;
        RECT 274.020 3519.700 277.020 3529.000 ;
        RECT 364.020 3519.700 367.020 3529.000 ;
        RECT 454.020 3519.700 457.020 3529.000 ;
        RECT 544.020 3519.700 547.020 3529.000 ;
        RECT 634.020 3519.700 637.020 3529.000 ;
        RECT 724.020 3519.700 727.020 3529.000 ;
        RECT 814.020 3519.700 817.020 3529.000 ;
        RECT 904.020 3519.700 907.020 3529.000 ;
        RECT 994.020 3519.700 997.020 3529.000 ;
        RECT 1084.020 3519.700 1087.020 3529.000 ;
        RECT 1174.020 3519.700 1177.020 3529.000 ;
        RECT 1264.020 3519.700 1267.020 3529.000 ;
        RECT 1354.020 3519.700 1357.020 3529.000 ;
        RECT 1444.020 3519.700 1447.020 3529.000 ;
        RECT 1534.020 3519.700 1537.020 3529.000 ;
        RECT 1624.020 3519.700 1627.020 3529.000 ;
        RECT 1714.020 3519.700 1717.020 3529.000 ;
        RECT 1804.020 3519.700 1807.020 3529.000 ;
        RECT 1894.020 3519.700 1897.020 3529.000 ;
        RECT 1984.020 3519.700 1987.020 3529.000 ;
        RECT 2074.020 3519.700 2077.020 3529.000 ;
        RECT 2164.020 3519.700 2167.020 3529.000 ;
        RECT 2254.020 3519.700 2257.020 3529.000 ;
        RECT 2344.020 3519.700 2347.020 3529.000 ;
        RECT 2434.020 3519.700 2437.020 3529.000 ;
        RECT 2524.020 3519.700 2527.020 3529.000 ;
        RECT 2614.020 3519.700 2617.020 3529.000 ;
        RECT 2704.020 3519.700 2707.020 3529.000 ;
        RECT 2794.020 3519.700 2797.020 3529.000 ;
        RECT 2884.020 3519.700 2887.020 3529.000 ;
        RECT 4.020 -9.320 7.020 0.300 ;
        RECT 94.020 -9.320 97.020 0.300 ;
        RECT 184.020 -9.320 187.020 0.300 ;
        RECT 274.020 -9.320 277.020 0.300 ;
        RECT 364.020 -9.320 367.020 0.300 ;
        RECT 454.020 -9.320 457.020 0.300 ;
        RECT 544.020 -9.320 547.020 0.300 ;
        RECT 634.020 -9.320 637.020 0.300 ;
        RECT 724.020 -9.320 727.020 0.300 ;
        RECT 814.020 -9.320 817.020 0.300 ;
        RECT 904.020 -9.320 907.020 0.300 ;
        RECT 994.020 -9.320 997.020 0.300 ;
        RECT 1084.020 -9.320 1087.020 0.300 ;
        RECT 1174.020 -9.320 1177.020 0.300 ;
        RECT 1264.020 -9.320 1267.020 0.300 ;
        RECT 1354.020 -9.320 1357.020 0.300 ;
        RECT 1444.020 -9.320 1447.020 0.300 ;
        RECT 1534.020 -9.320 1537.020 0.300 ;
        RECT 1624.020 -9.320 1627.020 0.300 ;
        RECT 1714.020 -9.320 1717.020 0.300 ;
        RECT 1804.020 -9.320 1807.020 0.300 ;
        RECT 1894.020 -9.320 1897.020 0.300 ;
        RECT 1984.020 -9.320 1987.020 0.300 ;
        RECT 2074.020 -9.320 2077.020 0.300 ;
        RECT 2164.020 -9.320 2167.020 0.300 ;
        RECT 2254.020 -9.320 2257.020 0.300 ;
        RECT 2344.020 -9.320 2347.020 0.300 ;
        RECT 2434.020 -9.320 2437.020 0.300 ;
        RECT 2524.020 -9.320 2527.020 0.300 ;
        RECT 2614.020 -9.320 2617.020 0.300 ;
        RECT 2704.020 -9.320 2707.020 0.300 ;
        RECT 2794.020 -9.320 2797.020 0.300 ;
        RECT 2884.020 -9.320 2887.020 0.300 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 94.930 3523.010 96.110 3524.190 ;
        RECT 94.930 3521.410 96.110 3522.590 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 274.930 3523.010 276.110 3524.190 ;
        RECT 274.930 3521.410 276.110 3522.590 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 454.930 3523.010 456.110 3524.190 ;
        RECT 454.930 3521.410 456.110 3522.590 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 634.930 3523.010 636.110 3524.190 ;
        RECT 634.930 3521.410 636.110 3522.590 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 814.930 3523.010 816.110 3524.190 ;
        RECT 814.930 3521.410 816.110 3522.590 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 994.930 3523.010 996.110 3524.190 ;
        RECT 994.930 3521.410 996.110 3522.590 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1174.930 3523.010 1176.110 3524.190 ;
        RECT 1174.930 3521.410 1176.110 3522.590 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1354.930 3523.010 1356.110 3524.190 ;
        RECT 1354.930 3521.410 1356.110 3522.590 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1534.930 3523.010 1536.110 3524.190 ;
        RECT 1534.930 3521.410 1536.110 3522.590 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1714.930 3523.010 1716.110 3524.190 ;
        RECT 1714.930 3521.410 1716.110 3522.590 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1894.930 3523.010 1896.110 3524.190 ;
        RECT 1894.930 3521.410 1896.110 3522.590 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 2074.930 3523.010 2076.110 3524.190 ;
        RECT 2074.930 3521.410 2076.110 3522.590 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2254.930 3523.010 2256.110 3524.190 ;
        RECT 2254.930 3521.410 2256.110 3522.590 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2434.930 3523.010 2436.110 3524.190 ;
        RECT 2434.930 3521.410 2436.110 3522.590 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2614.930 3523.010 2616.110 3524.190 ;
        RECT 2614.930 3521.410 2616.110 3522.590 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2794.930 3523.010 2796.110 3524.190 ;
        RECT 2794.930 3521.410 2796.110 3522.590 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT -9.070 3430.850 -7.890 3432.030 ;
        RECT -9.070 3429.250 -7.890 3430.430 ;
        RECT -9.070 3340.850 -7.890 3342.030 ;
        RECT -9.070 3339.250 -7.890 3340.430 ;
        RECT -9.070 3250.850 -7.890 3252.030 ;
        RECT -9.070 3249.250 -7.890 3250.430 ;
        RECT -9.070 3160.850 -7.890 3162.030 ;
        RECT -9.070 3159.250 -7.890 3160.430 ;
        RECT -9.070 3070.850 -7.890 3072.030 ;
        RECT -9.070 3069.250 -7.890 3070.430 ;
        RECT -9.070 2980.850 -7.890 2982.030 ;
        RECT -9.070 2979.250 -7.890 2980.430 ;
        RECT -9.070 2890.850 -7.890 2892.030 ;
        RECT -9.070 2889.250 -7.890 2890.430 ;
        RECT -9.070 2800.850 -7.890 2802.030 ;
        RECT -9.070 2799.250 -7.890 2800.430 ;
        RECT -9.070 2710.850 -7.890 2712.030 ;
        RECT -9.070 2709.250 -7.890 2710.430 ;
        RECT -9.070 2620.850 -7.890 2622.030 ;
        RECT -9.070 2619.250 -7.890 2620.430 ;
        RECT -9.070 2530.850 -7.890 2532.030 ;
        RECT -9.070 2529.250 -7.890 2530.430 ;
        RECT -9.070 2440.850 -7.890 2442.030 ;
        RECT -9.070 2439.250 -7.890 2440.430 ;
        RECT -9.070 2350.850 -7.890 2352.030 ;
        RECT -9.070 2349.250 -7.890 2350.430 ;
        RECT -9.070 2260.850 -7.890 2262.030 ;
        RECT -9.070 2259.250 -7.890 2260.430 ;
        RECT -9.070 2170.850 -7.890 2172.030 ;
        RECT -9.070 2169.250 -7.890 2170.430 ;
        RECT -9.070 2080.850 -7.890 2082.030 ;
        RECT -9.070 2079.250 -7.890 2080.430 ;
        RECT -9.070 1990.850 -7.890 1992.030 ;
        RECT -9.070 1989.250 -7.890 1990.430 ;
        RECT -9.070 1900.850 -7.890 1902.030 ;
        RECT -9.070 1899.250 -7.890 1900.430 ;
        RECT -9.070 1810.850 -7.890 1812.030 ;
        RECT -9.070 1809.250 -7.890 1810.430 ;
        RECT -9.070 1720.850 -7.890 1722.030 ;
        RECT -9.070 1719.250 -7.890 1720.430 ;
        RECT -9.070 1630.850 -7.890 1632.030 ;
        RECT -9.070 1629.250 -7.890 1630.430 ;
        RECT -9.070 1540.850 -7.890 1542.030 ;
        RECT -9.070 1539.250 -7.890 1540.430 ;
        RECT -9.070 1450.850 -7.890 1452.030 ;
        RECT -9.070 1449.250 -7.890 1450.430 ;
        RECT -9.070 1360.850 -7.890 1362.030 ;
        RECT -9.070 1359.250 -7.890 1360.430 ;
        RECT -9.070 1270.850 -7.890 1272.030 ;
        RECT -9.070 1269.250 -7.890 1270.430 ;
        RECT -9.070 1180.850 -7.890 1182.030 ;
        RECT -9.070 1179.250 -7.890 1180.430 ;
        RECT -9.070 1090.850 -7.890 1092.030 ;
        RECT -9.070 1089.250 -7.890 1090.430 ;
        RECT -9.070 1000.850 -7.890 1002.030 ;
        RECT -9.070 999.250 -7.890 1000.430 ;
        RECT -9.070 910.850 -7.890 912.030 ;
        RECT -9.070 909.250 -7.890 910.430 ;
        RECT -9.070 820.850 -7.890 822.030 ;
        RECT -9.070 819.250 -7.890 820.430 ;
        RECT -9.070 730.850 -7.890 732.030 ;
        RECT -9.070 729.250 -7.890 730.430 ;
        RECT -9.070 640.850 -7.890 642.030 ;
        RECT -9.070 639.250 -7.890 640.430 ;
        RECT -9.070 550.850 -7.890 552.030 ;
        RECT -9.070 549.250 -7.890 550.430 ;
        RECT -9.070 460.850 -7.890 462.030 ;
        RECT -9.070 459.250 -7.890 460.430 ;
        RECT -9.070 370.850 -7.890 372.030 ;
        RECT -9.070 369.250 -7.890 370.430 ;
        RECT -9.070 280.850 -7.890 282.030 ;
        RECT -9.070 279.250 -7.890 280.430 ;
        RECT -9.070 190.850 -7.890 192.030 ;
        RECT -9.070 189.250 -7.890 190.430 ;
        RECT -9.070 100.850 -7.890 102.030 ;
        RECT -9.070 99.250 -7.890 100.430 ;
        RECT -9.070 10.850 -7.890 12.030 ;
        RECT -9.070 9.250 -7.890 10.430 ;
        RECT 2927.510 3430.850 2928.690 3432.030 ;
        RECT 2927.510 3429.250 2928.690 3430.430 ;
        RECT 2927.510 3340.850 2928.690 3342.030 ;
        RECT 2927.510 3339.250 2928.690 3340.430 ;
        RECT 2927.510 3250.850 2928.690 3252.030 ;
        RECT 2927.510 3249.250 2928.690 3250.430 ;
        RECT 2927.510 3160.850 2928.690 3162.030 ;
        RECT 2927.510 3159.250 2928.690 3160.430 ;
        RECT 2927.510 3070.850 2928.690 3072.030 ;
        RECT 2927.510 3069.250 2928.690 3070.430 ;
        RECT 2927.510 2980.850 2928.690 2982.030 ;
        RECT 2927.510 2979.250 2928.690 2980.430 ;
        RECT 2927.510 2890.850 2928.690 2892.030 ;
        RECT 2927.510 2889.250 2928.690 2890.430 ;
        RECT 2927.510 2800.850 2928.690 2802.030 ;
        RECT 2927.510 2799.250 2928.690 2800.430 ;
        RECT 2927.510 2710.850 2928.690 2712.030 ;
        RECT 2927.510 2709.250 2928.690 2710.430 ;
        RECT 2927.510 2620.850 2928.690 2622.030 ;
        RECT 2927.510 2619.250 2928.690 2620.430 ;
        RECT 2927.510 2530.850 2928.690 2532.030 ;
        RECT 2927.510 2529.250 2928.690 2530.430 ;
        RECT 2927.510 2440.850 2928.690 2442.030 ;
        RECT 2927.510 2439.250 2928.690 2440.430 ;
        RECT 2927.510 2350.850 2928.690 2352.030 ;
        RECT 2927.510 2349.250 2928.690 2350.430 ;
        RECT 2927.510 2260.850 2928.690 2262.030 ;
        RECT 2927.510 2259.250 2928.690 2260.430 ;
        RECT 2927.510 2170.850 2928.690 2172.030 ;
        RECT 2927.510 2169.250 2928.690 2170.430 ;
        RECT 2927.510 2080.850 2928.690 2082.030 ;
        RECT 2927.510 2079.250 2928.690 2080.430 ;
        RECT 2927.510 1990.850 2928.690 1992.030 ;
        RECT 2927.510 1989.250 2928.690 1990.430 ;
        RECT 2927.510 1900.850 2928.690 1902.030 ;
        RECT 2927.510 1899.250 2928.690 1900.430 ;
        RECT 2927.510 1810.850 2928.690 1812.030 ;
        RECT 2927.510 1809.250 2928.690 1810.430 ;
        RECT 2927.510 1720.850 2928.690 1722.030 ;
        RECT 2927.510 1719.250 2928.690 1720.430 ;
        RECT 2927.510 1630.850 2928.690 1632.030 ;
        RECT 2927.510 1629.250 2928.690 1630.430 ;
        RECT 2927.510 1540.850 2928.690 1542.030 ;
        RECT 2927.510 1539.250 2928.690 1540.430 ;
        RECT 2927.510 1450.850 2928.690 1452.030 ;
        RECT 2927.510 1449.250 2928.690 1450.430 ;
        RECT 2927.510 1360.850 2928.690 1362.030 ;
        RECT 2927.510 1359.250 2928.690 1360.430 ;
        RECT 2927.510 1270.850 2928.690 1272.030 ;
        RECT 2927.510 1269.250 2928.690 1270.430 ;
        RECT 2927.510 1180.850 2928.690 1182.030 ;
        RECT 2927.510 1179.250 2928.690 1180.430 ;
        RECT 2927.510 1090.850 2928.690 1092.030 ;
        RECT 2927.510 1089.250 2928.690 1090.430 ;
        RECT 2927.510 1000.850 2928.690 1002.030 ;
        RECT 2927.510 999.250 2928.690 1000.430 ;
        RECT 2927.510 910.850 2928.690 912.030 ;
        RECT 2927.510 909.250 2928.690 910.430 ;
        RECT 2927.510 820.850 2928.690 822.030 ;
        RECT 2927.510 819.250 2928.690 820.430 ;
        RECT 2927.510 730.850 2928.690 732.030 ;
        RECT 2927.510 729.250 2928.690 730.430 ;
        RECT 2927.510 640.850 2928.690 642.030 ;
        RECT 2927.510 639.250 2928.690 640.430 ;
        RECT 2927.510 550.850 2928.690 552.030 ;
        RECT 2927.510 549.250 2928.690 550.430 ;
        RECT 2927.510 460.850 2928.690 462.030 ;
        RECT 2927.510 459.250 2928.690 460.430 ;
        RECT 2927.510 370.850 2928.690 372.030 ;
        RECT 2927.510 369.250 2928.690 370.430 ;
        RECT 2927.510 280.850 2928.690 282.030 ;
        RECT 2927.510 279.250 2928.690 280.430 ;
        RECT 2927.510 190.850 2928.690 192.030 ;
        RECT 2927.510 189.250 2928.690 190.430 ;
        RECT 2927.510 100.850 2928.690 102.030 ;
        RECT 2927.510 99.250 2928.690 100.430 ;
        RECT 2927.510 10.850 2928.690 12.030 ;
        RECT 2927.510 9.250 2928.690 10.430 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 94.930 -2.910 96.110 -1.730 ;
        RECT 94.930 -4.510 96.110 -3.330 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 274.930 -2.910 276.110 -1.730 ;
        RECT 274.930 -4.510 276.110 -3.330 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 454.930 -2.910 456.110 -1.730 ;
        RECT 454.930 -4.510 456.110 -3.330 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 634.930 -2.910 636.110 -1.730 ;
        RECT 634.930 -4.510 636.110 -3.330 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 814.930 -2.910 816.110 -1.730 ;
        RECT 814.930 -4.510 816.110 -3.330 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 994.930 -2.910 996.110 -1.730 ;
        RECT 994.930 -4.510 996.110 -3.330 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1174.930 -2.910 1176.110 -1.730 ;
        RECT 1174.930 -4.510 1176.110 -3.330 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1354.930 -2.910 1356.110 -1.730 ;
        RECT 1354.930 -4.510 1356.110 -3.330 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1534.930 -2.910 1536.110 -1.730 ;
        RECT 1534.930 -4.510 1536.110 -3.330 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1714.930 -2.910 1716.110 -1.730 ;
        RECT 1714.930 -4.510 1716.110 -3.330 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1894.930 -2.910 1896.110 -1.730 ;
        RECT 1894.930 -4.510 1896.110 -3.330 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2074.930 -2.910 2076.110 -1.730 ;
        RECT 2074.930 -4.510 2076.110 -3.330 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2254.930 -2.910 2256.110 -1.730 ;
        RECT 2254.930 -4.510 2256.110 -3.330 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2434.930 -2.910 2436.110 -1.730 ;
        RECT 2434.930 -4.510 2436.110 -3.330 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2614.930 -2.910 2616.110 -1.730 ;
        RECT 2614.930 -4.510 2616.110 -3.330 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2794.930 -2.910 2796.110 -1.730 ;
        RECT 2794.930 -4.510 2796.110 -3.330 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 94.020 3524.300 97.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 274.020 3524.300 277.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 454.020 3524.300 457.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 634.020 3524.300 637.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 814.020 3524.300 817.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 994.020 3524.300 997.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1174.020 3524.300 1177.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1354.020 3524.300 1357.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1534.020 3524.300 1537.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1714.020 3524.300 1717.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1894.020 3524.300 1897.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2074.020 3524.300 2077.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2254.020 3524.300 2257.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2434.020 3524.300 2437.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2614.020 3524.300 2617.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2794.020 3524.300 2797.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 94.020 3521.290 97.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 274.020 3521.290 277.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 454.020 3521.290 457.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 634.020 3521.290 637.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 814.020 3521.290 817.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 994.020 3521.290 997.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1174.020 3521.290 1177.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1354.020 3521.290 1357.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1534.020 3521.290 1537.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1714.020 3521.290 1717.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1894.020 3521.290 1897.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2074.020 3521.290 2077.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2254.020 3521.290 2257.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2434.020 3521.290 2437.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2614.020 3521.290 2617.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2794.020 3521.290 2797.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.140 -6.980 3432.150 ;
        RECT 2926.600 3432.140 2929.600 3432.150 ;
        RECT -14.680 3429.140 0.300 3432.140 ;
        RECT 2919.700 3429.140 2934.300 3432.140 ;
        RECT -9.980 3429.130 -6.980 3429.140 ;
        RECT 2926.600 3429.130 2929.600 3429.140 ;
        RECT -9.980 3342.140 -6.980 3342.150 ;
        RECT 2926.600 3342.140 2929.600 3342.150 ;
        RECT -14.680 3339.140 0.300 3342.140 ;
        RECT 2919.700 3339.140 2934.300 3342.140 ;
        RECT -9.980 3339.130 -6.980 3339.140 ;
        RECT 2926.600 3339.130 2929.600 3339.140 ;
        RECT -9.980 3252.140 -6.980 3252.150 ;
        RECT 2926.600 3252.140 2929.600 3252.150 ;
        RECT -14.680 3249.140 0.300 3252.140 ;
        RECT 2919.700 3249.140 2934.300 3252.140 ;
        RECT -9.980 3249.130 -6.980 3249.140 ;
        RECT 2926.600 3249.130 2929.600 3249.140 ;
        RECT -9.980 3162.140 -6.980 3162.150 ;
        RECT 2926.600 3162.140 2929.600 3162.150 ;
        RECT -14.680 3159.140 0.300 3162.140 ;
        RECT 2919.700 3159.140 2934.300 3162.140 ;
        RECT -9.980 3159.130 -6.980 3159.140 ;
        RECT 2926.600 3159.130 2929.600 3159.140 ;
        RECT -9.980 3072.140 -6.980 3072.150 ;
        RECT 2926.600 3072.140 2929.600 3072.150 ;
        RECT -14.680 3069.140 0.300 3072.140 ;
        RECT 2919.700 3069.140 2934.300 3072.140 ;
        RECT -9.980 3069.130 -6.980 3069.140 ;
        RECT 2926.600 3069.130 2929.600 3069.140 ;
        RECT -9.980 2982.140 -6.980 2982.150 ;
        RECT 2926.600 2982.140 2929.600 2982.150 ;
        RECT -14.680 2979.140 0.300 2982.140 ;
        RECT 2919.700 2979.140 2934.300 2982.140 ;
        RECT -9.980 2979.130 -6.980 2979.140 ;
        RECT 2926.600 2979.130 2929.600 2979.140 ;
        RECT -9.980 2892.140 -6.980 2892.150 ;
        RECT 2926.600 2892.140 2929.600 2892.150 ;
        RECT -14.680 2889.140 0.300 2892.140 ;
        RECT 2919.700 2889.140 2934.300 2892.140 ;
        RECT -9.980 2889.130 -6.980 2889.140 ;
        RECT 2926.600 2889.130 2929.600 2889.140 ;
        RECT -9.980 2802.140 -6.980 2802.150 ;
        RECT 2926.600 2802.140 2929.600 2802.150 ;
        RECT -14.680 2799.140 0.300 2802.140 ;
        RECT 2919.700 2799.140 2934.300 2802.140 ;
        RECT -9.980 2799.130 -6.980 2799.140 ;
        RECT 2926.600 2799.130 2929.600 2799.140 ;
        RECT -9.980 2712.140 -6.980 2712.150 ;
        RECT 2926.600 2712.140 2929.600 2712.150 ;
        RECT -14.680 2709.140 0.300 2712.140 ;
        RECT 2919.700 2709.140 2934.300 2712.140 ;
        RECT -9.980 2709.130 -6.980 2709.140 ;
        RECT 2926.600 2709.130 2929.600 2709.140 ;
        RECT -9.980 2622.140 -6.980 2622.150 ;
        RECT 2926.600 2622.140 2929.600 2622.150 ;
        RECT -14.680 2619.140 0.300 2622.140 ;
        RECT 2919.700 2619.140 2934.300 2622.140 ;
        RECT -9.980 2619.130 -6.980 2619.140 ;
        RECT 2926.600 2619.130 2929.600 2619.140 ;
        RECT -9.980 2532.140 -6.980 2532.150 ;
        RECT 2926.600 2532.140 2929.600 2532.150 ;
        RECT -14.680 2529.140 0.300 2532.140 ;
        RECT 2919.700 2529.140 2934.300 2532.140 ;
        RECT -9.980 2529.130 -6.980 2529.140 ;
        RECT 2926.600 2529.130 2929.600 2529.140 ;
        RECT -9.980 2442.140 -6.980 2442.150 ;
        RECT 2926.600 2442.140 2929.600 2442.150 ;
        RECT -14.680 2439.140 0.300 2442.140 ;
        RECT 2919.700 2439.140 2934.300 2442.140 ;
        RECT -9.980 2439.130 -6.980 2439.140 ;
        RECT 2926.600 2439.130 2929.600 2439.140 ;
        RECT -9.980 2352.140 -6.980 2352.150 ;
        RECT 2926.600 2352.140 2929.600 2352.150 ;
        RECT -14.680 2349.140 0.300 2352.140 ;
        RECT 2919.700 2349.140 2934.300 2352.140 ;
        RECT -9.980 2349.130 -6.980 2349.140 ;
        RECT 2926.600 2349.130 2929.600 2349.140 ;
        RECT -9.980 2262.140 -6.980 2262.150 ;
        RECT 2926.600 2262.140 2929.600 2262.150 ;
        RECT -14.680 2259.140 0.300 2262.140 ;
        RECT 2919.700 2259.140 2934.300 2262.140 ;
        RECT -9.980 2259.130 -6.980 2259.140 ;
        RECT 2926.600 2259.130 2929.600 2259.140 ;
        RECT -9.980 2172.140 -6.980 2172.150 ;
        RECT 2926.600 2172.140 2929.600 2172.150 ;
        RECT -14.680 2169.140 0.300 2172.140 ;
        RECT 2919.700 2169.140 2934.300 2172.140 ;
        RECT -9.980 2169.130 -6.980 2169.140 ;
        RECT 2926.600 2169.130 2929.600 2169.140 ;
        RECT -9.980 2082.140 -6.980 2082.150 ;
        RECT 2926.600 2082.140 2929.600 2082.150 ;
        RECT -14.680 2079.140 0.300 2082.140 ;
        RECT 2919.700 2079.140 2934.300 2082.140 ;
        RECT -9.980 2079.130 -6.980 2079.140 ;
        RECT 2926.600 2079.130 2929.600 2079.140 ;
        RECT -9.980 1992.140 -6.980 1992.150 ;
        RECT 2926.600 1992.140 2929.600 1992.150 ;
        RECT -14.680 1989.140 0.300 1992.140 ;
        RECT 2919.700 1989.140 2934.300 1992.140 ;
        RECT -9.980 1989.130 -6.980 1989.140 ;
        RECT 2926.600 1989.130 2929.600 1989.140 ;
        RECT -9.980 1902.140 -6.980 1902.150 ;
        RECT 2926.600 1902.140 2929.600 1902.150 ;
        RECT -14.680 1899.140 0.300 1902.140 ;
        RECT 2919.700 1899.140 2934.300 1902.140 ;
        RECT -9.980 1899.130 -6.980 1899.140 ;
        RECT 2926.600 1899.130 2929.600 1899.140 ;
        RECT -9.980 1812.140 -6.980 1812.150 ;
        RECT 2926.600 1812.140 2929.600 1812.150 ;
        RECT -14.680 1809.140 0.300 1812.140 ;
        RECT 2919.700 1809.140 2934.300 1812.140 ;
        RECT -9.980 1809.130 -6.980 1809.140 ;
        RECT 2926.600 1809.130 2929.600 1809.140 ;
        RECT -9.980 1722.140 -6.980 1722.150 ;
        RECT 2926.600 1722.140 2929.600 1722.150 ;
        RECT -14.680 1719.140 0.300 1722.140 ;
        RECT 2919.700 1719.140 2934.300 1722.140 ;
        RECT -9.980 1719.130 -6.980 1719.140 ;
        RECT 2926.600 1719.130 2929.600 1719.140 ;
        RECT -9.980 1632.140 -6.980 1632.150 ;
        RECT 2926.600 1632.140 2929.600 1632.150 ;
        RECT -14.680 1629.140 0.300 1632.140 ;
        RECT 2919.700 1629.140 2934.300 1632.140 ;
        RECT -9.980 1629.130 -6.980 1629.140 ;
        RECT 2926.600 1629.130 2929.600 1629.140 ;
        RECT -9.980 1542.140 -6.980 1542.150 ;
        RECT 2926.600 1542.140 2929.600 1542.150 ;
        RECT -14.680 1539.140 0.300 1542.140 ;
        RECT 2919.700 1539.140 2934.300 1542.140 ;
        RECT -9.980 1539.130 -6.980 1539.140 ;
        RECT 2926.600 1539.130 2929.600 1539.140 ;
        RECT -9.980 1452.140 -6.980 1452.150 ;
        RECT 2926.600 1452.140 2929.600 1452.150 ;
        RECT -14.680 1449.140 0.300 1452.140 ;
        RECT 2919.700 1449.140 2934.300 1452.140 ;
        RECT -9.980 1449.130 -6.980 1449.140 ;
        RECT 2926.600 1449.130 2929.600 1449.140 ;
        RECT -9.980 1362.140 -6.980 1362.150 ;
        RECT 2926.600 1362.140 2929.600 1362.150 ;
        RECT -14.680 1359.140 0.300 1362.140 ;
        RECT 2919.700 1359.140 2934.300 1362.140 ;
        RECT -9.980 1359.130 -6.980 1359.140 ;
        RECT 2926.600 1359.130 2929.600 1359.140 ;
        RECT -9.980 1272.140 -6.980 1272.150 ;
        RECT 2926.600 1272.140 2929.600 1272.150 ;
        RECT -14.680 1269.140 0.300 1272.140 ;
        RECT 2919.700 1269.140 2934.300 1272.140 ;
        RECT -9.980 1269.130 -6.980 1269.140 ;
        RECT 2926.600 1269.130 2929.600 1269.140 ;
        RECT -9.980 1182.140 -6.980 1182.150 ;
        RECT 2926.600 1182.140 2929.600 1182.150 ;
        RECT -14.680 1179.140 0.300 1182.140 ;
        RECT 2919.700 1179.140 2934.300 1182.140 ;
        RECT -9.980 1179.130 -6.980 1179.140 ;
        RECT 2926.600 1179.130 2929.600 1179.140 ;
        RECT -9.980 1092.140 -6.980 1092.150 ;
        RECT 2926.600 1092.140 2929.600 1092.150 ;
        RECT -14.680 1089.140 0.300 1092.140 ;
        RECT 2919.700 1089.140 2934.300 1092.140 ;
        RECT -9.980 1089.130 -6.980 1089.140 ;
        RECT 2926.600 1089.130 2929.600 1089.140 ;
        RECT -9.980 1002.140 -6.980 1002.150 ;
        RECT 2926.600 1002.140 2929.600 1002.150 ;
        RECT -14.680 999.140 0.300 1002.140 ;
        RECT 2919.700 999.140 2934.300 1002.140 ;
        RECT -9.980 999.130 -6.980 999.140 ;
        RECT 2926.600 999.130 2929.600 999.140 ;
        RECT -9.980 912.140 -6.980 912.150 ;
        RECT 2926.600 912.140 2929.600 912.150 ;
        RECT -14.680 909.140 0.300 912.140 ;
        RECT 2919.700 909.140 2934.300 912.140 ;
        RECT -9.980 909.130 -6.980 909.140 ;
        RECT 2926.600 909.130 2929.600 909.140 ;
        RECT -9.980 822.140 -6.980 822.150 ;
        RECT 2926.600 822.140 2929.600 822.150 ;
        RECT -14.680 819.140 0.300 822.140 ;
        RECT 2919.700 819.140 2934.300 822.140 ;
        RECT -9.980 819.130 -6.980 819.140 ;
        RECT 2926.600 819.130 2929.600 819.140 ;
        RECT -9.980 732.140 -6.980 732.150 ;
        RECT 2926.600 732.140 2929.600 732.150 ;
        RECT -14.680 729.140 0.300 732.140 ;
        RECT 2919.700 729.140 2934.300 732.140 ;
        RECT -9.980 729.130 -6.980 729.140 ;
        RECT 2926.600 729.130 2929.600 729.140 ;
        RECT -9.980 642.140 -6.980 642.150 ;
        RECT 2926.600 642.140 2929.600 642.150 ;
        RECT -14.680 639.140 0.300 642.140 ;
        RECT 2919.700 639.140 2934.300 642.140 ;
        RECT -9.980 639.130 -6.980 639.140 ;
        RECT 2926.600 639.130 2929.600 639.140 ;
        RECT -9.980 552.140 -6.980 552.150 ;
        RECT 2926.600 552.140 2929.600 552.150 ;
        RECT -14.680 549.140 0.300 552.140 ;
        RECT 2919.700 549.140 2934.300 552.140 ;
        RECT -9.980 549.130 -6.980 549.140 ;
        RECT 2926.600 549.130 2929.600 549.140 ;
        RECT -9.980 462.140 -6.980 462.150 ;
        RECT 2926.600 462.140 2929.600 462.150 ;
        RECT -14.680 459.140 0.300 462.140 ;
        RECT 2919.700 459.140 2934.300 462.140 ;
        RECT -9.980 459.130 -6.980 459.140 ;
        RECT 2926.600 459.130 2929.600 459.140 ;
        RECT -9.980 372.140 -6.980 372.150 ;
        RECT 2926.600 372.140 2929.600 372.150 ;
        RECT -14.680 369.140 0.300 372.140 ;
        RECT 2919.700 369.140 2934.300 372.140 ;
        RECT -9.980 369.130 -6.980 369.140 ;
        RECT 2926.600 369.130 2929.600 369.140 ;
        RECT -9.980 282.140 -6.980 282.150 ;
        RECT 2926.600 282.140 2929.600 282.150 ;
        RECT -14.680 279.140 0.300 282.140 ;
        RECT 2919.700 279.140 2934.300 282.140 ;
        RECT -9.980 279.130 -6.980 279.140 ;
        RECT 2926.600 279.130 2929.600 279.140 ;
        RECT -9.980 192.140 -6.980 192.150 ;
        RECT 2926.600 192.140 2929.600 192.150 ;
        RECT -14.680 189.140 0.300 192.140 ;
        RECT 2919.700 189.140 2934.300 192.140 ;
        RECT -9.980 189.130 -6.980 189.140 ;
        RECT 2926.600 189.130 2929.600 189.140 ;
        RECT -9.980 102.140 -6.980 102.150 ;
        RECT 2926.600 102.140 2929.600 102.150 ;
        RECT -14.680 99.140 0.300 102.140 ;
        RECT 2919.700 99.140 2934.300 102.140 ;
        RECT -9.980 99.130 -6.980 99.140 ;
        RECT 2926.600 99.130 2929.600 99.140 ;
        RECT -9.980 12.140 -6.980 12.150 ;
        RECT 2926.600 12.140 2929.600 12.150 ;
        RECT -14.680 9.140 0.300 12.140 ;
        RECT 2919.700 9.140 2934.300 12.140 ;
        RECT -9.980 9.130 -6.980 9.140 ;
        RECT 2926.600 9.130 2929.600 9.140 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 94.020 -1.620 97.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 274.020 -1.620 277.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 454.020 -1.620 457.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 634.020 -1.620 637.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 814.020 -1.620 817.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 994.020 -1.620 997.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1174.020 -1.620 1177.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1354.020 -1.620 1357.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1534.020 -1.620 1537.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1714.020 -1.620 1717.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1894.020 -1.620 1897.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2074.020 -1.620 2077.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2254.020 -1.620 2257.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2434.020 -1.620 2437.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2614.020 -1.620 2617.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2794.020 -1.620 2797.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 94.020 -4.630 97.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 274.020 -4.630 277.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 454.020 -4.630 457.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 634.020 -4.630 637.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 814.020 -4.630 817.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 994.020 -4.630 997.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1174.020 -4.630 1177.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1354.020 -4.630 1357.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1534.020 -4.630 1537.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1714.020 -4.630 1717.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1894.020 -4.630 1897.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2074.020 -4.630 2077.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2254.020 -4.630 2257.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2434.020 -4.630 2437.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2614.020 -4.630 2617.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2794.020 -4.630 2797.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 49.020 3519.700 52.020 3529.000 ;
        RECT 139.020 3519.700 142.020 3529.000 ;
        RECT 229.020 3519.700 232.020 3529.000 ;
        RECT 319.020 3519.700 322.020 3529.000 ;
        RECT 409.020 3519.700 412.020 3529.000 ;
        RECT 499.020 3519.700 502.020 3529.000 ;
        RECT 589.020 3519.700 592.020 3529.000 ;
        RECT 679.020 3519.700 682.020 3529.000 ;
        RECT 769.020 3519.700 772.020 3529.000 ;
        RECT 859.020 3519.700 862.020 3529.000 ;
        RECT 949.020 3519.700 952.020 3529.000 ;
        RECT 1039.020 3519.700 1042.020 3529.000 ;
        RECT 1129.020 3519.700 1132.020 3529.000 ;
        RECT 1219.020 3519.700 1222.020 3529.000 ;
        RECT 1309.020 3519.700 1312.020 3529.000 ;
        RECT 1399.020 3519.700 1402.020 3529.000 ;
        RECT 1489.020 3519.700 1492.020 3529.000 ;
        RECT 1579.020 3519.700 1582.020 3529.000 ;
        RECT 1669.020 3519.700 1672.020 3529.000 ;
        RECT 1759.020 3519.700 1762.020 3529.000 ;
        RECT 1849.020 3519.700 1852.020 3529.000 ;
        RECT 1939.020 3519.700 1942.020 3529.000 ;
        RECT 2029.020 3519.700 2032.020 3529.000 ;
        RECT 2119.020 3519.700 2122.020 3529.000 ;
        RECT 2209.020 3519.700 2212.020 3529.000 ;
        RECT 2299.020 3519.700 2302.020 3529.000 ;
        RECT 2389.020 3519.700 2392.020 3529.000 ;
        RECT 2479.020 3519.700 2482.020 3529.000 ;
        RECT 2569.020 3519.700 2572.020 3529.000 ;
        RECT 2659.020 3519.700 2662.020 3529.000 ;
        RECT 2749.020 3519.700 2752.020 3529.000 ;
        RECT 2839.020 3519.700 2842.020 3529.000 ;
        RECT 49.020 -9.320 52.020 0.300 ;
        RECT 139.020 -9.320 142.020 0.300 ;
        RECT 229.020 -9.320 232.020 0.300 ;
        RECT 319.020 -9.320 322.020 0.300 ;
        RECT 409.020 -9.320 412.020 0.300 ;
        RECT 499.020 -9.320 502.020 0.300 ;
        RECT 589.020 -9.320 592.020 0.300 ;
        RECT 679.020 -9.320 682.020 0.300 ;
        RECT 769.020 -9.320 772.020 0.300 ;
        RECT 859.020 -9.320 862.020 0.300 ;
        RECT 949.020 -9.320 952.020 0.300 ;
        RECT 1039.020 -9.320 1042.020 0.300 ;
        RECT 1129.020 -9.320 1132.020 0.300 ;
        RECT 1219.020 -9.320 1222.020 0.300 ;
        RECT 1309.020 -9.320 1312.020 0.300 ;
        RECT 1399.020 -9.320 1402.020 0.300 ;
        RECT 1489.020 -9.320 1492.020 0.300 ;
        RECT 1579.020 -9.320 1582.020 0.300 ;
        RECT 1669.020 -9.320 1672.020 0.300 ;
        RECT 1759.020 -9.320 1762.020 0.300 ;
        RECT 1849.020 -9.320 1852.020 0.300 ;
        RECT 1939.020 -9.320 1942.020 0.300 ;
        RECT 2029.020 -9.320 2032.020 0.300 ;
        RECT 2119.020 -9.320 2122.020 0.300 ;
        RECT 2209.020 -9.320 2212.020 0.300 ;
        RECT 2299.020 -9.320 2302.020 0.300 ;
        RECT 2389.020 -9.320 2392.020 0.300 ;
        RECT 2479.020 -9.320 2482.020 0.300 ;
        RECT 2569.020 -9.320 2572.020 0.300 ;
        RECT 2659.020 -9.320 2662.020 0.300 ;
        RECT 2749.020 -9.320 2752.020 0.300 ;
        RECT 2839.020 -9.320 2842.020 0.300 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT 49.930 3527.710 51.110 3528.890 ;
        RECT 49.930 3526.110 51.110 3527.290 ;
        RECT 139.930 3527.710 141.110 3528.890 ;
        RECT 139.930 3526.110 141.110 3527.290 ;
        RECT 229.930 3527.710 231.110 3528.890 ;
        RECT 229.930 3526.110 231.110 3527.290 ;
        RECT 319.930 3527.710 321.110 3528.890 ;
        RECT 319.930 3526.110 321.110 3527.290 ;
        RECT 409.930 3527.710 411.110 3528.890 ;
        RECT 409.930 3526.110 411.110 3527.290 ;
        RECT 499.930 3527.710 501.110 3528.890 ;
        RECT 499.930 3526.110 501.110 3527.290 ;
        RECT 589.930 3527.710 591.110 3528.890 ;
        RECT 589.930 3526.110 591.110 3527.290 ;
        RECT 679.930 3527.710 681.110 3528.890 ;
        RECT 679.930 3526.110 681.110 3527.290 ;
        RECT 769.930 3527.710 771.110 3528.890 ;
        RECT 769.930 3526.110 771.110 3527.290 ;
        RECT 859.930 3527.710 861.110 3528.890 ;
        RECT 859.930 3526.110 861.110 3527.290 ;
        RECT 949.930 3527.710 951.110 3528.890 ;
        RECT 949.930 3526.110 951.110 3527.290 ;
        RECT 1039.930 3527.710 1041.110 3528.890 ;
        RECT 1039.930 3526.110 1041.110 3527.290 ;
        RECT 1129.930 3527.710 1131.110 3528.890 ;
        RECT 1129.930 3526.110 1131.110 3527.290 ;
        RECT 1219.930 3527.710 1221.110 3528.890 ;
        RECT 1219.930 3526.110 1221.110 3527.290 ;
        RECT 1309.930 3527.710 1311.110 3528.890 ;
        RECT 1309.930 3526.110 1311.110 3527.290 ;
        RECT 1399.930 3527.710 1401.110 3528.890 ;
        RECT 1399.930 3526.110 1401.110 3527.290 ;
        RECT 1489.930 3527.710 1491.110 3528.890 ;
        RECT 1489.930 3526.110 1491.110 3527.290 ;
        RECT 1579.930 3527.710 1581.110 3528.890 ;
        RECT 1579.930 3526.110 1581.110 3527.290 ;
        RECT 1669.930 3527.710 1671.110 3528.890 ;
        RECT 1669.930 3526.110 1671.110 3527.290 ;
        RECT 1759.930 3527.710 1761.110 3528.890 ;
        RECT 1759.930 3526.110 1761.110 3527.290 ;
        RECT 1849.930 3527.710 1851.110 3528.890 ;
        RECT 1849.930 3526.110 1851.110 3527.290 ;
        RECT 1939.930 3527.710 1941.110 3528.890 ;
        RECT 1939.930 3526.110 1941.110 3527.290 ;
        RECT 2029.930 3527.710 2031.110 3528.890 ;
        RECT 2029.930 3526.110 2031.110 3527.290 ;
        RECT 2119.930 3527.710 2121.110 3528.890 ;
        RECT 2119.930 3526.110 2121.110 3527.290 ;
        RECT 2209.930 3527.710 2211.110 3528.890 ;
        RECT 2209.930 3526.110 2211.110 3527.290 ;
        RECT 2299.930 3527.710 2301.110 3528.890 ;
        RECT 2299.930 3526.110 2301.110 3527.290 ;
        RECT 2389.930 3527.710 2391.110 3528.890 ;
        RECT 2389.930 3526.110 2391.110 3527.290 ;
        RECT 2479.930 3527.710 2481.110 3528.890 ;
        RECT 2479.930 3526.110 2481.110 3527.290 ;
        RECT 2569.930 3527.710 2571.110 3528.890 ;
        RECT 2569.930 3526.110 2571.110 3527.290 ;
        RECT 2659.930 3527.710 2661.110 3528.890 ;
        RECT 2659.930 3526.110 2661.110 3527.290 ;
        RECT 2749.930 3527.710 2751.110 3528.890 ;
        RECT 2749.930 3526.110 2751.110 3527.290 ;
        RECT 2839.930 3527.710 2841.110 3528.890 ;
        RECT 2839.930 3526.110 2841.110 3527.290 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT -13.770 3475.850 -12.590 3477.030 ;
        RECT -13.770 3474.250 -12.590 3475.430 ;
        RECT -13.770 3385.850 -12.590 3387.030 ;
        RECT -13.770 3384.250 -12.590 3385.430 ;
        RECT -13.770 3295.850 -12.590 3297.030 ;
        RECT -13.770 3294.250 -12.590 3295.430 ;
        RECT -13.770 3205.850 -12.590 3207.030 ;
        RECT -13.770 3204.250 -12.590 3205.430 ;
        RECT -13.770 3115.850 -12.590 3117.030 ;
        RECT -13.770 3114.250 -12.590 3115.430 ;
        RECT -13.770 3025.850 -12.590 3027.030 ;
        RECT -13.770 3024.250 -12.590 3025.430 ;
        RECT -13.770 2935.850 -12.590 2937.030 ;
        RECT -13.770 2934.250 -12.590 2935.430 ;
        RECT -13.770 2845.850 -12.590 2847.030 ;
        RECT -13.770 2844.250 -12.590 2845.430 ;
        RECT -13.770 2755.850 -12.590 2757.030 ;
        RECT -13.770 2754.250 -12.590 2755.430 ;
        RECT -13.770 2665.850 -12.590 2667.030 ;
        RECT -13.770 2664.250 -12.590 2665.430 ;
        RECT -13.770 2575.850 -12.590 2577.030 ;
        RECT -13.770 2574.250 -12.590 2575.430 ;
        RECT -13.770 2485.850 -12.590 2487.030 ;
        RECT -13.770 2484.250 -12.590 2485.430 ;
        RECT -13.770 2395.850 -12.590 2397.030 ;
        RECT -13.770 2394.250 -12.590 2395.430 ;
        RECT -13.770 2305.850 -12.590 2307.030 ;
        RECT -13.770 2304.250 -12.590 2305.430 ;
        RECT -13.770 2215.850 -12.590 2217.030 ;
        RECT -13.770 2214.250 -12.590 2215.430 ;
        RECT -13.770 2125.850 -12.590 2127.030 ;
        RECT -13.770 2124.250 -12.590 2125.430 ;
        RECT -13.770 2035.850 -12.590 2037.030 ;
        RECT -13.770 2034.250 -12.590 2035.430 ;
        RECT -13.770 1945.850 -12.590 1947.030 ;
        RECT -13.770 1944.250 -12.590 1945.430 ;
        RECT -13.770 1855.850 -12.590 1857.030 ;
        RECT -13.770 1854.250 -12.590 1855.430 ;
        RECT -13.770 1765.850 -12.590 1767.030 ;
        RECT -13.770 1764.250 -12.590 1765.430 ;
        RECT -13.770 1675.850 -12.590 1677.030 ;
        RECT -13.770 1674.250 -12.590 1675.430 ;
        RECT -13.770 1585.850 -12.590 1587.030 ;
        RECT -13.770 1584.250 -12.590 1585.430 ;
        RECT -13.770 1495.850 -12.590 1497.030 ;
        RECT -13.770 1494.250 -12.590 1495.430 ;
        RECT -13.770 1405.850 -12.590 1407.030 ;
        RECT -13.770 1404.250 -12.590 1405.430 ;
        RECT -13.770 1315.850 -12.590 1317.030 ;
        RECT -13.770 1314.250 -12.590 1315.430 ;
        RECT -13.770 1225.850 -12.590 1227.030 ;
        RECT -13.770 1224.250 -12.590 1225.430 ;
        RECT -13.770 1135.850 -12.590 1137.030 ;
        RECT -13.770 1134.250 -12.590 1135.430 ;
        RECT -13.770 1045.850 -12.590 1047.030 ;
        RECT -13.770 1044.250 -12.590 1045.430 ;
        RECT -13.770 955.850 -12.590 957.030 ;
        RECT -13.770 954.250 -12.590 955.430 ;
        RECT -13.770 865.850 -12.590 867.030 ;
        RECT -13.770 864.250 -12.590 865.430 ;
        RECT -13.770 775.850 -12.590 777.030 ;
        RECT -13.770 774.250 -12.590 775.430 ;
        RECT -13.770 685.850 -12.590 687.030 ;
        RECT -13.770 684.250 -12.590 685.430 ;
        RECT -13.770 595.850 -12.590 597.030 ;
        RECT -13.770 594.250 -12.590 595.430 ;
        RECT -13.770 505.850 -12.590 507.030 ;
        RECT -13.770 504.250 -12.590 505.430 ;
        RECT -13.770 415.850 -12.590 417.030 ;
        RECT -13.770 414.250 -12.590 415.430 ;
        RECT -13.770 325.850 -12.590 327.030 ;
        RECT -13.770 324.250 -12.590 325.430 ;
        RECT -13.770 235.850 -12.590 237.030 ;
        RECT -13.770 234.250 -12.590 235.430 ;
        RECT -13.770 145.850 -12.590 147.030 ;
        RECT -13.770 144.250 -12.590 145.430 ;
        RECT -13.770 55.850 -12.590 57.030 ;
        RECT -13.770 54.250 -12.590 55.430 ;
        RECT 2932.210 3475.850 2933.390 3477.030 ;
        RECT 2932.210 3474.250 2933.390 3475.430 ;
        RECT 2932.210 3385.850 2933.390 3387.030 ;
        RECT 2932.210 3384.250 2933.390 3385.430 ;
        RECT 2932.210 3295.850 2933.390 3297.030 ;
        RECT 2932.210 3294.250 2933.390 3295.430 ;
        RECT 2932.210 3205.850 2933.390 3207.030 ;
        RECT 2932.210 3204.250 2933.390 3205.430 ;
        RECT 2932.210 3115.850 2933.390 3117.030 ;
        RECT 2932.210 3114.250 2933.390 3115.430 ;
        RECT 2932.210 3025.850 2933.390 3027.030 ;
        RECT 2932.210 3024.250 2933.390 3025.430 ;
        RECT 2932.210 2935.850 2933.390 2937.030 ;
        RECT 2932.210 2934.250 2933.390 2935.430 ;
        RECT 2932.210 2845.850 2933.390 2847.030 ;
        RECT 2932.210 2844.250 2933.390 2845.430 ;
        RECT 2932.210 2755.850 2933.390 2757.030 ;
        RECT 2932.210 2754.250 2933.390 2755.430 ;
        RECT 2932.210 2665.850 2933.390 2667.030 ;
        RECT 2932.210 2664.250 2933.390 2665.430 ;
        RECT 2932.210 2575.850 2933.390 2577.030 ;
        RECT 2932.210 2574.250 2933.390 2575.430 ;
        RECT 2932.210 2485.850 2933.390 2487.030 ;
        RECT 2932.210 2484.250 2933.390 2485.430 ;
        RECT 2932.210 2395.850 2933.390 2397.030 ;
        RECT 2932.210 2394.250 2933.390 2395.430 ;
        RECT 2932.210 2305.850 2933.390 2307.030 ;
        RECT 2932.210 2304.250 2933.390 2305.430 ;
        RECT 2932.210 2215.850 2933.390 2217.030 ;
        RECT 2932.210 2214.250 2933.390 2215.430 ;
        RECT 2932.210 2125.850 2933.390 2127.030 ;
        RECT 2932.210 2124.250 2933.390 2125.430 ;
        RECT 2932.210 2035.850 2933.390 2037.030 ;
        RECT 2932.210 2034.250 2933.390 2035.430 ;
        RECT 2932.210 1945.850 2933.390 1947.030 ;
        RECT 2932.210 1944.250 2933.390 1945.430 ;
        RECT 2932.210 1855.850 2933.390 1857.030 ;
        RECT 2932.210 1854.250 2933.390 1855.430 ;
        RECT 2932.210 1765.850 2933.390 1767.030 ;
        RECT 2932.210 1764.250 2933.390 1765.430 ;
        RECT 2932.210 1675.850 2933.390 1677.030 ;
        RECT 2932.210 1674.250 2933.390 1675.430 ;
        RECT 2932.210 1585.850 2933.390 1587.030 ;
        RECT 2932.210 1584.250 2933.390 1585.430 ;
        RECT 2932.210 1495.850 2933.390 1497.030 ;
        RECT 2932.210 1494.250 2933.390 1495.430 ;
        RECT 2932.210 1405.850 2933.390 1407.030 ;
        RECT 2932.210 1404.250 2933.390 1405.430 ;
        RECT 2932.210 1315.850 2933.390 1317.030 ;
        RECT 2932.210 1314.250 2933.390 1315.430 ;
        RECT 2932.210 1225.850 2933.390 1227.030 ;
        RECT 2932.210 1224.250 2933.390 1225.430 ;
        RECT 2932.210 1135.850 2933.390 1137.030 ;
        RECT 2932.210 1134.250 2933.390 1135.430 ;
        RECT 2932.210 1045.850 2933.390 1047.030 ;
        RECT 2932.210 1044.250 2933.390 1045.430 ;
        RECT 2932.210 955.850 2933.390 957.030 ;
        RECT 2932.210 954.250 2933.390 955.430 ;
        RECT 2932.210 865.850 2933.390 867.030 ;
        RECT 2932.210 864.250 2933.390 865.430 ;
        RECT 2932.210 775.850 2933.390 777.030 ;
        RECT 2932.210 774.250 2933.390 775.430 ;
        RECT 2932.210 685.850 2933.390 687.030 ;
        RECT 2932.210 684.250 2933.390 685.430 ;
        RECT 2932.210 595.850 2933.390 597.030 ;
        RECT 2932.210 594.250 2933.390 595.430 ;
        RECT 2932.210 505.850 2933.390 507.030 ;
        RECT 2932.210 504.250 2933.390 505.430 ;
        RECT 2932.210 415.850 2933.390 417.030 ;
        RECT 2932.210 414.250 2933.390 415.430 ;
        RECT 2932.210 325.850 2933.390 327.030 ;
        RECT 2932.210 324.250 2933.390 325.430 ;
        RECT 2932.210 235.850 2933.390 237.030 ;
        RECT 2932.210 234.250 2933.390 235.430 ;
        RECT 2932.210 145.850 2933.390 147.030 ;
        RECT 2932.210 144.250 2933.390 145.430 ;
        RECT 2932.210 55.850 2933.390 57.030 ;
        RECT 2932.210 54.250 2933.390 55.430 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 49.930 -7.610 51.110 -6.430 ;
        RECT 49.930 -9.210 51.110 -8.030 ;
        RECT 139.930 -7.610 141.110 -6.430 ;
        RECT 139.930 -9.210 141.110 -8.030 ;
        RECT 229.930 -7.610 231.110 -6.430 ;
        RECT 229.930 -9.210 231.110 -8.030 ;
        RECT 319.930 -7.610 321.110 -6.430 ;
        RECT 319.930 -9.210 321.110 -8.030 ;
        RECT 409.930 -7.610 411.110 -6.430 ;
        RECT 409.930 -9.210 411.110 -8.030 ;
        RECT 499.930 -7.610 501.110 -6.430 ;
        RECT 499.930 -9.210 501.110 -8.030 ;
        RECT 589.930 -7.610 591.110 -6.430 ;
        RECT 589.930 -9.210 591.110 -8.030 ;
        RECT 679.930 -7.610 681.110 -6.430 ;
        RECT 679.930 -9.210 681.110 -8.030 ;
        RECT 769.930 -7.610 771.110 -6.430 ;
        RECT 769.930 -9.210 771.110 -8.030 ;
        RECT 859.930 -7.610 861.110 -6.430 ;
        RECT 859.930 -9.210 861.110 -8.030 ;
        RECT 949.930 -7.610 951.110 -6.430 ;
        RECT 949.930 -9.210 951.110 -8.030 ;
        RECT 1039.930 -7.610 1041.110 -6.430 ;
        RECT 1039.930 -9.210 1041.110 -8.030 ;
        RECT 1129.930 -7.610 1131.110 -6.430 ;
        RECT 1129.930 -9.210 1131.110 -8.030 ;
        RECT 1219.930 -7.610 1221.110 -6.430 ;
        RECT 1219.930 -9.210 1221.110 -8.030 ;
        RECT 1309.930 -7.610 1311.110 -6.430 ;
        RECT 1309.930 -9.210 1311.110 -8.030 ;
        RECT 1399.930 -7.610 1401.110 -6.430 ;
        RECT 1399.930 -9.210 1401.110 -8.030 ;
        RECT 1489.930 -7.610 1491.110 -6.430 ;
        RECT 1489.930 -9.210 1491.110 -8.030 ;
        RECT 1579.930 -7.610 1581.110 -6.430 ;
        RECT 1579.930 -9.210 1581.110 -8.030 ;
        RECT 1669.930 -7.610 1671.110 -6.430 ;
        RECT 1669.930 -9.210 1671.110 -8.030 ;
        RECT 1759.930 -7.610 1761.110 -6.430 ;
        RECT 1759.930 -9.210 1761.110 -8.030 ;
        RECT 1849.930 -7.610 1851.110 -6.430 ;
        RECT 1849.930 -9.210 1851.110 -8.030 ;
        RECT 1939.930 -7.610 1941.110 -6.430 ;
        RECT 1939.930 -9.210 1941.110 -8.030 ;
        RECT 2029.930 -7.610 2031.110 -6.430 ;
        RECT 2029.930 -9.210 2031.110 -8.030 ;
        RECT 2119.930 -7.610 2121.110 -6.430 ;
        RECT 2119.930 -9.210 2121.110 -8.030 ;
        RECT 2209.930 -7.610 2211.110 -6.430 ;
        RECT 2209.930 -9.210 2211.110 -8.030 ;
        RECT 2299.930 -7.610 2301.110 -6.430 ;
        RECT 2299.930 -9.210 2301.110 -8.030 ;
        RECT 2389.930 -7.610 2391.110 -6.430 ;
        RECT 2389.930 -9.210 2391.110 -8.030 ;
        RECT 2479.930 -7.610 2481.110 -6.430 ;
        RECT 2479.930 -9.210 2481.110 -8.030 ;
        RECT 2569.930 -7.610 2571.110 -6.430 ;
        RECT 2569.930 -9.210 2571.110 -8.030 ;
        RECT 2659.930 -7.610 2661.110 -6.430 ;
        RECT 2659.930 -9.210 2661.110 -8.030 ;
        RECT 2749.930 -7.610 2751.110 -6.430 ;
        RECT 2749.930 -9.210 2751.110 -8.030 ;
        RECT 2839.930 -7.610 2841.110 -6.430 ;
        RECT 2839.930 -9.210 2841.110 -8.030 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 49.020 3529.000 52.020 3529.010 ;
        RECT 139.020 3529.000 142.020 3529.010 ;
        RECT 229.020 3529.000 232.020 3529.010 ;
        RECT 319.020 3529.000 322.020 3529.010 ;
        RECT 409.020 3529.000 412.020 3529.010 ;
        RECT 499.020 3529.000 502.020 3529.010 ;
        RECT 589.020 3529.000 592.020 3529.010 ;
        RECT 679.020 3529.000 682.020 3529.010 ;
        RECT 769.020 3529.000 772.020 3529.010 ;
        RECT 859.020 3529.000 862.020 3529.010 ;
        RECT 949.020 3529.000 952.020 3529.010 ;
        RECT 1039.020 3529.000 1042.020 3529.010 ;
        RECT 1129.020 3529.000 1132.020 3529.010 ;
        RECT 1219.020 3529.000 1222.020 3529.010 ;
        RECT 1309.020 3529.000 1312.020 3529.010 ;
        RECT 1399.020 3529.000 1402.020 3529.010 ;
        RECT 1489.020 3529.000 1492.020 3529.010 ;
        RECT 1579.020 3529.000 1582.020 3529.010 ;
        RECT 1669.020 3529.000 1672.020 3529.010 ;
        RECT 1759.020 3529.000 1762.020 3529.010 ;
        RECT 1849.020 3529.000 1852.020 3529.010 ;
        RECT 1939.020 3529.000 1942.020 3529.010 ;
        RECT 2029.020 3529.000 2032.020 3529.010 ;
        RECT 2119.020 3529.000 2122.020 3529.010 ;
        RECT 2209.020 3529.000 2212.020 3529.010 ;
        RECT 2299.020 3529.000 2302.020 3529.010 ;
        RECT 2389.020 3529.000 2392.020 3529.010 ;
        RECT 2479.020 3529.000 2482.020 3529.010 ;
        RECT 2569.020 3529.000 2572.020 3529.010 ;
        RECT 2659.020 3529.000 2662.020 3529.010 ;
        RECT 2749.020 3529.000 2752.020 3529.010 ;
        RECT 2839.020 3529.000 2842.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 49.020 3525.990 52.020 3526.000 ;
        RECT 139.020 3525.990 142.020 3526.000 ;
        RECT 229.020 3525.990 232.020 3526.000 ;
        RECT 319.020 3525.990 322.020 3526.000 ;
        RECT 409.020 3525.990 412.020 3526.000 ;
        RECT 499.020 3525.990 502.020 3526.000 ;
        RECT 589.020 3525.990 592.020 3526.000 ;
        RECT 679.020 3525.990 682.020 3526.000 ;
        RECT 769.020 3525.990 772.020 3526.000 ;
        RECT 859.020 3525.990 862.020 3526.000 ;
        RECT 949.020 3525.990 952.020 3526.000 ;
        RECT 1039.020 3525.990 1042.020 3526.000 ;
        RECT 1129.020 3525.990 1132.020 3526.000 ;
        RECT 1219.020 3525.990 1222.020 3526.000 ;
        RECT 1309.020 3525.990 1312.020 3526.000 ;
        RECT 1399.020 3525.990 1402.020 3526.000 ;
        RECT 1489.020 3525.990 1492.020 3526.000 ;
        RECT 1579.020 3525.990 1582.020 3526.000 ;
        RECT 1669.020 3525.990 1672.020 3526.000 ;
        RECT 1759.020 3525.990 1762.020 3526.000 ;
        RECT 1849.020 3525.990 1852.020 3526.000 ;
        RECT 1939.020 3525.990 1942.020 3526.000 ;
        RECT 2029.020 3525.990 2032.020 3526.000 ;
        RECT 2119.020 3525.990 2122.020 3526.000 ;
        RECT 2209.020 3525.990 2212.020 3526.000 ;
        RECT 2299.020 3525.990 2302.020 3526.000 ;
        RECT 2389.020 3525.990 2392.020 3526.000 ;
        RECT 2479.020 3525.990 2482.020 3526.000 ;
        RECT 2569.020 3525.990 2572.020 3526.000 ;
        RECT 2659.020 3525.990 2662.020 3526.000 ;
        RECT 2749.020 3525.990 2752.020 3526.000 ;
        RECT 2839.020 3525.990 2842.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3477.140 -11.680 3477.150 ;
        RECT 2931.300 3477.140 2934.300 3477.150 ;
        RECT -14.680 3474.140 0.300 3477.140 ;
        RECT 2919.700 3474.140 2934.300 3477.140 ;
        RECT -14.680 3474.130 -11.680 3474.140 ;
        RECT 2931.300 3474.130 2934.300 3474.140 ;
        RECT -14.680 3387.140 -11.680 3387.150 ;
        RECT 2931.300 3387.140 2934.300 3387.150 ;
        RECT -14.680 3384.140 0.300 3387.140 ;
        RECT 2919.700 3384.140 2934.300 3387.140 ;
        RECT -14.680 3384.130 -11.680 3384.140 ;
        RECT 2931.300 3384.130 2934.300 3384.140 ;
        RECT -14.680 3297.140 -11.680 3297.150 ;
        RECT 2931.300 3297.140 2934.300 3297.150 ;
        RECT -14.680 3294.140 0.300 3297.140 ;
        RECT 2919.700 3294.140 2934.300 3297.140 ;
        RECT -14.680 3294.130 -11.680 3294.140 ;
        RECT 2931.300 3294.130 2934.300 3294.140 ;
        RECT -14.680 3207.140 -11.680 3207.150 ;
        RECT 2931.300 3207.140 2934.300 3207.150 ;
        RECT -14.680 3204.140 0.300 3207.140 ;
        RECT 2919.700 3204.140 2934.300 3207.140 ;
        RECT -14.680 3204.130 -11.680 3204.140 ;
        RECT 2931.300 3204.130 2934.300 3204.140 ;
        RECT -14.680 3117.140 -11.680 3117.150 ;
        RECT 2931.300 3117.140 2934.300 3117.150 ;
        RECT -14.680 3114.140 0.300 3117.140 ;
        RECT 2919.700 3114.140 2934.300 3117.140 ;
        RECT -14.680 3114.130 -11.680 3114.140 ;
        RECT 2931.300 3114.130 2934.300 3114.140 ;
        RECT -14.680 3027.140 -11.680 3027.150 ;
        RECT 2931.300 3027.140 2934.300 3027.150 ;
        RECT -14.680 3024.140 0.300 3027.140 ;
        RECT 2919.700 3024.140 2934.300 3027.140 ;
        RECT -14.680 3024.130 -11.680 3024.140 ;
        RECT 2931.300 3024.130 2934.300 3024.140 ;
        RECT -14.680 2937.140 -11.680 2937.150 ;
        RECT 2931.300 2937.140 2934.300 2937.150 ;
        RECT -14.680 2934.140 0.300 2937.140 ;
        RECT 2919.700 2934.140 2934.300 2937.140 ;
        RECT -14.680 2934.130 -11.680 2934.140 ;
        RECT 2931.300 2934.130 2934.300 2934.140 ;
        RECT -14.680 2847.140 -11.680 2847.150 ;
        RECT 2931.300 2847.140 2934.300 2847.150 ;
        RECT -14.680 2844.140 0.300 2847.140 ;
        RECT 2919.700 2844.140 2934.300 2847.140 ;
        RECT -14.680 2844.130 -11.680 2844.140 ;
        RECT 2931.300 2844.130 2934.300 2844.140 ;
        RECT -14.680 2757.140 -11.680 2757.150 ;
        RECT 2931.300 2757.140 2934.300 2757.150 ;
        RECT -14.680 2754.140 0.300 2757.140 ;
        RECT 2919.700 2754.140 2934.300 2757.140 ;
        RECT -14.680 2754.130 -11.680 2754.140 ;
        RECT 2931.300 2754.130 2934.300 2754.140 ;
        RECT -14.680 2667.140 -11.680 2667.150 ;
        RECT 2931.300 2667.140 2934.300 2667.150 ;
        RECT -14.680 2664.140 0.300 2667.140 ;
        RECT 2919.700 2664.140 2934.300 2667.140 ;
        RECT -14.680 2664.130 -11.680 2664.140 ;
        RECT 2931.300 2664.130 2934.300 2664.140 ;
        RECT -14.680 2577.140 -11.680 2577.150 ;
        RECT 2931.300 2577.140 2934.300 2577.150 ;
        RECT -14.680 2574.140 0.300 2577.140 ;
        RECT 2919.700 2574.140 2934.300 2577.140 ;
        RECT -14.680 2574.130 -11.680 2574.140 ;
        RECT 2931.300 2574.130 2934.300 2574.140 ;
        RECT -14.680 2487.140 -11.680 2487.150 ;
        RECT 2931.300 2487.140 2934.300 2487.150 ;
        RECT -14.680 2484.140 0.300 2487.140 ;
        RECT 2919.700 2484.140 2934.300 2487.140 ;
        RECT -14.680 2484.130 -11.680 2484.140 ;
        RECT 2931.300 2484.130 2934.300 2484.140 ;
        RECT -14.680 2397.140 -11.680 2397.150 ;
        RECT 2931.300 2397.140 2934.300 2397.150 ;
        RECT -14.680 2394.140 0.300 2397.140 ;
        RECT 2919.700 2394.140 2934.300 2397.140 ;
        RECT -14.680 2394.130 -11.680 2394.140 ;
        RECT 2931.300 2394.130 2934.300 2394.140 ;
        RECT -14.680 2307.140 -11.680 2307.150 ;
        RECT 2931.300 2307.140 2934.300 2307.150 ;
        RECT -14.680 2304.140 0.300 2307.140 ;
        RECT 2919.700 2304.140 2934.300 2307.140 ;
        RECT -14.680 2304.130 -11.680 2304.140 ;
        RECT 2931.300 2304.130 2934.300 2304.140 ;
        RECT -14.680 2217.140 -11.680 2217.150 ;
        RECT 2931.300 2217.140 2934.300 2217.150 ;
        RECT -14.680 2214.140 0.300 2217.140 ;
        RECT 2919.700 2214.140 2934.300 2217.140 ;
        RECT -14.680 2214.130 -11.680 2214.140 ;
        RECT 2931.300 2214.130 2934.300 2214.140 ;
        RECT -14.680 2127.140 -11.680 2127.150 ;
        RECT 2931.300 2127.140 2934.300 2127.150 ;
        RECT -14.680 2124.140 0.300 2127.140 ;
        RECT 2919.700 2124.140 2934.300 2127.140 ;
        RECT -14.680 2124.130 -11.680 2124.140 ;
        RECT 2931.300 2124.130 2934.300 2124.140 ;
        RECT -14.680 2037.140 -11.680 2037.150 ;
        RECT 2931.300 2037.140 2934.300 2037.150 ;
        RECT -14.680 2034.140 0.300 2037.140 ;
        RECT 2919.700 2034.140 2934.300 2037.140 ;
        RECT -14.680 2034.130 -11.680 2034.140 ;
        RECT 2931.300 2034.130 2934.300 2034.140 ;
        RECT -14.680 1947.140 -11.680 1947.150 ;
        RECT 2931.300 1947.140 2934.300 1947.150 ;
        RECT -14.680 1944.140 0.300 1947.140 ;
        RECT 2919.700 1944.140 2934.300 1947.140 ;
        RECT -14.680 1944.130 -11.680 1944.140 ;
        RECT 2931.300 1944.130 2934.300 1944.140 ;
        RECT -14.680 1857.140 -11.680 1857.150 ;
        RECT 2931.300 1857.140 2934.300 1857.150 ;
        RECT -14.680 1854.140 0.300 1857.140 ;
        RECT 2919.700 1854.140 2934.300 1857.140 ;
        RECT -14.680 1854.130 -11.680 1854.140 ;
        RECT 2931.300 1854.130 2934.300 1854.140 ;
        RECT -14.680 1767.140 -11.680 1767.150 ;
        RECT 2931.300 1767.140 2934.300 1767.150 ;
        RECT -14.680 1764.140 0.300 1767.140 ;
        RECT 2919.700 1764.140 2934.300 1767.140 ;
        RECT -14.680 1764.130 -11.680 1764.140 ;
        RECT 2931.300 1764.130 2934.300 1764.140 ;
        RECT -14.680 1677.140 -11.680 1677.150 ;
        RECT 2931.300 1677.140 2934.300 1677.150 ;
        RECT -14.680 1674.140 0.300 1677.140 ;
        RECT 2919.700 1674.140 2934.300 1677.140 ;
        RECT -14.680 1674.130 -11.680 1674.140 ;
        RECT 2931.300 1674.130 2934.300 1674.140 ;
        RECT -14.680 1587.140 -11.680 1587.150 ;
        RECT 2931.300 1587.140 2934.300 1587.150 ;
        RECT -14.680 1584.140 0.300 1587.140 ;
        RECT 2919.700 1584.140 2934.300 1587.140 ;
        RECT -14.680 1584.130 -11.680 1584.140 ;
        RECT 2931.300 1584.130 2934.300 1584.140 ;
        RECT -14.680 1497.140 -11.680 1497.150 ;
        RECT 2931.300 1497.140 2934.300 1497.150 ;
        RECT -14.680 1494.140 0.300 1497.140 ;
        RECT 2919.700 1494.140 2934.300 1497.140 ;
        RECT -14.680 1494.130 -11.680 1494.140 ;
        RECT 2931.300 1494.130 2934.300 1494.140 ;
        RECT -14.680 1407.140 -11.680 1407.150 ;
        RECT 2931.300 1407.140 2934.300 1407.150 ;
        RECT -14.680 1404.140 0.300 1407.140 ;
        RECT 2919.700 1404.140 2934.300 1407.140 ;
        RECT -14.680 1404.130 -11.680 1404.140 ;
        RECT 2931.300 1404.130 2934.300 1404.140 ;
        RECT -14.680 1317.140 -11.680 1317.150 ;
        RECT 2931.300 1317.140 2934.300 1317.150 ;
        RECT -14.680 1314.140 0.300 1317.140 ;
        RECT 2919.700 1314.140 2934.300 1317.140 ;
        RECT -14.680 1314.130 -11.680 1314.140 ;
        RECT 2931.300 1314.130 2934.300 1314.140 ;
        RECT -14.680 1227.140 -11.680 1227.150 ;
        RECT 2931.300 1227.140 2934.300 1227.150 ;
        RECT -14.680 1224.140 0.300 1227.140 ;
        RECT 2919.700 1224.140 2934.300 1227.140 ;
        RECT -14.680 1224.130 -11.680 1224.140 ;
        RECT 2931.300 1224.130 2934.300 1224.140 ;
        RECT -14.680 1137.140 -11.680 1137.150 ;
        RECT 2931.300 1137.140 2934.300 1137.150 ;
        RECT -14.680 1134.140 0.300 1137.140 ;
        RECT 2919.700 1134.140 2934.300 1137.140 ;
        RECT -14.680 1134.130 -11.680 1134.140 ;
        RECT 2931.300 1134.130 2934.300 1134.140 ;
        RECT -14.680 1047.140 -11.680 1047.150 ;
        RECT 2931.300 1047.140 2934.300 1047.150 ;
        RECT -14.680 1044.140 0.300 1047.140 ;
        RECT 2919.700 1044.140 2934.300 1047.140 ;
        RECT -14.680 1044.130 -11.680 1044.140 ;
        RECT 2931.300 1044.130 2934.300 1044.140 ;
        RECT -14.680 957.140 -11.680 957.150 ;
        RECT 2931.300 957.140 2934.300 957.150 ;
        RECT -14.680 954.140 0.300 957.140 ;
        RECT 2919.700 954.140 2934.300 957.140 ;
        RECT -14.680 954.130 -11.680 954.140 ;
        RECT 2931.300 954.130 2934.300 954.140 ;
        RECT -14.680 867.140 -11.680 867.150 ;
        RECT 2931.300 867.140 2934.300 867.150 ;
        RECT -14.680 864.140 0.300 867.140 ;
        RECT 2919.700 864.140 2934.300 867.140 ;
        RECT -14.680 864.130 -11.680 864.140 ;
        RECT 2931.300 864.130 2934.300 864.140 ;
        RECT -14.680 777.140 -11.680 777.150 ;
        RECT 2931.300 777.140 2934.300 777.150 ;
        RECT -14.680 774.140 0.300 777.140 ;
        RECT 2919.700 774.140 2934.300 777.140 ;
        RECT -14.680 774.130 -11.680 774.140 ;
        RECT 2931.300 774.130 2934.300 774.140 ;
        RECT -14.680 687.140 -11.680 687.150 ;
        RECT 2931.300 687.140 2934.300 687.150 ;
        RECT -14.680 684.140 0.300 687.140 ;
        RECT 2919.700 684.140 2934.300 687.140 ;
        RECT -14.680 684.130 -11.680 684.140 ;
        RECT 2931.300 684.130 2934.300 684.140 ;
        RECT -14.680 597.140 -11.680 597.150 ;
        RECT 2931.300 597.140 2934.300 597.150 ;
        RECT -14.680 594.140 0.300 597.140 ;
        RECT 2919.700 594.140 2934.300 597.140 ;
        RECT -14.680 594.130 -11.680 594.140 ;
        RECT 2931.300 594.130 2934.300 594.140 ;
        RECT -14.680 507.140 -11.680 507.150 ;
        RECT 2931.300 507.140 2934.300 507.150 ;
        RECT -14.680 504.140 0.300 507.140 ;
        RECT 2919.700 504.140 2934.300 507.140 ;
        RECT -14.680 504.130 -11.680 504.140 ;
        RECT 2931.300 504.130 2934.300 504.140 ;
        RECT -14.680 417.140 -11.680 417.150 ;
        RECT 2931.300 417.140 2934.300 417.150 ;
        RECT -14.680 414.140 0.300 417.140 ;
        RECT 2919.700 414.140 2934.300 417.140 ;
        RECT -14.680 414.130 -11.680 414.140 ;
        RECT 2931.300 414.130 2934.300 414.140 ;
        RECT -14.680 327.140 -11.680 327.150 ;
        RECT 2931.300 327.140 2934.300 327.150 ;
        RECT -14.680 324.140 0.300 327.140 ;
        RECT 2919.700 324.140 2934.300 327.140 ;
        RECT -14.680 324.130 -11.680 324.140 ;
        RECT 2931.300 324.130 2934.300 324.140 ;
        RECT -14.680 237.140 -11.680 237.150 ;
        RECT 2931.300 237.140 2934.300 237.150 ;
        RECT -14.680 234.140 0.300 237.140 ;
        RECT 2919.700 234.140 2934.300 237.140 ;
        RECT -14.680 234.130 -11.680 234.140 ;
        RECT 2931.300 234.130 2934.300 234.140 ;
        RECT -14.680 147.140 -11.680 147.150 ;
        RECT 2931.300 147.140 2934.300 147.150 ;
        RECT -14.680 144.140 0.300 147.140 ;
        RECT 2919.700 144.140 2934.300 147.140 ;
        RECT -14.680 144.130 -11.680 144.140 ;
        RECT 2931.300 144.130 2934.300 144.140 ;
        RECT -14.680 57.140 -11.680 57.150 ;
        RECT 2931.300 57.140 2934.300 57.150 ;
        RECT -14.680 54.140 0.300 57.140 ;
        RECT 2919.700 54.140 2934.300 57.140 ;
        RECT -14.680 54.130 -11.680 54.140 ;
        RECT 2931.300 54.130 2934.300 54.140 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 49.020 -6.320 52.020 -6.310 ;
        RECT 139.020 -6.320 142.020 -6.310 ;
        RECT 229.020 -6.320 232.020 -6.310 ;
        RECT 319.020 -6.320 322.020 -6.310 ;
        RECT 409.020 -6.320 412.020 -6.310 ;
        RECT 499.020 -6.320 502.020 -6.310 ;
        RECT 589.020 -6.320 592.020 -6.310 ;
        RECT 679.020 -6.320 682.020 -6.310 ;
        RECT 769.020 -6.320 772.020 -6.310 ;
        RECT 859.020 -6.320 862.020 -6.310 ;
        RECT 949.020 -6.320 952.020 -6.310 ;
        RECT 1039.020 -6.320 1042.020 -6.310 ;
        RECT 1129.020 -6.320 1132.020 -6.310 ;
        RECT 1219.020 -6.320 1222.020 -6.310 ;
        RECT 1309.020 -6.320 1312.020 -6.310 ;
        RECT 1399.020 -6.320 1402.020 -6.310 ;
        RECT 1489.020 -6.320 1492.020 -6.310 ;
        RECT 1579.020 -6.320 1582.020 -6.310 ;
        RECT 1669.020 -6.320 1672.020 -6.310 ;
        RECT 1759.020 -6.320 1762.020 -6.310 ;
        RECT 1849.020 -6.320 1852.020 -6.310 ;
        RECT 1939.020 -6.320 1942.020 -6.310 ;
        RECT 2029.020 -6.320 2032.020 -6.310 ;
        RECT 2119.020 -6.320 2122.020 -6.310 ;
        RECT 2209.020 -6.320 2212.020 -6.310 ;
        RECT 2299.020 -6.320 2302.020 -6.310 ;
        RECT 2389.020 -6.320 2392.020 -6.310 ;
        RECT 2479.020 -6.320 2482.020 -6.310 ;
        RECT 2569.020 -6.320 2572.020 -6.310 ;
        RECT 2659.020 -6.320 2662.020 -6.310 ;
        RECT 2749.020 -6.320 2752.020 -6.310 ;
        RECT 2839.020 -6.320 2842.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 49.020 -9.330 52.020 -9.320 ;
        RECT 139.020 -9.330 142.020 -9.320 ;
        RECT 229.020 -9.330 232.020 -9.320 ;
        RECT 319.020 -9.330 322.020 -9.320 ;
        RECT 409.020 -9.330 412.020 -9.320 ;
        RECT 499.020 -9.330 502.020 -9.320 ;
        RECT 589.020 -9.330 592.020 -9.320 ;
        RECT 679.020 -9.330 682.020 -9.320 ;
        RECT 769.020 -9.330 772.020 -9.320 ;
        RECT 859.020 -9.330 862.020 -9.320 ;
        RECT 949.020 -9.330 952.020 -9.320 ;
        RECT 1039.020 -9.330 1042.020 -9.320 ;
        RECT 1129.020 -9.330 1132.020 -9.320 ;
        RECT 1219.020 -9.330 1222.020 -9.320 ;
        RECT 1309.020 -9.330 1312.020 -9.320 ;
        RECT 1399.020 -9.330 1402.020 -9.320 ;
        RECT 1489.020 -9.330 1492.020 -9.320 ;
        RECT 1579.020 -9.330 1582.020 -9.320 ;
        RECT 1669.020 -9.330 1672.020 -9.320 ;
        RECT 1759.020 -9.330 1762.020 -9.320 ;
        RECT 1849.020 -9.330 1852.020 -9.320 ;
        RECT 1939.020 -9.330 1942.020 -9.320 ;
        RECT 2029.020 -9.330 2032.020 -9.320 ;
        RECT 2119.020 -9.330 2122.020 -9.320 ;
        RECT 2209.020 -9.330 2212.020 -9.320 ;
        RECT 2299.020 -9.330 2302.020 -9.320 ;
        RECT 2389.020 -9.330 2392.020 -9.320 ;
        RECT 2479.020 -9.330 2482.020 -9.320 ;
        RECT 2569.020 -9.330 2572.020 -9.320 ;
        RECT 2659.020 -9.330 2662.020 -9.320 ;
        RECT 2749.020 -9.330 2752.020 -9.320 ;
        RECT 2839.020 -9.330 2842.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 3519.700 25.020 3538.400 ;
        RECT 112.020 3519.700 115.020 3538.400 ;
        RECT 202.020 3519.700 205.020 3538.400 ;
        RECT 292.020 3519.700 295.020 3538.400 ;
        RECT 382.020 3519.700 385.020 3538.400 ;
        RECT 472.020 3519.700 475.020 3538.400 ;
        RECT 562.020 3519.700 565.020 3538.400 ;
        RECT 652.020 3519.700 655.020 3538.400 ;
        RECT 742.020 3519.700 745.020 3538.400 ;
        RECT 832.020 3519.700 835.020 3538.400 ;
        RECT 922.020 3519.700 925.020 3538.400 ;
        RECT 1012.020 3519.700 1015.020 3538.400 ;
        RECT 1102.020 3519.700 1105.020 3538.400 ;
        RECT 1192.020 3519.700 1195.020 3538.400 ;
        RECT 1282.020 3519.700 1285.020 3538.400 ;
        RECT 1372.020 3519.700 1375.020 3538.400 ;
        RECT 1462.020 3519.700 1465.020 3538.400 ;
        RECT 1552.020 3519.700 1555.020 3538.400 ;
        RECT 1642.020 3519.700 1645.020 3538.400 ;
        RECT 1732.020 3519.700 1735.020 3538.400 ;
        RECT 1822.020 3519.700 1825.020 3538.400 ;
        RECT 1912.020 3519.700 1915.020 3538.400 ;
        RECT 2002.020 3519.700 2005.020 3538.400 ;
        RECT 2092.020 3519.700 2095.020 3538.400 ;
        RECT 2182.020 3519.700 2185.020 3538.400 ;
        RECT 2272.020 3519.700 2275.020 3538.400 ;
        RECT 2362.020 3519.700 2365.020 3538.400 ;
        RECT 2452.020 3519.700 2455.020 3538.400 ;
        RECT 2542.020 3519.700 2545.020 3538.400 ;
        RECT 2632.020 3519.700 2635.020 3538.400 ;
        RECT 2722.020 3519.700 2725.020 3538.400 ;
        RECT 2812.020 3519.700 2815.020 3538.400 ;
        RECT 2902.020 3519.700 2905.020 3538.400 ;
        RECT 22.020 -18.720 25.020 0.300 ;
        RECT 112.020 -18.720 115.020 0.300 ;
        RECT 202.020 -18.720 205.020 0.300 ;
        RECT 292.020 -18.720 295.020 0.300 ;
        RECT 382.020 -18.720 385.020 0.300 ;
        RECT 472.020 -18.720 475.020 0.300 ;
        RECT 562.020 -18.720 565.020 0.300 ;
        RECT 652.020 -18.720 655.020 0.300 ;
        RECT 742.020 -18.720 745.020 0.300 ;
        RECT 832.020 -18.720 835.020 0.300 ;
        RECT 922.020 -18.720 925.020 0.300 ;
        RECT 1012.020 -18.720 1015.020 0.300 ;
        RECT 1102.020 -18.720 1105.020 0.300 ;
        RECT 1192.020 -18.720 1195.020 0.300 ;
        RECT 1282.020 -18.720 1285.020 0.300 ;
        RECT 1372.020 -18.720 1375.020 0.300 ;
        RECT 1462.020 -18.720 1465.020 0.300 ;
        RECT 1552.020 -18.720 1555.020 0.300 ;
        RECT 1642.020 -18.720 1645.020 0.300 ;
        RECT 1732.020 -18.720 1735.020 0.300 ;
        RECT 1822.020 -18.720 1825.020 0.300 ;
        RECT 1912.020 -18.720 1915.020 0.300 ;
        RECT 2002.020 -18.720 2005.020 0.300 ;
        RECT 2092.020 -18.720 2095.020 0.300 ;
        RECT 2182.020 -18.720 2185.020 0.300 ;
        RECT 2272.020 -18.720 2275.020 0.300 ;
        RECT 2362.020 -18.720 2365.020 0.300 ;
        RECT 2452.020 -18.720 2455.020 0.300 ;
        RECT 2542.020 -18.720 2545.020 0.300 ;
        RECT 2632.020 -18.720 2635.020 0.300 ;
        RECT 2722.020 -18.720 2725.020 0.300 ;
        RECT 2812.020 -18.720 2815.020 0.300 ;
        RECT 2902.020 -18.720 2905.020 0.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 112.930 3532.410 114.110 3533.590 ;
        RECT 112.930 3530.810 114.110 3531.990 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 292.930 3532.410 294.110 3533.590 ;
        RECT 292.930 3530.810 294.110 3531.990 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 472.930 3532.410 474.110 3533.590 ;
        RECT 472.930 3530.810 474.110 3531.990 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 652.930 3532.410 654.110 3533.590 ;
        RECT 652.930 3530.810 654.110 3531.990 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 832.930 3532.410 834.110 3533.590 ;
        RECT 832.930 3530.810 834.110 3531.990 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 1012.930 3532.410 1014.110 3533.590 ;
        RECT 1012.930 3530.810 1014.110 3531.990 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1192.930 3532.410 1194.110 3533.590 ;
        RECT 1192.930 3530.810 1194.110 3531.990 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1372.930 3532.410 1374.110 3533.590 ;
        RECT 1372.930 3530.810 1374.110 3531.990 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1552.930 3532.410 1554.110 3533.590 ;
        RECT 1552.930 3530.810 1554.110 3531.990 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1732.930 3532.410 1734.110 3533.590 ;
        RECT 1732.930 3530.810 1734.110 3531.990 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1912.930 3532.410 1914.110 3533.590 ;
        RECT 1912.930 3530.810 1914.110 3531.990 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2092.930 3532.410 2094.110 3533.590 ;
        RECT 2092.930 3530.810 2094.110 3531.990 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2272.930 3532.410 2274.110 3533.590 ;
        RECT 2272.930 3530.810 2274.110 3531.990 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2452.930 3532.410 2454.110 3533.590 ;
        RECT 2452.930 3530.810 2454.110 3531.990 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2632.930 3532.410 2634.110 3533.590 ;
        RECT 2632.930 3530.810 2634.110 3531.990 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2812.930 3532.410 2814.110 3533.590 ;
        RECT 2812.930 3530.810 2814.110 3531.990 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3359.090 -17.290 3360.270 ;
        RECT -18.470 3357.490 -17.290 3358.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3179.090 -17.290 3180.270 ;
        RECT -18.470 3177.490 -17.290 3178.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2999.090 -17.290 3000.270 ;
        RECT -18.470 2997.490 -17.290 2998.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2819.090 -17.290 2820.270 ;
        RECT -18.470 2817.490 -17.290 2818.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2639.090 -17.290 2640.270 ;
        RECT -18.470 2637.490 -17.290 2638.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2459.090 -17.290 2460.270 ;
        RECT -18.470 2457.490 -17.290 2458.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2279.090 -17.290 2280.270 ;
        RECT -18.470 2277.490 -17.290 2278.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2099.090 -17.290 2100.270 ;
        RECT -18.470 2097.490 -17.290 2098.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1919.090 -17.290 1920.270 ;
        RECT -18.470 1917.490 -17.290 1918.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1739.090 -17.290 1740.270 ;
        RECT -18.470 1737.490 -17.290 1738.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1559.090 -17.290 1560.270 ;
        RECT -18.470 1557.490 -17.290 1558.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1379.090 -17.290 1380.270 ;
        RECT -18.470 1377.490 -17.290 1378.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1199.090 -17.290 1200.270 ;
        RECT -18.470 1197.490 -17.290 1198.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 1019.090 -17.290 1020.270 ;
        RECT -18.470 1017.490 -17.290 1018.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 839.090 -17.290 840.270 ;
        RECT -18.470 837.490 -17.290 838.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 659.090 -17.290 660.270 ;
        RECT -18.470 657.490 -17.290 658.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 479.090 -17.290 480.270 ;
        RECT -18.470 477.490 -17.290 478.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 299.090 -17.290 300.270 ;
        RECT -18.470 297.490 -17.290 298.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 119.090 -17.290 120.270 ;
        RECT -18.470 117.490 -17.290 118.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3359.090 2938.090 3360.270 ;
        RECT 2936.910 3357.490 2938.090 3358.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3179.090 2938.090 3180.270 ;
        RECT 2936.910 3177.490 2938.090 3178.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2999.090 2938.090 3000.270 ;
        RECT 2936.910 2997.490 2938.090 2998.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2819.090 2938.090 2820.270 ;
        RECT 2936.910 2817.490 2938.090 2818.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2639.090 2938.090 2640.270 ;
        RECT 2936.910 2637.490 2938.090 2638.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2459.090 2938.090 2460.270 ;
        RECT 2936.910 2457.490 2938.090 2458.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2279.090 2938.090 2280.270 ;
        RECT 2936.910 2277.490 2938.090 2278.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2099.090 2938.090 2100.270 ;
        RECT 2936.910 2097.490 2938.090 2098.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1919.090 2938.090 1920.270 ;
        RECT 2936.910 1917.490 2938.090 1918.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1739.090 2938.090 1740.270 ;
        RECT 2936.910 1737.490 2938.090 1738.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1559.090 2938.090 1560.270 ;
        RECT 2936.910 1557.490 2938.090 1558.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1379.090 2938.090 1380.270 ;
        RECT 2936.910 1377.490 2938.090 1378.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1199.090 2938.090 1200.270 ;
        RECT 2936.910 1197.490 2938.090 1198.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 1019.090 2938.090 1020.270 ;
        RECT 2936.910 1017.490 2938.090 1018.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 839.090 2938.090 840.270 ;
        RECT 2936.910 837.490 2938.090 838.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 659.090 2938.090 660.270 ;
        RECT 2936.910 657.490 2938.090 658.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 479.090 2938.090 480.270 ;
        RECT 2936.910 477.490 2938.090 478.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 299.090 2938.090 300.270 ;
        RECT 2936.910 297.490 2938.090 298.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 119.090 2938.090 120.270 ;
        RECT 2936.910 117.490 2938.090 118.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 112.930 -12.310 114.110 -11.130 ;
        RECT 112.930 -13.910 114.110 -12.730 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 292.930 -12.310 294.110 -11.130 ;
        RECT 292.930 -13.910 294.110 -12.730 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 472.930 -12.310 474.110 -11.130 ;
        RECT 472.930 -13.910 474.110 -12.730 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 652.930 -12.310 654.110 -11.130 ;
        RECT 652.930 -13.910 654.110 -12.730 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 832.930 -12.310 834.110 -11.130 ;
        RECT 832.930 -13.910 834.110 -12.730 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1012.930 -12.310 1014.110 -11.130 ;
        RECT 1012.930 -13.910 1014.110 -12.730 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1192.930 -12.310 1194.110 -11.130 ;
        RECT 1192.930 -13.910 1194.110 -12.730 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1372.930 -12.310 1374.110 -11.130 ;
        RECT 1372.930 -13.910 1374.110 -12.730 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1552.930 -12.310 1554.110 -11.130 ;
        RECT 1552.930 -13.910 1554.110 -12.730 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1732.930 -12.310 1734.110 -11.130 ;
        RECT 1732.930 -13.910 1734.110 -12.730 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 1912.930 -12.310 1914.110 -11.130 ;
        RECT 1912.930 -13.910 1914.110 -12.730 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2092.930 -12.310 2094.110 -11.130 ;
        RECT 2092.930 -13.910 2094.110 -12.730 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2272.930 -12.310 2274.110 -11.130 ;
        RECT 2272.930 -13.910 2274.110 -12.730 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2452.930 -12.310 2454.110 -11.130 ;
        RECT 2452.930 -13.910 2454.110 -12.730 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2632.930 -12.310 2634.110 -11.130 ;
        RECT 2632.930 -13.910 2634.110 -12.730 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2812.930 -12.310 2814.110 -11.130 ;
        RECT 2812.930 -13.910 2814.110 -12.730 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 112.020 3533.700 115.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 292.020 3533.700 295.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 472.020 3533.700 475.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 652.020 3533.700 655.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 832.020 3533.700 835.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1012.020 3533.700 1015.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1192.020 3533.700 1195.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1372.020 3533.700 1375.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1552.020 3533.700 1555.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1732.020 3533.700 1735.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 1912.020 3533.700 1915.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2092.020 3533.700 2095.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2272.020 3533.700 2275.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2452.020 3533.700 2455.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2632.020 3533.700 2635.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2812.020 3533.700 2815.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 112.020 3530.690 115.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 292.020 3530.690 295.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 472.020 3530.690 475.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 652.020 3530.690 655.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 832.020 3530.690 835.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1012.020 3530.690 1015.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1192.020 3530.690 1195.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1372.020 3530.690 1375.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1552.020 3530.690 1555.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1732.020 3530.690 1735.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 1912.020 3530.690 1915.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2092.020 3530.690 2095.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2272.020 3530.690 2275.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2452.020 3530.690 2455.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2632.020 3530.690 2635.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2812.020 3530.690 2815.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 0.300 3450.380 ;
        RECT 2919.700 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3360.380 -16.380 3360.390 ;
        RECT 2936.000 3360.380 2939.000 3360.390 ;
        RECT -24.080 3357.380 0.300 3360.380 ;
        RECT 2919.700 3357.380 2943.700 3360.380 ;
        RECT -19.380 3357.370 -16.380 3357.380 ;
        RECT 2936.000 3357.370 2939.000 3357.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 0.300 3270.380 ;
        RECT 2919.700 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3180.380 -16.380 3180.390 ;
        RECT 2936.000 3180.380 2939.000 3180.390 ;
        RECT -24.080 3177.380 0.300 3180.380 ;
        RECT 2919.700 3177.380 2943.700 3180.380 ;
        RECT -19.380 3177.370 -16.380 3177.380 ;
        RECT 2936.000 3177.370 2939.000 3177.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 0.300 3090.380 ;
        RECT 2919.700 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 3000.380 -16.380 3000.390 ;
        RECT 2936.000 3000.380 2939.000 3000.390 ;
        RECT -24.080 2997.380 0.300 3000.380 ;
        RECT 2919.700 2997.380 2943.700 3000.380 ;
        RECT -19.380 2997.370 -16.380 2997.380 ;
        RECT 2936.000 2997.370 2939.000 2997.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 0.300 2910.380 ;
        RECT 2919.700 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2820.380 -16.380 2820.390 ;
        RECT 2936.000 2820.380 2939.000 2820.390 ;
        RECT -24.080 2817.380 0.300 2820.380 ;
        RECT 2919.700 2817.380 2943.700 2820.380 ;
        RECT -19.380 2817.370 -16.380 2817.380 ;
        RECT 2936.000 2817.370 2939.000 2817.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 0.300 2730.380 ;
        RECT 2919.700 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2640.380 -16.380 2640.390 ;
        RECT 2936.000 2640.380 2939.000 2640.390 ;
        RECT -24.080 2637.380 0.300 2640.380 ;
        RECT 2919.700 2637.380 2943.700 2640.380 ;
        RECT -19.380 2637.370 -16.380 2637.380 ;
        RECT 2936.000 2637.370 2939.000 2637.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 0.300 2550.380 ;
        RECT 2919.700 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2460.380 -16.380 2460.390 ;
        RECT 2936.000 2460.380 2939.000 2460.390 ;
        RECT -24.080 2457.380 0.300 2460.380 ;
        RECT 2919.700 2457.380 2943.700 2460.380 ;
        RECT -19.380 2457.370 -16.380 2457.380 ;
        RECT 2936.000 2457.370 2939.000 2457.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 0.300 2370.380 ;
        RECT 2919.700 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2280.380 -16.380 2280.390 ;
        RECT 2936.000 2280.380 2939.000 2280.390 ;
        RECT -24.080 2277.380 0.300 2280.380 ;
        RECT 2919.700 2277.380 2943.700 2280.380 ;
        RECT -19.380 2277.370 -16.380 2277.380 ;
        RECT 2936.000 2277.370 2939.000 2277.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 0.300 2190.380 ;
        RECT 2919.700 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2100.380 -16.380 2100.390 ;
        RECT 2936.000 2100.380 2939.000 2100.390 ;
        RECT -24.080 2097.380 0.300 2100.380 ;
        RECT 2919.700 2097.380 2943.700 2100.380 ;
        RECT -19.380 2097.370 -16.380 2097.380 ;
        RECT 2936.000 2097.370 2939.000 2097.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 0.300 2010.380 ;
        RECT 2919.700 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1920.380 -16.380 1920.390 ;
        RECT 2936.000 1920.380 2939.000 1920.390 ;
        RECT -24.080 1917.380 0.300 1920.380 ;
        RECT 2919.700 1917.380 2943.700 1920.380 ;
        RECT -19.380 1917.370 -16.380 1917.380 ;
        RECT 2936.000 1917.370 2939.000 1917.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 0.300 1830.380 ;
        RECT 2919.700 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1740.380 -16.380 1740.390 ;
        RECT 2936.000 1740.380 2939.000 1740.390 ;
        RECT -24.080 1737.380 0.300 1740.380 ;
        RECT 2919.700 1737.380 2943.700 1740.380 ;
        RECT -19.380 1737.370 -16.380 1737.380 ;
        RECT 2936.000 1737.370 2939.000 1737.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 0.300 1650.380 ;
        RECT 2919.700 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1560.380 -16.380 1560.390 ;
        RECT 2936.000 1560.380 2939.000 1560.390 ;
        RECT -24.080 1557.380 0.300 1560.380 ;
        RECT 2919.700 1557.380 2943.700 1560.380 ;
        RECT -19.380 1557.370 -16.380 1557.380 ;
        RECT 2936.000 1557.370 2939.000 1557.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 0.300 1470.380 ;
        RECT 2919.700 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1380.380 -16.380 1380.390 ;
        RECT 2936.000 1380.380 2939.000 1380.390 ;
        RECT -24.080 1377.380 0.300 1380.380 ;
        RECT 2919.700 1377.380 2943.700 1380.380 ;
        RECT -19.380 1377.370 -16.380 1377.380 ;
        RECT 2936.000 1377.370 2939.000 1377.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 0.300 1290.380 ;
        RECT 2919.700 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1200.380 -16.380 1200.390 ;
        RECT 2936.000 1200.380 2939.000 1200.390 ;
        RECT -24.080 1197.380 0.300 1200.380 ;
        RECT 2919.700 1197.380 2943.700 1200.380 ;
        RECT -19.380 1197.370 -16.380 1197.380 ;
        RECT 2936.000 1197.370 2939.000 1197.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 0.300 1110.380 ;
        RECT 2919.700 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 1020.380 -16.380 1020.390 ;
        RECT 2936.000 1020.380 2939.000 1020.390 ;
        RECT -24.080 1017.380 0.300 1020.380 ;
        RECT 2919.700 1017.380 2943.700 1020.380 ;
        RECT -19.380 1017.370 -16.380 1017.380 ;
        RECT 2936.000 1017.370 2939.000 1017.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 0.300 930.380 ;
        RECT 2919.700 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 840.380 -16.380 840.390 ;
        RECT 2936.000 840.380 2939.000 840.390 ;
        RECT -24.080 837.380 0.300 840.380 ;
        RECT 2919.700 837.380 2943.700 840.380 ;
        RECT -19.380 837.370 -16.380 837.380 ;
        RECT 2936.000 837.370 2939.000 837.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 0.300 750.380 ;
        RECT 2919.700 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 660.380 -16.380 660.390 ;
        RECT 2936.000 660.380 2939.000 660.390 ;
        RECT -24.080 657.380 0.300 660.380 ;
        RECT 2919.700 657.380 2943.700 660.380 ;
        RECT -19.380 657.370 -16.380 657.380 ;
        RECT 2936.000 657.370 2939.000 657.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 0.300 570.380 ;
        RECT 2919.700 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 480.380 -16.380 480.390 ;
        RECT 2936.000 480.380 2939.000 480.390 ;
        RECT -24.080 477.380 0.300 480.380 ;
        RECT 2919.700 477.380 2943.700 480.380 ;
        RECT -19.380 477.370 -16.380 477.380 ;
        RECT 2936.000 477.370 2939.000 477.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 0.300 390.380 ;
        RECT 2919.700 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 300.380 -16.380 300.390 ;
        RECT 2936.000 300.380 2939.000 300.390 ;
        RECT -24.080 297.380 0.300 300.380 ;
        RECT 2919.700 297.380 2943.700 300.380 ;
        RECT -19.380 297.370 -16.380 297.380 ;
        RECT 2936.000 297.370 2939.000 297.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 0.300 210.380 ;
        RECT 2919.700 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 120.380 -16.380 120.390 ;
        RECT 2936.000 120.380 2939.000 120.390 ;
        RECT -24.080 117.380 0.300 120.380 ;
        RECT 2919.700 117.380 2943.700 120.380 ;
        RECT -19.380 117.370 -16.380 117.380 ;
        RECT 2936.000 117.370 2939.000 117.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 0.300 30.380 ;
        RECT 2919.700 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 112.020 -11.020 115.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 292.020 -11.020 295.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 472.020 -11.020 475.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 652.020 -11.020 655.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 832.020 -11.020 835.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1012.020 -11.020 1015.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1192.020 -11.020 1195.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1372.020 -11.020 1375.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1552.020 -11.020 1555.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1732.020 -11.020 1735.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 1912.020 -11.020 1915.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2092.020 -11.020 2095.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2272.020 -11.020 2275.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2452.020 -11.020 2455.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2632.020 -11.020 2635.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2812.020 -11.020 2815.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 112.020 -14.030 115.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 292.020 -14.030 295.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 472.020 -14.030 475.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 652.020 -14.030 655.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 832.020 -14.030 835.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1012.020 -14.030 1015.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1192.020 -14.030 1195.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1372.020 -14.030 1375.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1552.020 -14.030 1555.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1732.020 -14.030 1735.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 1912.020 -14.030 1915.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2092.020 -14.030 2095.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2272.020 -14.030 2275.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2452.020 -14.030 2455.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2632.020 -14.030 2635.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2812.020 -14.030 2815.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 67.020 3519.700 70.020 3538.400 ;
        RECT 157.020 3519.700 160.020 3538.400 ;
        RECT 247.020 3519.700 250.020 3538.400 ;
        RECT 337.020 3519.700 340.020 3538.400 ;
        RECT 427.020 3519.700 430.020 3538.400 ;
        RECT 517.020 3519.700 520.020 3538.400 ;
        RECT 607.020 3519.700 610.020 3538.400 ;
        RECT 697.020 3519.700 700.020 3538.400 ;
        RECT 787.020 3519.700 790.020 3538.400 ;
        RECT 877.020 3519.700 880.020 3538.400 ;
        RECT 967.020 3519.700 970.020 3538.400 ;
        RECT 1057.020 3519.700 1060.020 3538.400 ;
        RECT 1147.020 3519.700 1150.020 3538.400 ;
        RECT 1237.020 3519.700 1240.020 3538.400 ;
        RECT 1327.020 3519.700 1330.020 3538.400 ;
        RECT 1417.020 3519.700 1420.020 3538.400 ;
        RECT 1507.020 3519.700 1510.020 3538.400 ;
        RECT 1597.020 3519.700 1600.020 3538.400 ;
        RECT 1687.020 3519.700 1690.020 3538.400 ;
        RECT 1777.020 3519.700 1780.020 3538.400 ;
        RECT 1867.020 3519.700 1870.020 3538.400 ;
        RECT 1957.020 3519.700 1960.020 3538.400 ;
        RECT 2047.020 3519.700 2050.020 3538.400 ;
        RECT 2137.020 3519.700 2140.020 3538.400 ;
        RECT 2227.020 3519.700 2230.020 3538.400 ;
        RECT 2317.020 3519.700 2320.020 3538.400 ;
        RECT 2407.020 3519.700 2410.020 3538.400 ;
        RECT 2497.020 3519.700 2500.020 3538.400 ;
        RECT 2587.020 3519.700 2590.020 3538.400 ;
        RECT 2677.020 3519.700 2680.020 3538.400 ;
        RECT 2767.020 3519.700 2770.020 3538.400 ;
        RECT 2857.020 3519.700 2860.020 3538.400 ;
        RECT 67.020 -18.720 70.020 0.300 ;
        RECT 157.020 -18.720 160.020 0.300 ;
        RECT 247.020 -18.720 250.020 0.300 ;
        RECT 337.020 -18.720 340.020 0.300 ;
        RECT 427.020 -18.720 430.020 0.300 ;
        RECT 517.020 -18.720 520.020 0.300 ;
        RECT 607.020 -18.720 610.020 0.300 ;
        RECT 697.020 -18.720 700.020 0.300 ;
        RECT 787.020 -18.720 790.020 0.300 ;
        RECT 877.020 -18.720 880.020 0.300 ;
        RECT 967.020 -18.720 970.020 0.300 ;
        RECT 1057.020 -18.720 1060.020 0.300 ;
        RECT 1147.020 -18.720 1150.020 0.300 ;
        RECT 1237.020 -18.720 1240.020 0.300 ;
        RECT 1327.020 -18.720 1330.020 0.300 ;
        RECT 1417.020 -18.720 1420.020 0.300 ;
        RECT 1507.020 -18.720 1510.020 0.300 ;
        RECT 1597.020 -18.720 1600.020 0.300 ;
        RECT 1687.020 -18.720 1690.020 0.300 ;
        RECT 1777.020 -18.720 1780.020 0.300 ;
        RECT 1867.020 -18.720 1870.020 0.300 ;
        RECT 1957.020 -18.720 1960.020 0.300 ;
        RECT 2047.020 -18.720 2050.020 0.300 ;
        RECT 2137.020 -18.720 2140.020 0.300 ;
        RECT 2227.020 -18.720 2230.020 0.300 ;
        RECT 2317.020 -18.720 2320.020 0.300 ;
        RECT 2407.020 -18.720 2410.020 0.300 ;
        RECT 2497.020 -18.720 2500.020 0.300 ;
        RECT 2587.020 -18.720 2590.020 0.300 ;
        RECT 2677.020 -18.720 2680.020 0.300 ;
        RECT 2767.020 -18.720 2770.020 0.300 ;
        RECT 2857.020 -18.720 2860.020 0.300 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 67.930 3537.110 69.110 3538.290 ;
        RECT 67.930 3535.510 69.110 3536.690 ;
        RECT 157.930 3537.110 159.110 3538.290 ;
        RECT 157.930 3535.510 159.110 3536.690 ;
        RECT 247.930 3537.110 249.110 3538.290 ;
        RECT 247.930 3535.510 249.110 3536.690 ;
        RECT 337.930 3537.110 339.110 3538.290 ;
        RECT 337.930 3535.510 339.110 3536.690 ;
        RECT 427.930 3537.110 429.110 3538.290 ;
        RECT 427.930 3535.510 429.110 3536.690 ;
        RECT 517.930 3537.110 519.110 3538.290 ;
        RECT 517.930 3535.510 519.110 3536.690 ;
        RECT 607.930 3537.110 609.110 3538.290 ;
        RECT 607.930 3535.510 609.110 3536.690 ;
        RECT 697.930 3537.110 699.110 3538.290 ;
        RECT 697.930 3535.510 699.110 3536.690 ;
        RECT 787.930 3537.110 789.110 3538.290 ;
        RECT 787.930 3535.510 789.110 3536.690 ;
        RECT 877.930 3537.110 879.110 3538.290 ;
        RECT 877.930 3535.510 879.110 3536.690 ;
        RECT 967.930 3537.110 969.110 3538.290 ;
        RECT 967.930 3535.510 969.110 3536.690 ;
        RECT 1057.930 3537.110 1059.110 3538.290 ;
        RECT 1057.930 3535.510 1059.110 3536.690 ;
        RECT 1147.930 3537.110 1149.110 3538.290 ;
        RECT 1147.930 3535.510 1149.110 3536.690 ;
        RECT 1237.930 3537.110 1239.110 3538.290 ;
        RECT 1237.930 3535.510 1239.110 3536.690 ;
        RECT 1327.930 3537.110 1329.110 3538.290 ;
        RECT 1327.930 3535.510 1329.110 3536.690 ;
        RECT 1417.930 3537.110 1419.110 3538.290 ;
        RECT 1417.930 3535.510 1419.110 3536.690 ;
        RECT 1507.930 3537.110 1509.110 3538.290 ;
        RECT 1507.930 3535.510 1509.110 3536.690 ;
        RECT 1597.930 3537.110 1599.110 3538.290 ;
        RECT 1597.930 3535.510 1599.110 3536.690 ;
        RECT 1687.930 3537.110 1689.110 3538.290 ;
        RECT 1687.930 3535.510 1689.110 3536.690 ;
        RECT 1777.930 3537.110 1779.110 3538.290 ;
        RECT 1777.930 3535.510 1779.110 3536.690 ;
        RECT 1867.930 3537.110 1869.110 3538.290 ;
        RECT 1867.930 3535.510 1869.110 3536.690 ;
        RECT 1957.930 3537.110 1959.110 3538.290 ;
        RECT 1957.930 3535.510 1959.110 3536.690 ;
        RECT 2047.930 3537.110 2049.110 3538.290 ;
        RECT 2047.930 3535.510 2049.110 3536.690 ;
        RECT 2137.930 3537.110 2139.110 3538.290 ;
        RECT 2137.930 3535.510 2139.110 3536.690 ;
        RECT 2227.930 3537.110 2229.110 3538.290 ;
        RECT 2227.930 3535.510 2229.110 3536.690 ;
        RECT 2317.930 3537.110 2319.110 3538.290 ;
        RECT 2317.930 3535.510 2319.110 3536.690 ;
        RECT 2407.930 3537.110 2409.110 3538.290 ;
        RECT 2407.930 3535.510 2409.110 3536.690 ;
        RECT 2497.930 3537.110 2499.110 3538.290 ;
        RECT 2497.930 3535.510 2499.110 3536.690 ;
        RECT 2587.930 3537.110 2589.110 3538.290 ;
        RECT 2587.930 3535.510 2589.110 3536.690 ;
        RECT 2677.930 3537.110 2679.110 3538.290 ;
        RECT 2677.930 3535.510 2679.110 3536.690 ;
        RECT 2767.930 3537.110 2769.110 3538.290 ;
        RECT 2767.930 3535.510 2769.110 3536.690 ;
        RECT 2857.930 3537.110 2859.110 3538.290 ;
        RECT 2857.930 3535.510 2859.110 3536.690 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT -23.170 3494.090 -21.990 3495.270 ;
        RECT -23.170 3492.490 -21.990 3493.670 ;
        RECT -23.170 3404.090 -21.990 3405.270 ;
        RECT -23.170 3402.490 -21.990 3403.670 ;
        RECT -23.170 3314.090 -21.990 3315.270 ;
        RECT -23.170 3312.490 -21.990 3313.670 ;
        RECT -23.170 3224.090 -21.990 3225.270 ;
        RECT -23.170 3222.490 -21.990 3223.670 ;
        RECT -23.170 3134.090 -21.990 3135.270 ;
        RECT -23.170 3132.490 -21.990 3133.670 ;
        RECT -23.170 3044.090 -21.990 3045.270 ;
        RECT -23.170 3042.490 -21.990 3043.670 ;
        RECT -23.170 2954.090 -21.990 2955.270 ;
        RECT -23.170 2952.490 -21.990 2953.670 ;
        RECT -23.170 2864.090 -21.990 2865.270 ;
        RECT -23.170 2862.490 -21.990 2863.670 ;
        RECT -23.170 2774.090 -21.990 2775.270 ;
        RECT -23.170 2772.490 -21.990 2773.670 ;
        RECT -23.170 2684.090 -21.990 2685.270 ;
        RECT -23.170 2682.490 -21.990 2683.670 ;
        RECT -23.170 2594.090 -21.990 2595.270 ;
        RECT -23.170 2592.490 -21.990 2593.670 ;
        RECT -23.170 2504.090 -21.990 2505.270 ;
        RECT -23.170 2502.490 -21.990 2503.670 ;
        RECT -23.170 2414.090 -21.990 2415.270 ;
        RECT -23.170 2412.490 -21.990 2413.670 ;
        RECT -23.170 2324.090 -21.990 2325.270 ;
        RECT -23.170 2322.490 -21.990 2323.670 ;
        RECT -23.170 2234.090 -21.990 2235.270 ;
        RECT -23.170 2232.490 -21.990 2233.670 ;
        RECT -23.170 2144.090 -21.990 2145.270 ;
        RECT -23.170 2142.490 -21.990 2143.670 ;
        RECT -23.170 2054.090 -21.990 2055.270 ;
        RECT -23.170 2052.490 -21.990 2053.670 ;
        RECT -23.170 1964.090 -21.990 1965.270 ;
        RECT -23.170 1962.490 -21.990 1963.670 ;
        RECT -23.170 1874.090 -21.990 1875.270 ;
        RECT -23.170 1872.490 -21.990 1873.670 ;
        RECT -23.170 1784.090 -21.990 1785.270 ;
        RECT -23.170 1782.490 -21.990 1783.670 ;
        RECT -23.170 1694.090 -21.990 1695.270 ;
        RECT -23.170 1692.490 -21.990 1693.670 ;
        RECT -23.170 1604.090 -21.990 1605.270 ;
        RECT -23.170 1602.490 -21.990 1603.670 ;
        RECT -23.170 1514.090 -21.990 1515.270 ;
        RECT -23.170 1512.490 -21.990 1513.670 ;
        RECT -23.170 1424.090 -21.990 1425.270 ;
        RECT -23.170 1422.490 -21.990 1423.670 ;
        RECT -23.170 1334.090 -21.990 1335.270 ;
        RECT -23.170 1332.490 -21.990 1333.670 ;
        RECT -23.170 1244.090 -21.990 1245.270 ;
        RECT -23.170 1242.490 -21.990 1243.670 ;
        RECT -23.170 1154.090 -21.990 1155.270 ;
        RECT -23.170 1152.490 -21.990 1153.670 ;
        RECT -23.170 1064.090 -21.990 1065.270 ;
        RECT -23.170 1062.490 -21.990 1063.670 ;
        RECT -23.170 974.090 -21.990 975.270 ;
        RECT -23.170 972.490 -21.990 973.670 ;
        RECT -23.170 884.090 -21.990 885.270 ;
        RECT -23.170 882.490 -21.990 883.670 ;
        RECT -23.170 794.090 -21.990 795.270 ;
        RECT -23.170 792.490 -21.990 793.670 ;
        RECT -23.170 704.090 -21.990 705.270 ;
        RECT -23.170 702.490 -21.990 703.670 ;
        RECT -23.170 614.090 -21.990 615.270 ;
        RECT -23.170 612.490 -21.990 613.670 ;
        RECT -23.170 524.090 -21.990 525.270 ;
        RECT -23.170 522.490 -21.990 523.670 ;
        RECT -23.170 434.090 -21.990 435.270 ;
        RECT -23.170 432.490 -21.990 433.670 ;
        RECT -23.170 344.090 -21.990 345.270 ;
        RECT -23.170 342.490 -21.990 343.670 ;
        RECT -23.170 254.090 -21.990 255.270 ;
        RECT -23.170 252.490 -21.990 253.670 ;
        RECT -23.170 164.090 -21.990 165.270 ;
        RECT -23.170 162.490 -21.990 163.670 ;
        RECT -23.170 74.090 -21.990 75.270 ;
        RECT -23.170 72.490 -21.990 73.670 ;
        RECT 2941.610 3494.090 2942.790 3495.270 ;
        RECT 2941.610 3492.490 2942.790 3493.670 ;
        RECT 2941.610 3404.090 2942.790 3405.270 ;
        RECT 2941.610 3402.490 2942.790 3403.670 ;
        RECT 2941.610 3314.090 2942.790 3315.270 ;
        RECT 2941.610 3312.490 2942.790 3313.670 ;
        RECT 2941.610 3224.090 2942.790 3225.270 ;
        RECT 2941.610 3222.490 2942.790 3223.670 ;
        RECT 2941.610 3134.090 2942.790 3135.270 ;
        RECT 2941.610 3132.490 2942.790 3133.670 ;
        RECT 2941.610 3044.090 2942.790 3045.270 ;
        RECT 2941.610 3042.490 2942.790 3043.670 ;
        RECT 2941.610 2954.090 2942.790 2955.270 ;
        RECT 2941.610 2952.490 2942.790 2953.670 ;
        RECT 2941.610 2864.090 2942.790 2865.270 ;
        RECT 2941.610 2862.490 2942.790 2863.670 ;
        RECT 2941.610 2774.090 2942.790 2775.270 ;
        RECT 2941.610 2772.490 2942.790 2773.670 ;
        RECT 2941.610 2684.090 2942.790 2685.270 ;
        RECT 2941.610 2682.490 2942.790 2683.670 ;
        RECT 2941.610 2594.090 2942.790 2595.270 ;
        RECT 2941.610 2592.490 2942.790 2593.670 ;
        RECT 2941.610 2504.090 2942.790 2505.270 ;
        RECT 2941.610 2502.490 2942.790 2503.670 ;
        RECT 2941.610 2414.090 2942.790 2415.270 ;
        RECT 2941.610 2412.490 2942.790 2413.670 ;
        RECT 2941.610 2324.090 2942.790 2325.270 ;
        RECT 2941.610 2322.490 2942.790 2323.670 ;
        RECT 2941.610 2234.090 2942.790 2235.270 ;
        RECT 2941.610 2232.490 2942.790 2233.670 ;
        RECT 2941.610 2144.090 2942.790 2145.270 ;
        RECT 2941.610 2142.490 2942.790 2143.670 ;
        RECT 2941.610 2054.090 2942.790 2055.270 ;
        RECT 2941.610 2052.490 2942.790 2053.670 ;
        RECT 2941.610 1964.090 2942.790 1965.270 ;
        RECT 2941.610 1962.490 2942.790 1963.670 ;
        RECT 2941.610 1874.090 2942.790 1875.270 ;
        RECT 2941.610 1872.490 2942.790 1873.670 ;
        RECT 2941.610 1784.090 2942.790 1785.270 ;
        RECT 2941.610 1782.490 2942.790 1783.670 ;
        RECT 2941.610 1694.090 2942.790 1695.270 ;
        RECT 2941.610 1692.490 2942.790 1693.670 ;
        RECT 2941.610 1604.090 2942.790 1605.270 ;
        RECT 2941.610 1602.490 2942.790 1603.670 ;
        RECT 2941.610 1514.090 2942.790 1515.270 ;
        RECT 2941.610 1512.490 2942.790 1513.670 ;
        RECT 2941.610 1424.090 2942.790 1425.270 ;
        RECT 2941.610 1422.490 2942.790 1423.670 ;
        RECT 2941.610 1334.090 2942.790 1335.270 ;
        RECT 2941.610 1332.490 2942.790 1333.670 ;
        RECT 2941.610 1244.090 2942.790 1245.270 ;
        RECT 2941.610 1242.490 2942.790 1243.670 ;
        RECT 2941.610 1154.090 2942.790 1155.270 ;
        RECT 2941.610 1152.490 2942.790 1153.670 ;
        RECT 2941.610 1064.090 2942.790 1065.270 ;
        RECT 2941.610 1062.490 2942.790 1063.670 ;
        RECT 2941.610 974.090 2942.790 975.270 ;
        RECT 2941.610 972.490 2942.790 973.670 ;
        RECT 2941.610 884.090 2942.790 885.270 ;
        RECT 2941.610 882.490 2942.790 883.670 ;
        RECT 2941.610 794.090 2942.790 795.270 ;
        RECT 2941.610 792.490 2942.790 793.670 ;
        RECT 2941.610 704.090 2942.790 705.270 ;
        RECT 2941.610 702.490 2942.790 703.670 ;
        RECT 2941.610 614.090 2942.790 615.270 ;
        RECT 2941.610 612.490 2942.790 613.670 ;
        RECT 2941.610 524.090 2942.790 525.270 ;
        RECT 2941.610 522.490 2942.790 523.670 ;
        RECT 2941.610 434.090 2942.790 435.270 ;
        RECT 2941.610 432.490 2942.790 433.670 ;
        RECT 2941.610 344.090 2942.790 345.270 ;
        RECT 2941.610 342.490 2942.790 343.670 ;
        RECT 2941.610 254.090 2942.790 255.270 ;
        RECT 2941.610 252.490 2942.790 253.670 ;
        RECT 2941.610 164.090 2942.790 165.270 ;
        RECT 2941.610 162.490 2942.790 163.670 ;
        RECT 2941.610 74.090 2942.790 75.270 ;
        RECT 2941.610 72.490 2942.790 73.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 67.930 -17.010 69.110 -15.830 ;
        RECT 67.930 -18.610 69.110 -17.430 ;
        RECT 157.930 -17.010 159.110 -15.830 ;
        RECT 157.930 -18.610 159.110 -17.430 ;
        RECT 247.930 -17.010 249.110 -15.830 ;
        RECT 247.930 -18.610 249.110 -17.430 ;
        RECT 337.930 -17.010 339.110 -15.830 ;
        RECT 337.930 -18.610 339.110 -17.430 ;
        RECT 427.930 -17.010 429.110 -15.830 ;
        RECT 427.930 -18.610 429.110 -17.430 ;
        RECT 517.930 -17.010 519.110 -15.830 ;
        RECT 517.930 -18.610 519.110 -17.430 ;
        RECT 607.930 -17.010 609.110 -15.830 ;
        RECT 607.930 -18.610 609.110 -17.430 ;
        RECT 697.930 -17.010 699.110 -15.830 ;
        RECT 697.930 -18.610 699.110 -17.430 ;
        RECT 787.930 -17.010 789.110 -15.830 ;
        RECT 787.930 -18.610 789.110 -17.430 ;
        RECT 877.930 -17.010 879.110 -15.830 ;
        RECT 877.930 -18.610 879.110 -17.430 ;
        RECT 967.930 -17.010 969.110 -15.830 ;
        RECT 967.930 -18.610 969.110 -17.430 ;
        RECT 1057.930 -17.010 1059.110 -15.830 ;
        RECT 1057.930 -18.610 1059.110 -17.430 ;
        RECT 1147.930 -17.010 1149.110 -15.830 ;
        RECT 1147.930 -18.610 1149.110 -17.430 ;
        RECT 1237.930 -17.010 1239.110 -15.830 ;
        RECT 1237.930 -18.610 1239.110 -17.430 ;
        RECT 1327.930 -17.010 1329.110 -15.830 ;
        RECT 1327.930 -18.610 1329.110 -17.430 ;
        RECT 1417.930 -17.010 1419.110 -15.830 ;
        RECT 1417.930 -18.610 1419.110 -17.430 ;
        RECT 1507.930 -17.010 1509.110 -15.830 ;
        RECT 1507.930 -18.610 1509.110 -17.430 ;
        RECT 1597.930 -17.010 1599.110 -15.830 ;
        RECT 1597.930 -18.610 1599.110 -17.430 ;
        RECT 1687.930 -17.010 1689.110 -15.830 ;
        RECT 1687.930 -18.610 1689.110 -17.430 ;
        RECT 1777.930 -17.010 1779.110 -15.830 ;
        RECT 1777.930 -18.610 1779.110 -17.430 ;
        RECT 1867.930 -17.010 1869.110 -15.830 ;
        RECT 1867.930 -18.610 1869.110 -17.430 ;
        RECT 1957.930 -17.010 1959.110 -15.830 ;
        RECT 1957.930 -18.610 1959.110 -17.430 ;
        RECT 2047.930 -17.010 2049.110 -15.830 ;
        RECT 2047.930 -18.610 2049.110 -17.430 ;
        RECT 2137.930 -17.010 2139.110 -15.830 ;
        RECT 2137.930 -18.610 2139.110 -17.430 ;
        RECT 2227.930 -17.010 2229.110 -15.830 ;
        RECT 2227.930 -18.610 2229.110 -17.430 ;
        RECT 2317.930 -17.010 2319.110 -15.830 ;
        RECT 2317.930 -18.610 2319.110 -17.430 ;
        RECT 2407.930 -17.010 2409.110 -15.830 ;
        RECT 2407.930 -18.610 2409.110 -17.430 ;
        RECT 2497.930 -17.010 2499.110 -15.830 ;
        RECT 2497.930 -18.610 2499.110 -17.430 ;
        RECT 2587.930 -17.010 2589.110 -15.830 ;
        RECT 2587.930 -18.610 2589.110 -17.430 ;
        RECT 2677.930 -17.010 2679.110 -15.830 ;
        RECT 2677.930 -18.610 2679.110 -17.430 ;
        RECT 2767.930 -17.010 2769.110 -15.830 ;
        RECT 2767.930 -18.610 2769.110 -17.430 ;
        RECT 2857.930 -17.010 2859.110 -15.830 ;
        RECT 2857.930 -18.610 2859.110 -17.430 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 67.020 3538.400 70.020 3538.410 ;
        RECT 157.020 3538.400 160.020 3538.410 ;
        RECT 247.020 3538.400 250.020 3538.410 ;
        RECT 337.020 3538.400 340.020 3538.410 ;
        RECT 427.020 3538.400 430.020 3538.410 ;
        RECT 517.020 3538.400 520.020 3538.410 ;
        RECT 607.020 3538.400 610.020 3538.410 ;
        RECT 697.020 3538.400 700.020 3538.410 ;
        RECT 787.020 3538.400 790.020 3538.410 ;
        RECT 877.020 3538.400 880.020 3538.410 ;
        RECT 967.020 3538.400 970.020 3538.410 ;
        RECT 1057.020 3538.400 1060.020 3538.410 ;
        RECT 1147.020 3538.400 1150.020 3538.410 ;
        RECT 1237.020 3538.400 1240.020 3538.410 ;
        RECT 1327.020 3538.400 1330.020 3538.410 ;
        RECT 1417.020 3538.400 1420.020 3538.410 ;
        RECT 1507.020 3538.400 1510.020 3538.410 ;
        RECT 1597.020 3538.400 1600.020 3538.410 ;
        RECT 1687.020 3538.400 1690.020 3538.410 ;
        RECT 1777.020 3538.400 1780.020 3538.410 ;
        RECT 1867.020 3538.400 1870.020 3538.410 ;
        RECT 1957.020 3538.400 1960.020 3538.410 ;
        RECT 2047.020 3538.400 2050.020 3538.410 ;
        RECT 2137.020 3538.400 2140.020 3538.410 ;
        RECT 2227.020 3538.400 2230.020 3538.410 ;
        RECT 2317.020 3538.400 2320.020 3538.410 ;
        RECT 2407.020 3538.400 2410.020 3538.410 ;
        RECT 2497.020 3538.400 2500.020 3538.410 ;
        RECT 2587.020 3538.400 2590.020 3538.410 ;
        RECT 2677.020 3538.400 2680.020 3538.410 ;
        RECT 2767.020 3538.400 2770.020 3538.410 ;
        RECT 2857.020 3538.400 2860.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 67.020 3535.390 70.020 3535.400 ;
        RECT 157.020 3535.390 160.020 3535.400 ;
        RECT 247.020 3535.390 250.020 3535.400 ;
        RECT 337.020 3535.390 340.020 3535.400 ;
        RECT 427.020 3535.390 430.020 3535.400 ;
        RECT 517.020 3535.390 520.020 3535.400 ;
        RECT 607.020 3535.390 610.020 3535.400 ;
        RECT 697.020 3535.390 700.020 3535.400 ;
        RECT 787.020 3535.390 790.020 3535.400 ;
        RECT 877.020 3535.390 880.020 3535.400 ;
        RECT 967.020 3535.390 970.020 3535.400 ;
        RECT 1057.020 3535.390 1060.020 3535.400 ;
        RECT 1147.020 3535.390 1150.020 3535.400 ;
        RECT 1237.020 3535.390 1240.020 3535.400 ;
        RECT 1327.020 3535.390 1330.020 3535.400 ;
        RECT 1417.020 3535.390 1420.020 3535.400 ;
        RECT 1507.020 3535.390 1510.020 3535.400 ;
        RECT 1597.020 3535.390 1600.020 3535.400 ;
        RECT 1687.020 3535.390 1690.020 3535.400 ;
        RECT 1777.020 3535.390 1780.020 3535.400 ;
        RECT 1867.020 3535.390 1870.020 3535.400 ;
        RECT 1957.020 3535.390 1960.020 3535.400 ;
        RECT 2047.020 3535.390 2050.020 3535.400 ;
        RECT 2137.020 3535.390 2140.020 3535.400 ;
        RECT 2227.020 3535.390 2230.020 3535.400 ;
        RECT 2317.020 3535.390 2320.020 3535.400 ;
        RECT 2407.020 3535.390 2410.020 3535.400 ;
        RECT 2497.020 3535.390 2500.020 3535.400 ;
        RECT 2587.020 3535.390 2590.020 3535.400 ;
        RECT 2677.020 3535.390 2680.020 3535.400 ;
        RECT 2767.020 3535.390 2770.020 3535.400 ;
        RECT 2857.020 3535.390 2860.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3495.380 -21.080 3495.390 ;
        RECT 2940.700 3495.380 2943.700 3495.390 ;
        RECT -24.080 3492.380 0.300 3495.380 ;
        RECT 2919.700 3492.380 2943.700 3495.380 ;
        RECT -24.080 3492.370 -21.080 3492.380 ;
        RECT 2940.700 3492.370 2943.700 3492.380 ;
        RECT -24.080 3405.380 -21.080 3405.390 ;
        RECT 2940.700 3405.380 2943.700 3405.390 ;
        RECT -24.080 3402.380 0.300 3405.380 ;
        RECT 2919.700 3402.380 2943.700 3405.380 ;
        RECT -24.080 3402.370 -21.080 3402.380 ;
        RECT 2940.700 3402.370 2943.700 3402.380 ;
        RECT -24.080 3315.380 -21.080 3315.390 ;
        RECT 2940.700 3315.380 2943.700 3315.390 ;
        RECT -24.080 3312.380 0.300 3315.380 ;
        RECT 2919.700 3312.380 2943.700 3315.380 ;
        RECT -24.080 3312.370 -21.080 3312.380 ;
        RECT 2940.700 3312.370 2943.700 3312.380 ;
        RECT -24.080 3225.380 -21.080 3225.390 ;
        RECT 2940.700 3225.380 2943.700 3225.390 ;
        RECT -24.080 3222.380 0.300 3225.380 ;
        RECT 2919.700 3222.380 2943.700 3225.380 ;
        RECT -24.080 3222.370 -21.080 3222.380 ;
        RECT 2940.700 3222.370 2943.700 3222.380 ;
        RECT -24.080 3135.380 -21.080 3135.390 ;
        RECT 2940.700 3135.380 2943.700 3135.390 ;
        RECT -24.080 3132.380 0.300 3135.380 ;
        RECT 2919.700 3132.380 2943.700 3135.380 ;
        RECT -24.080 3132.370 -21.080 3132.380 ;
        RECT 2940.700 3132.370 2943.700 3132.380 ;
        RECT -24.080 3045.380 -21.080 3045.390 ;
        RECT 2940.700 3045.380 2943.700 3045.390 ;
        RECT -24.080 3042.380 0.300 3045.380 ;
        RECT 2919.700 3042.380 2943.700 3045.380 ;
        RECT -24.080 3042.370 -21.080 3042.380 ;
        RECT 2940.700 3042.370 2943.700 3042.380 ;
        RECT -24.080 2955.380 -21.080 2955.390 ;
        RECT 2940.700 2955.380 2943.700 2955.390 ;
        RECT -24.080 2952.380 0.300 2955.380 ;
        RECT 2919.700 2952.380 2943.700 2955.380 ;
        RECT -24.080 2952.370 -21.080 2952.380 ;
        RECT 2940.700 2952.370 2943.700 2952.380 ;
        RECT -24.080 2865.380 -21.080 2865.390 ;
        RECT 2940.700 2865.380 2943.700 2865.390 ;
        RECT -24.080 2862.380 0.300 2865.380 ;
        RECT 2919.700 2862.380 2943.700 2865.380 ;
        RECT -24.080 2862.370 -21.080 2862.380 ;
        RECT 2940.700 2862.370 2943.700 2862.380 ;
        RECT -24.080 2775.380 -21.080 2775.390 ;
        RECT 2940.700 2775.380 2943.700 2775.390 ;
        RECT -24.080 2772.380 0.300 2775.380 ;
        RECT 2919.700 2772.380 2943.700 2775.380 ;
        RECT -24.080 2772.370 -21.080 2772.380 ;
        RECT 2940.700 2772.370 2943.700 2772.380 ;
        RECT -24.080 2685.380 -21.080 2685.390 ;
        RECT 2940.700 2685.380 2943.700 2685.390 ;
        RECT -24.080 2682.380 0.300 2685.380 ;
        RECT 2919.700 2682.380 2943.700 2685.380 ;
        RECT -24.080 2682.370 -21.080 2682.380 ;
        RECT 2940.700 2682.370 2943.700 2682.380 ;
        RECT -24.080 2595.380 -21.080 2595.390 ;
        RECT 2940.700 2595.380 2943.700 2595.390 ;
        RECT -24.080 2592.380 0.300 2595.380 ;
        RECT 2919.700 2592.380 2943.700 2595.380 ;
        RECT -24.080 2592.370 -21.080 2592.380 ;
        RECT 2940.700 2592.370 2943.700 2592.380 ;
        RECT -24.080 2505.380 -21.080 2505.390 ;
        RECT 2940.700 2505.380 2943.700 2505.390 ;
        RECT -24.080 2502.380 0.300 2505.380 ;
        RECT 2919.700 2502.380 2943.700 2505.380 ;
        RECT -24.080 2502.370 -21.080 2502.380 ;
        RECT 2940.700 2502.370 2943.700 2502.380 ;
        RECT -24.080 2415.380 -21.080 2415.390 ;
        RECT 2940.700 2415.380 2943.700 2415.390 ;
        RECT -24.080 2412.380 0.300 2415.380 ;
        RECT 2919.700 2412.380 2943.700 2415.380 ;
        RECT -24.080 2412.370 -21.080 2412.380 ;
        RECT 2940.700 2412.370 2943.700 2412.380 ;
        RECT -24.080 2325.380 -21.080 2325.390 ;
        RECT 2940.700 2325.380 2943.700 2325.390 ;
        RECT -24.080 2322.380 0.300 2325.380 ;
        RECT 2919.700 2322.380 2943.700 2325.380 ;
        RECT -24.080 2322.370 -21.080 2322.380 ;
        RECT 2940.700 2322.370 2943.700 2322.380 ;
        RECT -24.080 2235.380 -21.080 2235.390 ;
        RECT 2940.700 2235.380 2943.700 2235.390 ;
        RECT -24.080 2232.380 0.300 2235.380 ;
        RECT 2919.700 2232.380 2943.700 2235.380 ;
        RECT -24.080 2232.370 -21.080 2232.380 ;
        RECT 2940.700 2232.370 2943.700 2232.380 ;
        RECT -24.080 2145.380 -21.080 2145.390 ;
        RECT 2940.700 2145.380 2943.700 2145.390 ;
        RECT -24.080 2142.380 0.300 2145.380 ;
        RECT 2919.700 2142.380 2943.700 2145.380 ;
        RECT -24.080 2142.370 -21.080 2142.380 ;
        RECT 2940.700 2142.370 2943.700 2142.380 ;
        RECT -24.080 2055.380 -21.080 2055.390 ;
        RECT 2940.700 2055.380 2943.700 2055.390 ;
        RECT -24.080 2052.380 0.300 2055.380 ;
        RECT 2919.700 2052.380 2943.700 2055.380 ;
        RECT -24.080 2052.370 -21.080 2052.380 ;
        RECT 2940.700 2052.370 2943.700 2052.380 ;
        RECT -24.080 1965.380 -21.080 1965.390 ;
        RECT 2940.700 1965.380 2943.700 1965.390 ;
        RECT -24.080 1962.380 0.300 1965.380 ;
        RECT 2919.700 1962.380 2943.700 1965.380 ;
        RECT -24.080 1962.370 -21.080 1962.380 ;
        RECT 2940.700 1962.370 2943.700 1962.380 ;
        RECT -24.080 1875.380 -21.080 1875.390 ;
        RECT 2940.700 1875.380 2943.700 1875.390 ;
        RECT -24.080 1872.380 0.300 1875.380 ;
        RECT 2919.700 1872.380 2943.700 1875.380 ;
        RECT -24.080 1872.370 -21.080 1872.380 ;
        RECT 2940.700 1872.370 2943.700 1872.380 ;
        RECT -24.080 1785.380 -21.080 1785.390 ;
        RECT 2940.700 1785.380 2943.700 1785.390 ;
        RECT -24.080 1782.380 0.300 1785.380 ;
        RECT 2919.700 1782.380 2943.700 1785.380 ;
        RECT -24.080 1782.370 -21.080 1782.380 ;
        RECT 2940.700 1782.370 2943.700 1782.380 ;
        RECT -24.080 1695.380 -21.080 1695.390 ;
        RECT 2940.700 1695.380 2943.700 1695.390 ;
        RECT -24.080 1692.380 0.300 1695.380 ;
        RECT 2919.700 1692.380 2943.700 1695.380 ;
        RECT -24.080 1692.370 -21.080 1692.380 ;
        RECT 2940.700 1692.370 2943.700 1692.380 ;
        RECT -24.080 1605.380 -21.080 1605.390 ;
        RECT 2940.700 1605.380 2943.700 1605.390 ;
        RECT -24.080 1602.380 0.300 1605.380 ;
        RECT 2919.700 1602.380 2943.700 1605.380 ;
        RECT -24.080 1602.370 -21.080 1602.380 ;
        RECT 2940.700 1602.370 2943.700 1602.380 ;
        RECT -24.080 1515.380 -21.080 1515.390 ;
        RECT 2940.700 1515.380 2943.700 1515.390 ;
        RECT -24.080 1512.380 0.300 1515.380 ;
        RECT 2919.700 1512.380 2943.700 1515.380 ;
        RECT -24.080 1512.370 -21.080 1512.380 ;
        RECT 2940.700 1512.370 2943.700 1512.380 ;
        RECT -24.080 1425.380 -21.080 1425.390 ;
        RECT 2940.700 1425.380 2943.700 1425.390 ;
        RECT -24.080 1422.380 0.300 1425.380 ;
        RECT 2919.700 1422.380 2943.700 1425.380 ;
        RECT -24.080 1422.370 -21.080 1422.380 ;
        RECT 2940.700 1422.370 2943.700 1422.380 ;
        RECT -24.080 1335.380 -21.080 1335.390 ;
        RECT 2940.700 1335.380 2943.700 1335.390 ;
        RECT -24.080 1332.380 0.300 1335.380 ;
        RECT 2919.700 1332.380 2943.700 1335.380 ;
        RECT -24.080 1332.370 -21.080 1332.380 ;
        RECT 2940.700 1332.370 2943.700 1332.380 ;
        RECT -24.080 1245.380 -21.080 1245.390 ;
        RECT 2940.700 1245.380 2943.700 1245.390 ;
        RECT -24.080 1242.380 0.300 1245.380 ;
        RECT 2919.700 1242.380 2943.700 1245.380 ;
        RECT -24.080 1242.370 -21.080 1242.380 ;
        RECT 2940.700 1242.370 2943.700 1242.380 ;
        RECT -24.080 1155.380 -21.080 1155.390 ;
        RECT 2940.700 1155.380 2943.700 1155.390 ;
        RECT -24.080 1152.380 0.300 1155.380 ;
        RECT 2919.700 1152.380 2943.700 1155.380 ;
        RECT -24.080 1152.370 -21.080 1152.380 ;
        RECT 2940.700 1152.370 2943.700 1152.380 ;
        RECT -24.080 1065.380 -21.080 1065.390 ;
        RECT 2940.700 1065.380 2943.700 1065.390 ;
        RECT -24.080 1062.380 0.300 1065.380 ;
        RECT 2919.700 1062.380 2943.700 1065.380 ;
        RECT -24.080 1062.370 -21.080 1062.380 ;
        RECT 2940.700 1062.370 2943.700 1062.380 ;
        RECT -24.080 975.380 -21.080 975.390 ;
        RECT 2940.700 975.380 2943.700 975.390 ;
        RECT -24.080 972.380 0.300 975.380 ;
        RECT 2919.700 972.380 2943.700 975.380 ;
        RECT -24.080 972.370 -21.080 972.380 ;
        RECT 2940.700 972.370 2943.700 972.380 ;
        RECT -24.080 885.380 -21.080 885.390 ;
        RECT 2940.700 885.380 2943.700 885.390 ;
        RECT -24.080 882.380 0.300 885.380 ;
        RECT 2919.700 882.380 2943.700 885.380 ;
        RECT -24.080 882.370 -21.080 882.380 ;
        RECT 2940.700 882.370 2943.700 882.380 ;
        RECT -24.080 795.380 -21.080 795.390 ;
        RECT 2940.700 795.380 2943.700 795.390 ;
        RECT -24.080 792.380 0.300 795.380 ;
        RECT 2919.700 792.380 2943.700 795.380 ;
        RECT -24.080 792.370 -21.080 792.380 ;
        RECT 2940.700 792.370 2943.700 792.380 ;
        RECT -24.080 705.380 -21.080 705.390 ;
        RECT 2940.700 705.380 2943.700 705.390 ;
        RECT -24.080 702.380 0.300 705.380 ;
        RECT 2919.700 702.380 2943.700 705.380 ;
        RECT -24.080 702.370 -21.080 702.380 ;
        RECT 2940.700 702.370 2943.700 702.380 ;
        RECT -24.080 615.380 -21.080 615.390 ;
        RECT 2940.700 615.380 2943.700 615.390 ;
        RECT -24.080 612.380 0.300 615.380 ;
        RECT 2919.700 612.380 2943.700 615.380 ;
        RECT -24.080 612.370 -21.080 612.380 ;
        RECT 2940.700 612.370 2943.700 612.380 ;
        RECT -24.080 525.380 -21.080 525.390 ;
        RECT 2940.700 525.380 2943.700 525.390 ;
        RECT -24.080 522.380 0.300 525.380 ;
        RECT 2919.700 522.380 2943.700 525.380 ;
        RECT -24.080 522.370 -21.080 522.380 ;
        RECT 2940.700 522.370 2943.700 522.380 ;
        RECT -24.080 435.380 -21.080 435.390 ;
        RECT 2940.700 435.380 2943.700 435.390 ;
        RECT -24.080 432.380 0.300 435.380 ;
        RECT 2919.700 432.380 2943.700 435.380 ;
        RECT -24.080 432.370 -21.080 432.380 ;
        RECT 2940.700 432.370 2943.700 432.380 ;
        RECT -24.080 345.380 -21.080 345.390 ;
        RECT 2940.700 345.380 2943.700 345.390 ;
        RECT -24.080 342.380 0.300 345.380 ;
        RECT 2919.700 342.380 2943.700 345.380 ;
        RECT -24.080 342.370 -21.080 342.380 ;
        RECT 2940.700 342.370 2943.700 342.380 ;
        RECT -24.080 255.380 -21.080 255.390 ;
        RECT 2940.700 255.380 2943.700 255.390 ;
        RECT -24.080 252.380 0.300 255.380 ;
        RECT 2919.700 252.380 2943.700 255.380 ;
        RECT -24.080 252.370 -21.080 252.380 ;
        RECT 2940.700 252.370 2943.700 252.380 ;
        RECT -24.080 165.380 -21.080 165.390 ;
        RECT 2940.700 165.380 2943.700 165.390 ;
        RECT -24.080 162.380 0.300 165.380 ;
        RECT 2919.700 162.380 2943.700 165.380 ;
        RECT -24.080 162.370 -21.080 162.380 ;
        RECT 2940.700 162.370 2943.700 162.380 ;
        RECT -24.080 75.380 -21.080 75.390 ;
        RECT 2940.700 75.380 2943.700 75.390 ;
        RECT -24.080 72.380 0.300 75.380 ;
        RECT 2919.700 72.380 2943.700 75.380 ;
        RECT -24.080 72.370 -21.080 72.380 ;
        RECT 2940.700 72.370 2943.700 72.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 67.020 -15.720 70.020 -15.710 ;
        RECT 157.020 -15.720 160.020 -15.710 ;
        RECT 247.020 -15.720 250.020 -15.710 ;
        RECT 337.020 -15.720 340.020 -15.710 ;
        RECT 427.020 -15.720 430.020 -15.710 ;
        RECT 517.020 -15.720 520.020 -15.710 ;
        RECT 607.020 -15.720 610.020 -15.710 ;
        RECT 697.020 -15.720 700.020 -15.710 ;
        RECT 787.020 -15.720 790.020 -15.710 ;
        RECT 877.020 -15.720 880.020 -15.710 ;
        RECT 967.020 -15.720 970.020 -15.710 ;
        RECT 1057.020 -15.720 1060.020 -15.710 ;
        RECT 1147.020 -15.720 1150.020 -15.710 ;
        RECT 1237.020 -15.720 1240.020 -15.710 ;
        RECT 1327.020 -15.720 1330.020 -15.710 ;
        RECT 1417.020 -15.720 1420.020 -15.710 ;
        RECT 1507.020 -15.720 1510.020 -15.710 ;
        RECT 1597.020 -15.720 1600.020 -15.710 ;
        RECT 1687.020 -15.720 1690.020 -15.710 ;
        RECT 1777.020 -15.720 1780.020 -15.710 ;
        RECT 1867.020 -15.720 1870.020 -15.710 ;
        RECT 1957.020 -15.720 1960.020 -15.710 ;
        RECT 2047.020 -15.720 2050.020 -15.710 ;
        RECT 2137.020 -15.720 2140.020 -15.710 ;
        RECT 2227.020 -15.720 2230.020 -15.710 ;
        RECT 2317.020 -15.720 2320.020 -15.710 ;
        RECT 2407.020 -15.720 2410.020 -15.710 ;
        RECT 2497.020 -15.720 2500.020 -15.710 ;
        RECT 2587.020 -15.720 2590.020 -15.710 ;
        RECT 2677.020 -15.720 2680.020 -15.710 ;
        RECT 2767.020 -15.720 2770.020 -15.710 ;
        RECT 2857.020 -15.720 2860.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 67.020 -18.730 70.020 -18.720 ;
        RECT 157.020 -18.730 160.020 -18.720 ;
        RECT 247.020 -18.730 250.020 -18.720 ;
        RECT 337.020 -18.730 340.020 -18.720 ;
        RECT 427.020 -18.730 430.020 -18.720 ;
        RECT 517.020 -18.730 520.020 -18.720 ;
        RECT 607.020 -18.730 610.020 -18.720 ;
        RECT 697.020 -18.730 700.020 -18.720 ;
        RECT 787.020 -18.730 790.020 -18.720 ;
        RECT 877.020 -18.730 880.020 -18.720 ;
        RECT 967.020 -18.730 970.020 -18.720 ;
        RECT 1057.020 -18.730 1060.020 -18.720 ;
        RECT 1147.020 -18.730 1150.020 -18.720 ;
        RECT 1237.020 -18.730 1240.020 -18.720 ;
        RECT 1327.020 -18.730 1330.020 -18.720 ;
        RECT 1417.020 -18.730 1420.020 -18.720 ;
        RECT 1507.020 -18.730 1510.020 -18.720 ;
        RECT 1597.020 -18.730 1600.020 -18.720 ;
        RECT 1687.020 -18.730 1690.020 -18.720 ;
        RECT 1777.020 -18.730 1780.020 -18.720 ;
        RECT 1867.020 -18.730 1870.020 -18.720 ;
        RECT 1957.020 -18.730 1960.020 -18.720 ;
        RECT 2047.020 -18.730 2050.020 -18.720 ;
        RECT 2137.020 -18.730 2140.020 -18.720 ;
        RECT 2227.020 -18.730 2230.020 -18.720 ;
        RECT 2317.020 -18.730 2320.020 -18.720 ;
        RECT 2407.020 -18.730 2410.020 -18.720 ;
        RECT 2497.020 -18.730 2500.020 -18.720 ;
        RECT 2587.020 -18.730 2590.020 -18.720 ;
        RECT 2677.020 -18.730 2680.020 -18.720 ;
        RECT 2767.020 -18.730 2770.020 -18.720 ;
        RECT 2857.020 -18.730 2860.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 3519.700 43.020 3547.800 ;
        RECT 130.020 3519.700 133.020 3547.800 ;
        RECT 220.020 3519.700 223.020 3547.800 ;
        RECT 310.020 3519.700 313.020 3547.800 ;
        RECT 400.020 3519.700 403.020 3547.800 ;
        RECT 490.020 3519.700 493.020 3547.800 ;
        RECT 580.020 3519.700 583.020 3547.800 ;
        RECT 670.020 3519.700 673.020 3547.800 ;
        RECT 760.020 3519.700 763.020 3547.800 ;
        RECT 850.020 3519.700 853.020 3547.800 ;
        RECT 940.020 3519.700 943.020 3547.800 ;
        RECT 1030.020 3519.700 1033.020 3547.800 ;
        RECT 1120.020 3519.700 1123.020 3547.800 ;
        RECT 1210.020 3519.700 1213.020 3547.800 ;
        RECT 1300.020 3519.700 1303.020 3547.800 ;
        RECT 1390.020 3519.700 1393.020 3547.800 ;
        RECT 1480.020 3519.700 1483.020 3547.800 ;
        RECT 1570.020 3519.700 1573.020 3547.800 ;
        RECT 1660.020 3519.700 1663.020 3547.800 ;
        RECT 1750.020 3519.700 1753.020 3547.800 ;
        RECT 1840.020 3519.700 1843.020 3547.800 ;
        RECT 1930.020 3519.700 1933.020 3547.800 ;
        RECT 2020.020 3519.700 2023.020 3547.800 ;
        RECT 2110.020 3519.700 2113.020 3547.800 ;
        RECT 2200.020 3519.700 2203.020 3547.800 ;
        RECT 2290.020 3519.700 2293.020 3547.800 ;
        RECT 2380.020 3519.700 2383.020 3547.800 ;
        RECT 2470.020 3519.700 2473.020 3547.800 ;
        RECT 2560.020 3519.700 2563.020 3547.800 ;
        RECT 2650.020 3519.700 2653.020 3547.800 ;
        RECT 2740.020 3519.700 2743.020 3547.800 ;
        RECT 2830.020 3519.700 2833.020 3547.800 ;
        RECT 40.020 -28.120 43.020 0.300 ;
        RECT 130.020 -28.120 133.020 0.300 ;
        RECT 220.020 -28.120 223.020 0.300 ;
        RECT 310.020 -28.120 313.020 0.300 ;
        RECT 400.020 -28.120 403.020 0.300 ;
        RECT 490.020 -28.120 493.020 0.300 ;
        RECT 580.020 -28.120 583.020 0.300 ;
        RECT 670.020 -28.120 673.020 0.300 ;
        RECT 760.020 -28.120 763.020 0.300 ;
        RECT 850.020 -28.120 853.020 0.300 ;
        RECT 940.020 -28.120 943.020 0.300 ;
        RECT 1030.020 -28.120 1033.020 0.300 ;
        RECT 1120.020 -28.120 1123.020 0.300 ;
        RECT 1210.020 -28.120 1213.020 0.300 ;
        RECT 1300.020 -28.120 1303.020 0.300 ;
        RECT 1390.020 -28.120 1393.020 0.300 ;
        RECT 1480.020 -28.120 1483.020 0.300 ;
        RECT 1570.020 -28.120 1573.020 0.300 ;
        RECT 1660.020 -28.120 1663.020 0.300 ;
        RECT 1750.020 -28.120 1753.020 0.300 ;
        RECT 1840.020 -28.120 1843.020 0.300 ;
        RECT 1930.020 -28.120 1933.020 0.300 ;
        RECT 2020.020 -28.120 2023.020 0.300 ;
        RECT 2110.020 -28.120 2113.020 0.300 ;
        RECT 2200.020 -28.120 2203.020 0.300 ;
        RECT 2290.020 -28.120 2293.020 0.300 ;
        RECT 2380.020 -28.120 2383.020 0.300 ;
        RECT 2470.020 -28.120 2473.020 0.300 ;
        RECT 2560.020 -28.120 2563.020 0.300 ;
        RECT 2650.020 -28.120 2653.020 0.300 ;
        RECT 2740.020 -28.120 2743.020 0.300 ;
        RECT 2830.020 -28.120 2833.020 0.300 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 130.930 3541.810 132.110 3542.990 ;
        RECT 130.930 3540.210 132.110 3541.390 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 310.930 3541.810 312.110 3542.990 ;
        RECT 310.930 3540.210 312.110 3541.390 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 490.930 3541.810 492.110 3542.990 ;
        RECT 490.930 3540.210 492.110 3541.390 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 670.930 3541.810 672.110 3542.990 ;
        RECT 670.930 3540.210 672.110 3541.390 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 850.930 3541.810 852.110 3542.990 ;
        RECT 850.930 3540.210 852.110 3541.390 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 1030.930 3541.810 1032.110 3542.990 ;
        RECT 1030.930 3540.210 1032.110 3541.390 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1210.930 3541.810 1212.110 3542.990 ;
        RECT 1210.930 3540.210 1212.110 3541.390 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1390.930 3541.810 1392.110 3542.990 ;
        RECT 1390.930 3540.210 1392.110 3541.390 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1570.930 3541.810 1572.110 3542.990 ;
        RECT 1570.930 3540.210 1572.110 3541.390 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1750.930 3541.810 1752.110 3542.990 ;
        RECT 1750.930 3540.210 1752.110 3541.390 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1930.930 3541.810 1932.110 3542.990 ;
        RECT 1930.930 3540.210 1932.110 3541.390 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2110.930 3541.810 2112.110 3542.990 ;
        RECT 2110.930 3540.210 2112.110 3541.390 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2290.930 3541.810 2292.110 3542.990 ;
        RECT 2290.930 3540.210 2292.110 3541.390 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2470.930 3541.810 2472.110 3542.990 ;
        RECT 2470.930 3540.210 2472.110 3541.390 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2650.930 3541.810 2652.110 3542.990 ;
        RECT 2650.930 3540.210 2652.110 3541.390 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2830.930 3541.810 2832.110 3542.990 ;
        RECT 2830.930 3540.210 2832.110 3541.390 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3377.090 -26.690 3378.270 ;
        RECT -27.870 3375.490 -26.690 3376.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3197.090 -26.690 3198.270 ;
        RECT -27.870 3195.490 -26.690 3196.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 3017.090 -26.690 3018.270 ;
        RECT -27.870 3015.490 -26.690 3016.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2837.090 -26.690 2838.270 ;
        RECT -27.870 2835.490 -26.690 2836.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2657.090 -26.690 2658.270 ;
        RECT -27.870 2655.490 -26.690 2656.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2477.090 -26.690 2478.270 ;
        RECT -27.870 2475.490 -26.690 2476.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2297.090 -26.690 2298.270 ;
        RECT -27.870 2295.490 -26.690 2296.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2117.090 -26.690 2118.270 ;
        RECT -27.870 2115.490 -26.690 2116.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1937.090 -26.690 1938.270 ;
        RECT -27.870 1935.490 -26.690 1936.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1757.090 -26.690 1758.270 ;
        RECT -27.870 1755.490 -26.690 1756.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1577.090 -26.690 1578.270 ;
        RECT -27.870 1575.490 -26.690 1576.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1397.090 -26.690 1398.270 ;
        RECT -27.870 1395.490 -26.690 1396.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1217.090 -26.690 1218.270 ;
        RECT -27.870 1215.490 -26.690 1216.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 1037.090 -26.690 1038.270 ;
        RECT -27.870 1035.490 -26.690 1036.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 857.090 -26.690 858.270 ;
        RECT -27.870 855.490 -26.690 856.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 677.090 -26.690 678.270 ;
        RECT -27.870 675.490 -26.690 676.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 497.090 -26.690 498.270 ;
        RECT -27.870 495.490 -26.690 496.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 317.090 -26.690 318.270 ;
        RECT -27.870 315.490 -26.690 316.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 137.090 -26.690 138.270 ;
        RECT -27.870 135.490 -26.690 136.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3377.090 2947.490 3378.270 ;
        RECT 2946.310 3375.490 2947.490 3376.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3197.090 2947.490 3198.270 ;
        RECT 2946.310 3195.490 2947.490 3196.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 3017.090 2947.490 3018.270 ;
        RECT 2946.310 3015.490 2947.490 3016.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2837.090 2947.490 2838.270 ;
        RECT 2946.310 2835.490 2947.490 2836.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2657.090 2947.490 2658.270 ;
        RECT 2946.310 2655.490 2947.490 2656.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2477.090 2947.490 2478.270 ;
        RECT 2946.310 2475.490 2947.490 2476.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2297.090 2947.490 2298.270 ;
        RECT 2946.310 2295.490 2947.490 2296.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2117.090 2947.490 2118.270 ;
        RECT 2946.310 2115.490 2947.490 2116.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1937.090 2947.490 1938.270 ;
        RECT 2946.310 1935.490 2947.490 1936.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1757.090 2947.490 1758.270 ;
        RECT 2946.310 1755.490 2947.490 1756.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1577.090 2947.490 1578.270 ;
        RECT 2946.310 1575.490 2947.490 1576.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1397.090 2947.490 1398.270 ;
        RECT 2946.310 1395.490 2947.490 1396.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1217.090 2947.490 1218.270 ;
        RECT 2946.310 1215.490 2947.490 1216.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 1037.090 2947.490 1038.270 ;
        RECT 2946.310 1035.490 2947.490 1036.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 857.090 2947.490 858.270 ;
        RECT 2946.310 855.490 2947.490 856.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 677.090 2947.490 678.270 ;
        RECT 2946.310 675.490 2947.490 676.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 497.090 2947.490 498.270 ;
        RECT 2946.310 495.490 2947.490 496.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 317.090 2947.490 318.270 ;
        RECT 2946.310 315.490 2947.490 316.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 137.090 2947.490 138.270 ;
        RECT 2946.310 135.490 2947.490 136.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 130.930 -21.710 132.110 -20.530 ;
        RECT 130.930 -23.310 132.110 -22.130 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 310.930 -21.710 312.110 -20.530 ;
        RECT 310.930 -23.310 312.110 -22.130 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 490.930 -21.710 492.110 -20.530 ;
        RECT 490.930 -23.310 492.110 -22.130 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 670.930 -21.710 672.110 -20.530 ;
        RECT 670.930 -23.310 672.110 -22.130 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 850.930 -21.710 852.110 -20.530 ;
        RECT 850.930 -23.310 852.110 -22.130 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1030.930 -21.710 1032.110 -20.530 ;
        RECT 1030.930 -23.310 1032.110 -22.130 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1210.930 -21.710 1212.110 -20.530 ;
        RECT 1210.930 -23.310 1212.110 -22.130 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1390.930 -21.710 1392.110 -20.530 ;
        RECT 1390.930 -23.310 1392.110 -22.130 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1570.930 -21.710 1572.110 -20.530 ;
        RECT 1570.930 -23.310 1572.110 -22.130 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1750.930 -21.710 1752.110 -20.530 ;
        RECT 1750.930 -23.310 1752.110 -22.130 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 1930.930 -21.710 1932.110 -20.530 ;
        RECT 1930.930 -23.310 1932.110 -22.130 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2110.930 -21.710 2112.110 -20.530 ;
        RECT 2110.930 -23.310 2112.110 -22.130 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2290.930 -21.710 2292.110 -20.530 ;
        RECT 2290.930 -23.310 2292.110 -22.130 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2470.930 -21.710 2472.110 -20.530 ;
        RECT 2470.930 -23.310 2472.110 -22.130 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2650.930 -21.710 2652.110 -20.530 ;
        RECT 2650.930 -23.310 2652.110 -22.130 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2830.930 -21.710 2832.110 -20.530 ;
        RECT 2830.930 -23.310 2832.110 -22.130 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 130.020 3543.100 133.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 310.020 3543.100 313.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 490.020 3543.100 493.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 670.020 3543.100 673.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 850.020 3543.100 853.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1030.020 3543.100 1033.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1210.020 3543.100 1213.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1390.020 3543.100 1393.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1570.020 3543.100 1573.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1750.020 3543.100 1753.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 1930.020 3543.100 1933.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2110.020 3543.100 2113.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2290.020 3543.100 2293.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2470.020 3543.100 2473.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2650.020 3543.100 2653.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2830.020 3543.100 2833.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 130.020 3540.090 133.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 310.020 3540.090 313.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 490.020 3540.090 493.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 670.020 3540.090 673.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 850.020 3540.090 853.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1030.020 3540.090 1033.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1210.020 3540.090 1213.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1390.020 3540.090 1393.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1570.020 3540.090 1573.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1750.020 3540.090 1753.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 1930.020 3540.090 1933.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2110.020 3540.090 2113.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2290.020 3540.090 2293.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2470.020 3540.090 2473.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2650.020 3540.090 2653.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2830.020 3540.090 2833.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 0.300 3468.380 ;
        RECT 2919.700 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3378.380 -25.780 3378.390 ;
        RECT 2945.400 3378.380 2948.400 3378.390 ;
        RECT -33.480 3375.380 0.300 3378.380 ;
        RECT 2919.700 3375.380 2953.100 3378.380 ;
        RECT -28.780 3375.370 -25.780 3375.380 ;
        RECT 2945.400 3375.370 2948.400 3375.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 0.300 3288.380 ;
        RECT 2919.700 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3198.380 -25.780 3198.390 ;
        RECT 2945.400 3198.380 2948.400 3198.390 ;
        RECT -33.480 3195.380 0.300 3198.380 ;
        RECT 2919.700 3195.380 2953.100 3198.380 ;
        RECT -28.780 3195.370 -25.780 3195.380 ;
        RECT 2945.400 3195.370 2948.400 3195.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 0.300 3108.380 ;
        RECT 2919.700 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 3018.380 -25.780 3018.390 ;
        RECT 2945.400 3018.380 2948.400 3018.390 ;
        RECT -33.480 3015.380 0.300 3018.380 ;
        RECT 2919.700 3015.380 2953.100 3018.380 ;
        RECT -28.780 3015.370 -25.780 3015.380 ;
        RECT 2945.400 3015.370 2948.400 3015.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 0.300 2928.380 ;
        RECT 2919.700 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2838.380 -25.780 2838.390 ;
        RECT 2945.400 2838.380 2948.400 2838.390 ;
        RECT -33.480 2835.380 0.300 2838.380 ;
        RECT 2919.700 2835.380 2953.100 2838.380 ;
        RECT -28.780 2835.370 -25.780 2835.380 ;
        RECT 2945.400 2835.370 2948.400 2835.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 0.300 2748.380 ;
        RECT 2919.700 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2658.380 -25.780 2658.390 ;
        RECT 2945.400 2658.380 2948.400 2658.390 ;
        RECT -33.480 2655.380 0.300 2658.380 ;
        RECT 2919.700 2655.380 2953.100 2658.380 ;
        RECT -28.780 2655.370 -25.780 2655.380 ;
        RECT 2945.400 2655.370 2948.400 2655.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 0.300 2568.380 ;
        RECT 2919.700 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2478.380 -25.780 2478.390 ;
        RECT 2945.400 2478.380 2948.400 2478.390 ;
        RECT -33.480 2475.380 0.300 2478.380 ;
        RECT 2919.700 2475.380 2953.100 2478.380 ;
        RECT -28.780 2475.370 -25.780 2475.380 ;
        RECT 2945.400 2475.370 2948.400 2475.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 0.300 2388.380 ;
        RECT 2919.700 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2298.380 -25.780 2298.390 ;
        RECT 2945.400 2298.380 2948.400 2298.390 ;
        RECT -33.480 2295.380 0.300 2298.380 ;
        RECT 2919.700 2295.380 2953.100 2298.380 ;
        RECT -28.780 2295.370 -25.780 2295.380 ;
        RECT 2945.400 2295.370 2948.400 2295.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 0.300 2208.380 ;
        RECT 2919.700 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2118.380 -25.780 2118.390 ;
        RECT 2945.400 2118.380 2948.400 2118.390 ;
        RECT -33.480 2115.380 0.300 2118.380 ;
        RECT 2919.700 2115.380 2953.100 2118.380 ;
        RECT -28.780 2115.370 -25.780 2115.380 ;
        RECT 2945.400 2115.370 2948.400 2115.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 0.300 2028.380 ;
        RECT 2919.700 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1938.380 -25.780 1938.390 ;
        RECT 2945.400 1938.380 2948.400 1938.390 ;
        RECT -33.480 1935.380 0.300 1938.380 ;
        RECT 2919.700 1935.380 2953.100 1938.380 ;
        RECT -28.780 1935.370 -25.780 1935.380 ;
        RECT 2945.400 1935.370 2948.400 1935.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 0.300 1848.380 ;
        RECT 2919.700 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1758.380 -25.780 1758.390 ;
        RECT 2945.400 1758.380 2948.400 1758.390 ;
        RECT -33.480 1755.380 0.300 1758.380 ;
        RECT 2919.700 1755.380 2953.100 1758.380 ;
        RECT -28.780 1755.370 -25.780 1755.380 ;
        RECT 2945.400 1755.370 2948.400 1755.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 0.300 1668.380 ;
        RECT 2919.700 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1578.380 -25.780 1578.390 ;
        RECT 2945.400 1578.380 2948.400 1578.390 ;
        RECT -33.480 1575.380 0.300 1578.380 ;
        RECT 2919.700 1575.380 2953.100 1578.380 ;
        RECT -28.780 1575.370 -25.780 1575.380 ;
        RECT 2945.400 1575.370 2948.400 1575.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 0.300 1488.380 ;
        RECT 2919.700 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1398.380 -25.780 1398.390 ;
        RECT 2945.400 1398.380 2948.400 1398.390 ;
        RECT -33.480 1395.380 0.300 1398.380 ;
        RECT 2919.700 1395.380 2953.100 1398.380 ;
        RECT -28.780 1395.370 -25.780 1395.380 ;
        RECT 2945.400 1395.370 2948.400 1395.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 0.300 1308.380 ;
        RECT 2919.700 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1218.380 -25.780 1218.390 ;
        RECT 2945.400 1218.380 2948.400 1218.390 ;
        RECT -33.480 1215.380 0.300 1218.380 ;
        RECT 2919.700 1215.380 2953.100 1218.380 ;
        RECT -28.780 1215.370 -25.780 1215.380 ;
        RECT 2945.400 1215.370 2948.400 1215.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 0.300 1128.380 ;
        RECT 2919.700 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 1038.380 -25.780 1038.390 ;
        RECT 2945.400 1038.380 2948.400 1038.390 ;
        RECT -33.480 1035.380 0.300 1038.380 ;
        RECT 2919.700 1035.380 2953.100 1038.380 ;
        RECT -28.780 1035.370 -25.780 1035.380 ;
        RECT 2945.400 1035.370 2948.400 1035.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 0.300 948.380 ;
        RECT 2919.700 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 858.380 -25.780 858.390 ;
        RECT 2945.400 858.380 2948.400 858.390 ;
        RECT -33.480 855.380 0.300 858.380 ;
        RECT 2919.700 855.380 2953.100 858.380 ;
        RECT -28.780 855.370 -25.780 855.380 ;
        RECT 2945.400 855.370 2948.400 855.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 0.300 768.380 ;
        RECT 2919.700 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 678.380 -25.780 678.390 ;
        RECT 2945.400 678.380 2948.400 678.390 ;
        RECT -33.480 675.380 0.300 678.380 ;
        RECT 2919.700 675.380 2953.100 678.380 ;
        RECT -28.780 675.370 -25.780 675.380 ;
        RECT 2945.400 675.370 2948.400 675.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 0.300 588.380 ;
        RECT 2919.700 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 498.380 -25.780 498.390 ;
        RECT 2945.400 498.380 2948.400 498.390 ;
        RECT -33.480 495.380 0.300 498.380 ;
        RECT 2919.700 495.380 2953.100 498.380 ;
        RECT -28.780 495.370 -25.780 495.380 ;
        RECT 2945.400 495.370 2948.400 495.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 0.300 408.380 ;
        RECT 2919.700 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 318.380 -25.780 318.390 ;
        RECT 2945.400 318.380 2948.400 318.390 ;
        RECT -33.480 315.380 0.300 318.380 ;
        RECT 2919.700 315.380 2953.100 318.380 ;
        RECT -28.780 315.370 -25.780 315.380 ;
        RECT 2945.400 315.370 2948.400 315.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 0.300 228.380 ;
        RECT 2919.700 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 138.380 -25.780 138.390 ;
        RECT 2945.400 138.380 2948.400 138.390 ;
        RECT -33.480 135.380 0.300 138.380 ;
        RECT 2919.700 135.380 2953.100 138.380 ;
        RECT -28.780 135.370 -25.780 135.380 ;
        RECT 2945.400 135.370 2948.400 135.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 0.300 48.380 ;
        RECT 2919.700 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 130.020 -20.420 133.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 310.020 -20.420 313.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 490.020 -20.420 493.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 670.020 -20.420 673.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 850.020 -20.420 853.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1030.020 -20.420 1033.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1210.020 -20.420 1213.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1390.020 -20.420 1393.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1570.020 -20.420 1573.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1750.020 -20.420 1753.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 1930.020 -20.420 1933.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2110.020 -20.420 2113.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2290.020 -20.420 2293.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2470.020 -20.420 2473.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2650.020 -20.420 2653.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2830.020 -20.420 2833.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 130.020 -23.430 133.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 310.020 -23.430 313.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 490.020 -23.430 493.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 670.020 -23.430 673.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 850.020 -23.430 853.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1030.020 -23.430 1033.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1210.020 -23.430 1213.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1390.020 -23.430 1393.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1570.020 -23.430 1573.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1750.020 -23.430 1753.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 1930.020 -23.430 1933.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2110.020 -23.430 2113.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2290.020 -23.430 2293.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2470.020 -23.430 2473.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2650.020 -23.430 2653.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2830.020 -23.430 2833.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 85.020 3519.700 88.020 3547.800 ;
        RECT 175.020 3519.700 178.020 3547.800 ;
        RECT 265.020 3519.700 268.020 3547.800 ;
        RECT 355.020 3519.700 358.020 3547.800 ;
        RECT 445.020 3519.700 448.020 3547.800 ;
        RECT 535.020 3519.700 538.020 3547.800 ;
        RECT 625.020 3519.700 628.020 3547.800 ;
        RECT 715.020 3519.700 718.020 3547.800 ;
        RECT 805.020 3519.700 808.020 3547.800 ;
        RECT 895.020 3519.700 898.020 3547.800 ;
        RECT 985.020 3519.700 988.020 3547.800 ;
        RECT 1075.020 3519.700 1078.020 3547.800 ;
        RECT 1165.020 3519.700 1168.020 3547.800 ;
        RECT 1255.020 3519.700 1258.020 3547.800 ;
        RECT 1345.020 3519.700 1348.020 3547.800 ;
        RECT 1435.020 3519.700 1438.020 3547.800 ;
        RECT 1525.020 3519.700 1528.020 3547.800 ;
        RECT 1615.020 3519.700 1618.020 3547.800 ;
        RECT 1705.020 3519.700 1708.020 3547.800 ;
        RECT 1795.020 3519.700 1798.020 3547.800 ;
        RECT 1885.020 3519.700 1888.020 3547.800 ;
        RECT 1975.020 3519.700 1978.020 3547.800 ;
        RECT 2065.020 3519.700 2068.020 3547.800 ;
        RECT 2155.020 3519.700 2158.020 3547.800 ;
        RECT 2245.020 3519.700 2248.020 3547.800 ;
        RECT 2335.020 3519.700 2338.020 3547.800 ;
        RECT 2425.020 3519.700 2428.020 3547.800 ;
        RECT 2515.020 3519.700 2518.020 3547.800 ;
        RECT 2605.020 3519.700 2608.020 3547.800 ;
        RECT 2695.020 3519.700 2698.020 3547.800 ;
        RECT 2785.020 3519.700 2788.020 3547.800 ;
        RECT 2875.020 3519.700 2878.020 3547.800 ;
        RECT 85.020 -28.120 88.020 0.300 ;
        RECT 175.020 -28.120 178.020 0.300 ;
        RECT 265.020 -28.120 268.020 0.300 ;
        RECT 355.020 -28.120 358.020 0.300 ;
        RECT 445.020 -28.120 448.020 0.300 ;
        RECT 535.020 -28.120 538.020 0.300 ;
        RECT 625.020 -28.120 628.020 0.300 ;
        RECT 715.020 -28.120 718.020 0.300 ;
        RECT 805.020 -28.120 808.020 0.300 ;
        RECT 895.020 -28.120 898.020 0.300 ;
        RECT 985.020 -28.120 988.020 0.300 ;
        RECT 1075.020 -28.120 1078.020 0.300 ;
        RECT 1165.020 -28.120 1168.020 0.300 ;
        RECT 1255.020 -28.120 1258.020 0.300 ;
        RECT 1345.020 -28.120 1348.020 0.300 ;
        RECT 1435.020 -28.120 1438.020 0.300 ;
        RECT 1525.020 -28.120 1528.020 0.300 ;
        RECT 1615.020 -28.120 1618.020 0.300 ;
        RECT 1705.020 -28.120 1708.020 0.300 ;
        RECT 1795.020 -28.120 1798.020 0.300 ;
        RECT 1885.020 -28.120 1888.020 0.300 ;
        RECT 1975.020 -28.120 1978.020 0.300 ;
        RECT 2065.020 -28.120 2068.020 0.300 ;
        RECT 2155.020 -28.120 2158.020 0.300 ;
        RECT 2245.020 -28.120 2248.020 0.300 ;
        RECT 2335.020 -28.120 2338.020 0.300 ;
        RECT 2425.020 -28.120 2428.020 0.300 ;
        RECT 2515.020 -28.120 2518.020 0.300 ;
        RECT 2605.020 -28.120 2608.020 0.300 ;
        RECT 2695.020 -28.120 2698.020 0.300 ;
        RECT 2785.020 -28.120 2788.020 0.300 ;
        RECT 2875.020 -28.120 2878.020 0.300 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 85.930 3546.510 87.110 3547.690 ;
        RECT 85.930 3544.910 87.110 3546.090 ;
        RECT 175.930 3546.510 177.110 3547.690 ;
        RECT 175.930 3544.910 177.110 3546.090 ;
        RECT 265.930 3546.510 267.110 3547.690 ;
        RECT 265.930 3544.910 267.110 3546.090 ;
        RECT 355.930 3546.510 357.110 3547.690 ;
        RECT 355.930 3544.910 357.110 3546.090 ;
        RECT 445.930 3546.510 447.110 3547.690 ;
        RECT 445.930 3544.910 447.110 3546.090 ;
        RECT 535.930 3546.510 537.110 3547.690 ;
        RECT 535.930 3544.910 537.110 3546.090 ;
        RECT 625.930 3546.510 627.110 3547.690 ;
        RECT 625.930 3544.910 627.110 3546.090 ;
        RECT 715.930 3546.510 717.110 3547.690 ;
        RECT 715.930 3544.910 717.110 3546.090 ;
        RECT 805.930 3546.510 807.110 3547.690 ;
        RECT 805.930 3544.910 807.110 3546.090 ;
        RECT 895.930 3546.510 897.110 3547.690 ;
        RECT 895.930 3544.910 897.110 3546.090 ;
        RECT 985.930 3546.510 987.110 3547.690 ;
        RECT 985.930 3544.910 987.110 3546.090 ;
        RECT 1075.930 3546.510 1077.110 3547.690 ;
        RECT 1075.930 3544.910 1077.110 3546.090 ;
        RECT 1165.930 3546.510 1167.110 3547.690 ;
        RECT 1165.930 3544.910 1167.110 3546.090 ;
        RECT 1255.930 3546.510 1257.110 3547.690 ;
        RECT 1255.930 3544.910 1257.110 3546.090 ;
        RECT 1345.930 3546.510 1347.110 3547.690 ;
        RECT 1345.930 3544.910 1347.110 3546.090 ;
        RECT 1435.930 3546.510 1437.110 3547.690 ;
        RECT 1435.930 3544.910 1437.110 3546.090 ;
        RECT 1525.930 3546.510 1527.110 3547.690 ;
        RECT 1525.930 3544.910 1527.110 3546.090 ;
        RECT 1615.930 3546.510 1617.110 3547.690 ;
        RECT 1615.930 3544.910 1617.110 3546.090 ;
        RECT 1705.930 3546.510 1707.110 3547.690 ;
        RECT 1705.930 3544.910 1707.110 3546.090 ;
        RECT 1795.930 3546.510 1797.110 3547.690 ;
        RECT 1795.930 3544.910 1797.110 3546.090 ;
        RECT 1885.930 3546.510 1887.110 3547.690 ;
        RECT 1885.930 3544.910 1887.110 3546.090 ;
        RECT 1975.930 3546.510 1977.110 3547.690 ;
        RECT 1975.930 3544.910 1977.110 3546.090 ;
        RECT 2065.930 3546.510 2067.110 3547.690 ;
        RECT 2065.930 3544.910 2067.110 3546.090 ;
        RECT 2155.930 3546.510 2157.110 3547.690 ;
        RECT 2155.930 3544.910 2157.110 3546.090 ;
        RECT 2245.930 3546.510 2247.110 3547.690 ;
        RECT 2245.930 3544.910 2247.110 3546.090 ;
        RECT 2335.930 3546.510 2337.110 3547.690 ;
        RECT 2335.930 3544.910 2337.110 3546.090 ;
        RECT 2425.930 3546.510 2427.110 3547.690 ;
        RECT 2425.930 3544.910 2427.110 3546.090 ;
        RECT 2515.930 3546.510 2517.110 3547.690 ;
        RECT 2515.930 3544.910 2517.110 3546.090 ;
        RECT 2605.930 3546.510 2607.110 3547.690 ;
        RECT 2605.930 3544.910 2607.110 3546.090 ;
        RECT 2695.930 3546.510 2697.110 3547.690 ;
        RECT 2695.930 3544.910 2697.110 3546.090 ;
        RECT 2785.930 3546.510 2787.110 3547.690 ;
        RECT 2785.930 3544.910 2787.110 3546.090 ;
        RECT 2875.930 3546.510 2877.110 3547.690 ;
        RECT 2875.930 3544.910 2877.110 3546.090 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT -32.570 3422.090 -31.390 3423.270 ;
        RECT -32.570 3420.490 -31.390 3421.670 ;
        RECT -32.570 3332.090 -31.390 3333.270 ;
        RECT -32.570 3330.490 -31.390 3331.670 ;
        RECT -32.570 3242.090 -31.390 3243.270 ;
        RECT -32.570 3240.490 -31.390 3241.670 ;
        RECT -32.570 3152.090 -31.390 3153.270 ;
        RECT -32.570 3150.490 -31.390 3151.670 ;
        RECT -32.570 3062.090 -31.390 3063.270 ;
        RECT -32.570 3060.490 -31.390 3061.670 ;
        RECT -32.570 2972.090 -31.390 2973.270 ;
        RECT -32.570 2970.490 -31.390 2971.670 ;
        RECT -32.570 2882.090 -31.390 2883.270 ;
        RECT -32.570 2880.490 -31.390 2881.670 ;
        RECT -32.570 2792.090 -31.390 2793.270 ;
        RECT -32.570 2790.490 -31.390 2791.670 ;
        RECT -32.570 2702.090 -31.390 2703.270 ;
        RECT -32.570 2700.490 -31.390 2701.670 ;
        RECT -32.570 2612.090 -31.390 2613.270 ;
        RECT -32.570 2610.490 -31.390 2611.670 ;
        RECT -32.570 2522.090 -31.390 2523.270 ;
        RECT -32.570 2520.490 -31.390 2521.670 ;
        RECT -32.570 2432.090 -31.390 2433.270 ;
        RECT -32.570 2430.490 -31.390 2431.670 ;
        RECT -32.570 2342.090 -31.390 2343.270 ;
        RECT -32.570 2340.490 -31.390 2341.670 ;
        RECT -32.570 2252.090 -31.390 2253.270 ;
        RECT -32.570 2250.490 -31.390 2251.670 ;
        RECT -32.570 2162.090 -31.390 2163.270 ;
        RECT -32.570 2160.490 -31.390 2161.670 ;
        RECT -32.570 2072.090 -31.390 2073.270 ;
        RECT -32.570 2070.490 -31.390 2071.670 ;
        RECT -32.570 1982.090 -31.390 1983.270 ;
        RECT -32.570 1980.490 -31.390 1981.670 ;
        RECT -32.570 1892.090 -31.390 1893.270 ;
        RECT -32.570 1890.490 -31.390 1891.670 ;
        RECT -32.570 1802.090 -31.390 1803.270 ;
        RECT -32.570 1800.490 -31.390 1801.670 ;
        RECT -32.570 1712.090 -31.390 1713.270 ;
        RECT -32.570 1710.490 -31.390 1711.670 ;
        RECT -32.570 1622.090 -31.390 1623.270 ;
        RECT -32.570 1620.490 -31.390 1621.670 ;
        RECT -32.570 1532.090 -31.390 1533.270 ;
        RECT -32.570 1530.490 -31.390 1531.670 ;
        RECT -32.570 1442.090 -31.390 1443.270 ;
        RECT -32.570 1440.490 -31.390 1441.670 ;
        RECT -32.570 1352.090 -31.390 1353.270 ;
        RECT -32.570 1350.490 -31.390 1351.670 ;
        RECT -32.570 1262.090 -31.390 1263.270 ;
        RECT -32.570 1260.490 -31.390 1261.670 ;
        RECT -32.570 1172.090 -31.390 1173.270 ;
        RECT -32.570 1170.490 -31.390 1171.670 ;
        RECT -32.570 1082.090 -31.390 1083.270 ;
        RECT -32.570 1080.490 -31.390 1081.670 ;
        RECT -32.570 992.090 -31.390 993.270 ;
        RECT -32.570 990.490 -31.390 991.670 ;
        RECT -32.570 902.090 -31.390 903.270 ;
        RECT -32.570 900.490 -31.390 901.670 ;
        RECT -32.570 812.090 -31.390 813.270 ;
        RECT -32.570 810.490 -31.390 811.670 ;
        RECT -32.570 722.090 -31.390 723.270 ;
        RECT -32.570 720.490 -31.390 721.670 ;
        RECT -32.570 632.090 -31.390 633.270 ;
        RECT -32.570 630.490 -31.390 631.670 ;
        RECT -32.570 542.090 -31.390 543.270 ;
        RECT -32.570 540.490 -31.390 541.670 ;
        RECT -32.570 452.090 -31.390 453.270 ;
        RECT -32.570 450.490 -31.390 451.670 ;
        RECT -32.570 362.090 -31.390 363.270 ;
        RECT -32.570 360.490 -31.390 361.670 ;
        RECT -32.570 272.090 -31.390 273.270 ;
        RECT -32.570 270.490 -31.390 271.670 ;
        RECT -32.570 182.090 -31.390 183.270 ;
        RECT -32.570 180.490 -31.390 181.670 ;
        RECT -32.570 92.090 -31.390 93.270 ;
        RECT -32.570 90.490 -31.390 91.670 ;
        RECT 2951.010 3422.090 2952.190 3423.270 ;
        RECT 2951.010 3420.490 2952.190 3421.670 ;
        RECT 2951.010 3332.090 2952.190 3333.270 ;
        RECT 2951.010 3330.490 2952.190 3331.670 ;
        RECT 2951.010 3242.090 2952.190 3243.270 ;
        RECT 2951.010 3240.490 2952.190 3241.670 ;
        RECT 2951.010 3152.090 2952.190 3153.270 ;
        RECT 2951.010 3150.490 2952.190 3151.670 ;
        RECT 2951.010 3062.090 2952.190 3063.270 ;
        RECT 2951.010 3060.490 2952.190 3061.670 ;
        RECT 2951.010 2972.090 2952.190 2973.270 ;
        RECT 2951.010 2970.490 2952.190 2971.670 ;
        RECT 2951.010 2882.090 2952.190 2883.270 ;
        RECT 2951.010 2880.490 2952.190 2881.670 ;
        RECT 2951.010 2792.090 2952.190 2793.270 ;
        RECT 2951.010 2790.490 2952.190 2791.670 ;
        RECT 2951.010 2702.090 2952.190 2703.270 ;
        RECT 2951.010 2700.490 2952.190 2701.670 ;
        RECT 2951.010 2612.090 2952.190 2613.270 ;
        RECT 2951.010 2610.490 2952.190 2611.670 ;
        RECT 2951.010 2522.090 2952.190 2523.270 ;
        RECT 2951.010 2520.490 2952.190 2521.670 ;
        RECT 2951.010 2432.090 2952.190 2433.270 ;
        RECT 2951.010 2430.490 2952.190 2431.670 ;
        RECT 2951.010 2342.090 2952.190 2343.270 ;
        RECT 2951.010 2340.490 2952.190 2341.670 ;
        RECT 2951.010 2252.090 2952.190 2253.270 ;
        RECT 2951.010 2250.490 2952.190 2251.670 ;
        RECT 2951.010 2162.090 2952.190 2163.270 ;
        RECT 2951.010 2160.490 2952.190 2161.670 ;
        RECT 2951.010 2072.090 2952.190 2073.270 ;
        RECT 2951.010 2070.490 2952.190 2071.670 ;
        RECT 2951.010 1982.090 2952.190 1983.270 ;
        RECT 2951.010 1980.490 2952.190 1981.670 ;
        RECT 2951.010 1892.090 2952.190 1893.270 ;
        RECT 2951.010 1890.490 2952.190 1891.670 ;
        RECT 2951.010 1802.090 2952.190 1803.270 ;
        RECT 2951.010 1800.490 2952.190 1801.670 ;
        RECT 2951.010 1712.090 2952.190 1713.270 ;
        RECT 2951.010 1710.490 2952.190 1711.670 ;
        RECT 2951.010 1622.090 2952.190 1623.270 ;
        RECT 2951.010 1620.490 2952.190 1621.670 ;
        RECT 2951.010 1532.090 2952.190 1533.270 ;
        RECT 2951.010 1530.490 2952.190 1531.670 ;
        RECT 2951.010 1442.090 2952.190 1443.270 ;
        RECT 2951.010 1440.490 2952.190 1441.670 ;
        RECT 2951.010 1352.090 2952.190 1353.270 ;
        RECT 2951.010 1350.490 2952.190 1351.670 ;
        RECT 2951.010 1262.090 2952.190 1263.270 ;
        RECT 2951.010 1260.490 2952.190 1261.670 ;
        RECT 2951.010 1172.090 2952.190 1173.270 ;
        RECT 2951.010 1170.490 2952.190 1171.670 ;
        RECT 2951.010 1082.090 2952.190 1083.270 ;
        RECT 2951.010 1080.490 2952.190 1081.670 ;
        RECT 2951.010 992.090 2952.190 993.270 ;
        RECT 2951.010 990.490 2952.190 991.670 ;
        RECT 2951.010 902.090 2952.190 903.270 ;
        RECT 2951.010 900.490 2952.190 901.670 ;
        RECT 2951.010 812.090 2952.190 813.270 ;
        RECT 2951.010 810.490 2952.190 811.670 ;
        RECT 2951.010 722.090 2952.190 723.270 ;
        RECT 2951.010 720.490 2952.190 721.670 ;
        RECT 2951.010 632.090 2952.190 633.270 ;
        RECT 2951.010 630.490 2952.190 631.670 ;
        RECT 2951.010 542.090 2952.190 543.270 ;
        RECT 2951.010 540.490 2952.190 541.670 ;
        RECT 2951.010 452.090 2952.190 453.270 ;
        RECT 2951.010 450.490 2952.190 451.670 ;
        RECT 2951.010 362.090 2952.190 363.270 ;
        RECT 2951.010 360.490 2952.190 361.670 ;
        RECT 2951.010 272.090 2952.190 273.270 ;
        RECT 2951.010 270.490 2952.190 271.670 ;
        RECT 2951.010 182.090 2952.190 183.270 ;
        RECT 2951.010 180.490 2952.190 181.670 ;
        RECT 2951.010 92.090 2952.190 93.270 ;
        RECT 2951.010 90.490 2952.190 91.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 85.930 -26.410 87.110 -25.230 ;
        RECT 85.930 -28.010 87.110 -26.830 ;
        RECT 175.930 -26.410 177.110 -25.230 ;
        RECT 175.930 -28.010 177.110 -26.830 ;
        RECT 265.930 -26.410 267.110 -25.230 ;
        RECT 265.930 -28.010 267.110 -26.830 ;
        RECT 355.930 -26.410 357.110 -25.230 ;
        RECT 355.930 -28.010 357.110 -26.830 ;
        RECT 445.930 -26.410 447.110 -25.230 ;
        RECT 445.930 -28.010 447.110 -26.830 ;
        RECT 535.930 -26.410 537.110 -25.230 ;
        RECT 535.930 -28.010 537.110 -26.830 ;
        RECT 625.930 -26.410 627.110 -25.230 ;
        RECT 625.930 -28.010 627.110 -26.830 ;
        RECT 715.930 -26.410 717.110 -25.230 ;
        RECT 715.930 -28.010 717.110 -26.830 ;
        RECT 805.930 -26.410 807.110 -25.230 ;
        RECT 805.930 -28.010 807.110 -26.830 ;
        RECT 895.930 -26.410 897.110 -25.230 ;
        RECT 895.930 -28.010 897.110 -26.830 ;
        RECT 985.930 -26.410 987.110 -25.230 ;
        RECT 985.930 -28.010 987.110 -26.830 ;
        RECT 1075.930 -26.410 1077.110 -25.230 ;
        RECT 1075.930 -28.010 1077.110 -26.830 ;
        RECT 1165.930 -26.410 1167.110 -25.230 ;
        RECT 1165.930 -28.010 1167.110 -26.830 ;
        RECT 1255.930 -26.410 1257.110 -25.230 ;
        RECT 1255.930 -28.010 1257.110 -26.830 ;
        RECT 1345.930 -26.410 1347.110 -25.230 ;
        RECT 1345.930 -28.010 1347.110 -26.830 ;
        RECT 1435.930 -26.410 1437.110 -25.230 ;
        RECT 1435.930 -28.010 1437.110 -26.830 ;
        RECT 1525.930 -26.410 1527.110 -25.230 ;
        RECT 1525.930 -28.010 1527.110 -26.830 ;
        RECT 1615.930 -26.410 1617.110 -25.230 ;
        RECT 1615.930 -28.010 1617.110 -26.830 ;
        RECT 1705.930 -26.410 1707.110 -25.230 ;
        RECT 1705.930 -28.010 1707.110 -26.830 ;
        RECT 1795.930 -26.410 1797.110 -25.230 ;
        RECT 1795.930 -28.010 1797.110 -26.830 ;
        RECT 1885.930 -26.410 1887.110 -25.230 ;
        RECT 1885.930 -28.010 1887.110 -26.830 ;
        RECT 1975.930 -26.410 1977.110 -25.230 ;
        RECT 1975.930 -28.010 1977.110 -26.830 ;
        RECT 2065.930 -26.410 2067.110 -25.230 ;
        RECT 2065.930 -28.010 2067.110 -26.830 ;
        RECT 2155.930 -26.410 2157.110 -25.230 ;
        RECT 2155.930 -28.010 2157.110 -26.830 ;
        RECT 2245.930 -26.410 2247.110 -25.230 ;
        RECT 2245.930 -28.010 2247.110 -26.830 ;
        RECT 2335.930 -26.410 2337.110 -25.230 ;
        RECT 2335.930 -28.010 2337.110 -26.830 ;
        RECT 2425.930 -26.410 2427.110 -25.230 ;
        RECT 2425.930 -28.010 2427.110 -26.830 ;
        RECT 2515.930 -26.410 2517.110 -25.230 ;
        RECT 2515.930 -28.010 2517.110 -26.830 ;
        RECT 2605.930 -26.410 2607.110 -25.230 ;
        RECT 2605.930 -28.010 2607.110 -26.830 ;
        RECT 2695.930 -26.410 2697.110 -25.230 ;
        RECT 2695.930 -28.010 2697.110 -26.830 ;
        RECT 2785.930 -26.410 2787.110 -25.230 ;
        RECT 2785.930 -28.010 2787.110 -26.830 ;
        RECT 2875.930 -26.410 2877.110 -25.230 ;
        RECT 2875.930 -28.010 2877.110 -26.830 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 85.020 3547.800 88.020 3547.810 ;
        RECT 175.020 3547.800 178.020 3547.810 ;
        RECT 265.020 3547.800 268.020 3547.810 ;
        RECT 355.020 3547.800 358.020 3547.810 ;
        RECT 445.020 3547.800 448.020 3547.810 ;
        RECT 535.020 3547.800 538.020 3547.810 ;
        RECT 625.020 3547.800 628.020 3547.810 ;
        RECT 715.020 3547.800 718.020 3547.810 ;
        RECT 805.020 3547.800 808.020 3547.810 ;
        RECT 895.020 3547.800 898.020 3547.810 ;
        RECT 985.020 3547.800 988.020 3547.810 ;
        RECT 1075.020 3547.800 1078.020 3547.810 ;
        RECT 1165.020 3547.800 1168.020 3547.810 ;
        RECT 1255.020 3547.800 1258.020 3547.810 ;
        RECT 1345.020 3547.800 1348.020 3547.810 ;
        RECT 1435.020 3547.800 1438.020 3547.810 ;
        RECT 1525.020 3547.800 1528.020 3547.810 ;
        RECT 1615.020 3547.800 1618.020 3547.810 ;
        RECT 1705.020 3547.800 1708.020 3547.810 ;
        RECT 1795.020 3547.800 1798.020 3547.810 ;
        RECT 1885.020 3547.800 1888.020 3547.810 ;
        RECT 1975.020 3547.800 1978.020 3547.810 ;
        RECT 2065.020 3547.800 2068.020 3547.810 ;
        RECT 2155.020 3547.800 2158.020 3547.810 ;
        RECT 2245.020 3547.800 2248.020 3547.810 ;
        RECT 2335.020 3547.800 2338.020 3547.810 ;
        RECT 2425.020 3547.800 2428.020 3547.810 ;
        RECT 2515.020 3547.800 2518.020 3547.810 ;
        RECT 2605.020 3547.800 2608.020 3547.810 ;
        RECT 2695.020 3547.800 2698.020 3547.810 ;
        RECT 2785.020 3547.800 2788.020 3547.810 ;
        RECT 2875.020 3547.800 2878.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 85.020 3544.790 88.020 3544.800 ;
        RECT 175.020 3544.790 178.020 3544.800 ;
        RECT 265.020 3544.790 268.020 3544.800 ;
        RECT 355.020 3544.790 358.020 3544.800 ;
        RECT 445.020 3544.790 448.020 3544.800 ;
        RECT 535.020 3544.790 538.020 3544.800 ;
        RECT 625.020 3544.790 628.020 3544.800 ;
        RECT 715.020 3544.790 718.020 3544.800 ;
        RECT 805.020 3544.790 808.020 3544.800 ;
        RECT 895.020 3544.790 898.020 3544.800 ;
        RECT 985.020 3544.790 988.020 3544.800 ;
        RECT 1075.020 3544.790 1078.020 3544.800 ;
        RECT 1165.020 3544.790 1168.020 3544.800 ;
        RECT 1255.020 3544.790 1258.020 3544.800 ;
        RECT 1345.020 3544.790 1348.020 3544.800 ;
        RECT 1435.020 3544.790 1438.020 3544.800 ;
        RECT 1525.020 3544.790 1528.020 3544.800 ;
        RECT 1615.020 3544.790 1618.020 3544.800 ;
        RECT 1705.020 3544.790 1708.020 3544.800 ;
        RECT 1795.020 3544.790 1798.020 3544.800 ;
        RECT 1885.020 3544.790 1888.020 3544.800 ;
        RECT 1975.020 3544.790 1978.020 3544.800 ;
        RECT 2065.020 3544.790 2068.020 3544.800 ;
        RECT 2155.020 3544.790 2158.020 3544.800 ;
        RECT 2245.020 3544.790 2248.020 3544.800 ;
        RECT 2335.020 3544.790 2338.020 3544.800 ;
        RECT 2425.020 3544.790 2428.020 3544.800 ;
        RECT 2515.020 3544.790 2518.020 3544.800 ;
        RECT 2605.020 3544.790 2608.020 3544.800 ;
        RECT 2695.020 3544.790 2698.020 3544.800 ;
        RECT 2785.020 3544.790 2788.020 3544.800 ;
        RECT 2875.020 3544.790 2878.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3423.380 -30.480 3423.390 ;
        RECT 2950.100 3423.380 2953.100 3423.390 ;
        RECT -33.480 3420.380 0.300 3423.380 ;
        RECT 2919.700 3420.380 2953.100 3423.380 ;
        RECT -33.480 3420.370 -30.480 3420.380 ;
        RECT 2950.100 3420.370 2953.100 3420.380 ;
        RECT -33.480 3333.380 -30.480 3333.390 ;
        RECT 2950.100 3333.380 2953.100 3333.390 ;
        RECT -33.480 3330.380 0.300 3333.380 ;
        RECT 2919.700 3330.380 2953.100 3333.380 ;
        RECT -33.480 3330.370 -30.480 3330.380 ;
        RECT 2950.100 3330.370 2953.100 3330.380 ;
        RECT -33.480 3243.380 -30.480 3243.390 ;
        RECT 2950.100 3243.380 2953.100 3243.390 ;
        RECT -33.480 3240.380 0.300 3243.380 ;
        RECT 2919.700 3240.380 2953.100 3243.380 ;
        RECT -33.480 3240.370 -30.480 3240.380 ;
        RECT 2950.100 3240.370 2953.100 3240.380 ;
        RECT -33.480 3153.380 -30.480 3153.390 ;
        RECT 2950.100 3153.380 2953.100 3153.390 ;
        RECT -33.480 3150.380 0.300 3153.380 ;
        RECT 2919.700 3150.380 2953.100 3153.380 ;
        RECT -33.480 3150.370 -30.480 3150.380 ;
        RECT 2950.100 3150.370 2953.100 3150.380 ;
        RECT -33.480 3063.380 -30.480 3063.390 ;
        RECT 2950.100 3063.380 2953.100 3063.390 ;
        RECT -33.480 3060.380 0.300 3063.380 ;
        RECT 2919.700 3060.380 2953.100 3063.380 ;
        RECT -33.480 3060.370 -30.480 3060.380 ;
        RECT 2950.100 3060.370 2953.100 3060.380 ;
        RECT -33.480 2973.380 -30.480 2973.390 ;
        RECT 2950.100 2973.380 2953.100 2973.390 ;
        RECT -33.480 2970.380 0.300 2973.380 ;
        RECT 2919.700 2970.380 2953.100 2973.380 ;
        RECT -33.480 2970.370 -30.480 2970.380 ;
        RECT 2950.100 2970.370 2953.100 2970.380 ;
        RECT -33.480 2883.380 -30.480 2883.390 ;
        RECT 2950.100 2883.380 2953.100 2883.390 ;
        RECT -33.480 2880.380 0.300 2883.380 ;
        RECT 2919.700 2880.380 2953.100 2883.380 ;
        RECT -33.480 2880.370 -30.480 2880.380 ;
        RECT 2950.100 2880.370 2953.100 2880.380 ;
        RECT -33.480 2793.380 -30.480 2793.390 ;
        RECT 2950.100 2793.380 2953.100 2793.390 ;
        RECT -33.480 2790.380 0.300 2793.380 ;
        RECT 2919.700 2790.380 2953.100 2793.380 ;
        RECT -33.480 2790.370 -30.480 2790.380 ;
        RECT 2950.100 2790.370 2953.100 2790.380 ;
        RECT -33.480 2703.380 -30.480 2703.390 ;
        RECT 2950.100 2703.380 2953.100 2703.390 ;
        RECT -33.480 2700.380 0.300 2703.380 ;
        RECT 2919.700 2700.380 2953.100 2703.380 ;
        RECT -33.480 2700.370 -30.480 2700.380 ;
        RECT 2950.100 2700.370 2953.100 2700.380 ;
        RECT -33.480 2613.380 -30.480 2613.390 ;
        RECT 2950.100 2613.380 2953.100 2613.390 ;
        RECT -33.480 2610.380 0.300 2613.380 ;
        RECT 2919.700 2610.380 2953.100 2613.380 ;
        RECT -33.480 2610.370 -30.480 2610.380 ;
        RECT 2950.100 2610.370 2953.100 2610.380 ;
        RECT -33.480 2523.380 -30.480 2523.390 ;
        RECT 2950.100 2523.380 2953.100 2523.390 ;
        RECT -33.480 2520.380 0.300 2523.380 ;
        RECT 2919.700 2520.380 2953.100 2523.380 ;
        RECT -33.480 2520.370 -30.480 2520.380 ;
        RECT 2950.100 2520.370 2953.100 2520.380 ;
        RECT -33.480 2433.380 -30.480 2433.390 ;
        RECT 2950.100 2433.380 2953.100 2433.390 ;
        RECT -33.480 2430.380 0.300 2433.380 ;
        RECT 2919.700 2430.380 2953.100 2433.380 ;
        RECT -33.480 2430.370 -30.480 2430.380 ;
        RECT 2950.100 2430.370 2953.100 2430.380 ;
        RECT -33.480 2343.380 -30.480 2343.390 ;
        RECT 2950.100 2343.380 2953.100 2343.390 ;
        RECT -33.480 2340.380 0.300 2343.380 ;
        RECT 2919.700 2340.380 2953.100 2343.380 ;
        RECT -33.480 2340.370 -30.480 2340.380 ;
        RECT 2950.100 2340.370 2953.100 2340.380 ;
        RECT -33.480 2253.380 -30.480 2253.390 ;
        RECT 2950.100 2253.380 2953.100 2253.390 ;
        RECT -33.480 2250.380 0.300 2253.380 ;
        RECT 2919.700 2250.380 2953.100 2253.380 ;
        RECT -33.480 2250.370 -30.480 2250.380 ;
        RECT 2950.100 2250.370 2953.100 2250.380 ;
        RECT -33.480 2163.380 -30.480 2163.390 ;
        RECT 2950.100 2163.380 2953.100 2163.390 ;
        RECT -33.480 2160.380 0.300 2163.380 ;
        RECT 2919.700 2160.380 2953.100 2163.380 ;
        RECT -33.480 2160.370 -30.480 2160.380 ;
        RECT 2950.100 2160.370 2953.100 2160.380 ;
        RECT -33.480 2073.380 -30.480 2073.390 ;
        RECT 2950.100 2073.380 2953.100 2073.390 ;
        RECT -33.480 2070.380 0.300 2073.380 ;
        RECT 2919.700 2070.380 2953.100 2073.380 ;
        RECT -33.480 2070.370 -30.480 2070.380 ;
        RECT 2950.100 2070.370 2953.100 2070.380 ;
        RECT -33.480 1983.380 -30.480 1983.390 ;
        RECT 2950.100 1983.380 2953.100 1983.390 ;
        RECT -33.480 1980.380 0.300 1983.380 ;
        RECT 2919.700 1980.380 2953.100 1983.380 ;
        RECT -33.480 1980.370 -30.480 1980.380 ;
        RECT 2950.100 1980.370 2953.100 1980.380 ;
        RECT -33.480 1893.380 -30.480 1893.390 ;
        RECT 2950.100 1893.380 2953.100 1893.390 ;
        RECT -33.480 1890.380 0.300 1893.380 ;
        RECT 2919.700 1890.380 2953.100 1893.380 ;
        RECT -33.480 1890.370 -30.480 1890.380 ;
        RECT 2950.100 1890.370 2953.100 1890.380 ;
        RECT -33.480 1803.380 -30.480 1803.390 ;
        RECT 2950.100 1803.380 2953.100 1803.390 ;
        RECT -33.480 1800.380 0.300 1803.380 ;
        RECT 2919.700 1800.380 2953.100 1803.380 ;
        RECT -33.480 1800.370 -30.480 1800.380 ;
        RECT 2950.100 1800.370 2953.100 1800.380 ;
        RECT -33.480 1713.380 -30.480 1713.390 ;
        RECT 2950.100 1713.380 2953.100 1713.390 ;
        RECT -33.480 1710.380 0.300 1713.380 ;
        RECT 2919.700 1710.380 2953.100 1713.380 ;
        RECT -33.480 1710.370 -30.480 1710.380 ;
        RECT 2950.100 1710.370 2953.100 1710.380 ;
        RECT -33.480 1623.380 -30.480 1623.390 ;
        RECT 2950.100 1623.380 2953.100 1623.390 ;
        RECT -33.480 1620.380 0.300 1623.380 ;
        RECT 2919.700 1620.380 2953.100 1623.380 ;
        RECT -33.480 1620.370 -30.480 1620.380 ;
        RECT 2950.100 1620.370 2953.100 1620.380 ;
        RECT -33.480 1533.380 -30.480 1533.390 ;
        RECT 2950.100 1533.380 2953.100 1533.390 ;
        RECT -33.480 1530.380 0.300 1533.380 ;
        RECT 2919.700 1530.380 2953.100 1533.380 ;
        RECT -33.480 1530.370 -30.480 1530.380 ;
        RECT 2950.100 1530.370 2953.100 1530.380 ;
        RECT -33.480 1443.380 -30.480 1443.390 ;
        RECT 2950.100 1443.380 2953.100 1443.390 ;
        RECT -33.480 1440.380 0.300 1443.380 ;
        RECT 2919.700 1440.380 2953.100 1443.380 ;
        RECT -33.480 1440.370 -30.480 1440.380 ;
        RECT 2950.100 1440.370 2953.100 1440.380 ;
        RECT -33.480 1353.380 -30.480 1353.390 ;
        RECT 2950.100 1353.380 2953.100 1353.390 ;
        RECT -33.480 1350.380 0.300 1353.380 ;
        RECT 2919.700 1350.380 2953.100 1353.380 ;
        RECT -33.480 1350.370 -30.480 1350.380 ;
        RECT 2950.100 1350.370 2953.100 1350.380 ;
        RECT -33.480 1263.380 -30.480 1263.390 ;
        RECT 2950.100 1263.380 2953.100 1263.390 ;
        RECT -33.480 1260.380 0.300 1263.380 ;
        RECT 2919.700 1260.380 2953.100 1263.380 ;
        RECT -33.480 1260.370 -30.480 1260.380 ;
        RECT 2950.100 1260.370 2953.100 1260.380 ;
        RECT -33.480 1173.380 -30.480 1173.390 ;
        RECT 2950.100 1173.380 2953.100 1173.390 ;
        RECT -33.480 1170.380 0.300 1173.380 ;
        RECT 2919.700 1170.380 2953.100 1173.380 ;
        RECT -33.480 1170.370 -30.480 1170.380 ;
        RECT 2950.100 1170.370 2953.100 1170.380 ;
        RECT -33.480 1083.380 -30.480 1083.390 ;
        RECT 2950.100 1083.380 2953.100 1083.390 ;
        RECT -33.480 1080.380 0.300 1083.380 ;
        RECT 2919.700 1080.380 2953.100 1083.380 ;
        RECT -33.480 1080.370 -30.480 1080.380 ;
        RECT 2950.100 1080.370 2953.100 1080.380 ;
        RECT -33.480 993.380 -30.480 993.390 ;
        RECT 2950.100 993.380 2953.100 993.390 ;
        RECT -33.480 990.380 0.300 993.380 ;
        RECT 2919.700 990.380 2953.100 993.380 ;
        RECT -33.480 990.370 -30.480 990.380 ;
        RECT 2950.100 990.370 2953.100 990.380 ;
        RECT -33.480 903.380 -30.480 903.390 ;
        RECT 2950.100 903.380 2953.100 903.390 ;
        RECT -33.480 900.380 0.300 903.380 ;
        RECT 2919.700 900.380 2953.100 903.380 ;
        RECT -33.480 900.370 -30.480 900.380 ;
        RECT 2950.100 900.370 2953.100 900.380 ;
        RECT -33.480 813.380 -30.480 813.390 ;
        RECT 2950.100 813.380 2953.100 813.390 ;
        RECT -33.480 810.380 0.300 813.380 ;
        RECT 2919.700 810.380 2953.100 813.380 ;
        RECT -33.480 810.370 -30.480 810.380 ;
        RECT 2950.100 810.370 2953.100 810.380 ;
        RECT -33.480 723.380 -30.480 723.390 ;
        RECT 2950.100 723.380 2953.100 723.390 ;
        RECT -33.480 720.380 0.300 723.380 ;
        RECT 2919.700 720.380 2953.100 723.380 ;
        RECT -33.480 720.370 -30.480 720.380 ;
        RECT 2950.100 720.370 2953.100 720.380 ;
        RECT -33.480 633.380 -30.480 633.390 ;
        RECT 2950.100 633.380 2953.100 633.390 ;
        RECT -33.480 630.380 0.300 633.380 ;
        RECT 2919.700 630.380 2953.100 633.380 ;
        RECT -33.480 630.370 -30.480 630.380 ;
        RECT 2950.100 630.370 2953.100 630.380 ;
        RECT -33.480 543.380 -30.480 543.390 ;
        RECT 2950.100 543.380 2953.100 543.390 ;
        RECT -33.480 540.380 0.300 543.380 ;
        RECT 2919.700 540.380 2953.100 543.380 ;
        RECT -33.480 540.370 -30.480 540.380 ;
        RECT 2950.100 540.370 2953.100 540.380 ;
        RECT -33.480 453.380 -30.480 453.390 ;
        RECT 2950.100 453.380 2953.100 453.390 ;
        RECT -33.480 450.380 0.300 453.380 ;
        RECT 2919.700 450.380 2953.100 453.380 ;
        RECT -33.480 450.370 -30.480 450.380 ;
        RECT 2950.100 450.370 2953.100 450.380 ;
        RECT -33.480 363.380 -30.480 363.390 ;
        RECT 2950.100 363.380 2953.100 363.390 ;
        RECT -33.480 360.380 0.300 363.380 ;
        RECT 2919.700 360.380 2953.100 363.380 ;
        RECT -33.480 360.370 -30.480 360.380 ;
        RECT 2950.100 360.370 2953.100 360.380 ;
        RECT -33.480 273.380 -30.480 273.390 ;
        RECT 2950.100 273.380 2953.100 273.390 ;
        RECT -33.480 270.380 0.300 273.380 ;
        RECT 2919.700 270.380 2953.100 273.380 ;
        RECT -33.480 270.370 -30.480 270.380 ;
        RECT 2950.100 270.370 2953.100 270.380 ;
        RECT -33.480 183.380 -30.480 183.390 ;
        RECT 2950.100 183.380 2953.100 183.390 ;
        RECT -33.480 180.380 0.300 183.380 ;
        RECT 2919.700 180.380 2953.100 183.380 ;
        RECT -33.480 180.370 -30.480 180.380 ;
        RECT 2950.100 180.370 2953.100 180.380 ;
        RECT -33.480 93.380 -30.480 93.390 ;
        RECT 2950.100 93.380 2953.100 93.390 ;
        RECT -33.480 90.380 0.300 93.380 ;
        RECT 2919.700 90.380 2953.100 93.380 ;
        RECT -33.480 90.370 -30.480 90.380 ;
        RECT 2950.100 90.370 2953.100 90.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 85.020 -25.120 88.020 -25.110 ;
        RECT 175.020 -25.120 178.020 -25.110 ;
        RECT 265.020 -25.120 268.020 -25.110 ;
        RECT 355.020 -25.120 358.020 -25.110 ;
        RECT 445.020 -25.120 448.020 -25.110 ;
        RECT 535.020 -25.120 538.020 -25.110 ;
        RECT 625.020 -25.120 628.020 -25.110 ;
        RECT 715.020 -25.120 718.020 -25.110 ;
        RECT 805.020 -25.120 808.020 -25.110 ;
        RECT 895.020 -25.120 898.020 -25.110 ;
        RECT 985.020 -25.120 988.020 -25.110 ;
        RECT 1075.020 -25.120 1078.020 -25.110 ;
        RECT 1165.020 -25.120 1168.020 -25.110 ;
        RECT 1255.020 -25.120 1258.020 -25.110 ;
        RECT 1345.020 -25.120 1348.020 -25.110 ;
        RECT 1435.020 -25.120 1438.020 -25.110 ;
        RECT 1525.020 -25.120 1528.020 -25.110 ;
        RECT 1615.020 -25.120 1618.020 -25.110 ;
        RECT 1705.020 -25.120 1708.020 -25.110 ;
        RECT 1795.020 -25.120 1798.020 -25.110 ;
        RECT 1885.020 -25.120 1888.020 -25.110 ;
        RECT 1975.020 -25.120 1978.020 -25.110 ;
        RECT 2065.020 -25.120 2068.020 -25.110 ;
        RECT 2155.020 -25.120 2158.020 -25.110 ;
        RECT 2245.020 -25.120 2248.020 -25.110 ;
        RECT 2335.020 -25.120 2338.020 -25.110 ;
        RECT 2425.020 -25.120 2428.020 -25.110 ;
        RECT 2515.020 -25.120 2518.020 -25.110 ;
        RECT 2605.020 -25.120 2608.020 -25.110 ;
        RECT 2695.020 -25.120 2698.020 -25.110 ;
        RECT 2785.020 -25.120 2788.020 -25.110 ;
        RECT 2875.020 -25.120 2878.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 85.020 -28.130 88.020 -28.120 ;
        RECT 175.020 -28.130 178.020 -28.120 ;
        RECT 265.020 -28.130 268.020 -28.120 ;
        RECT 355.020 -28.130 358.020 -28.120 ;
        RECT 445.020 -28.130 448.020 -28.120 ;
        RECT 535.020 -28.130 538.020 -28.120 ;
        RECT 625.020 -28.130 628.020 -28.120 ;
        RECT 715.020 -28.130 718.020 -28.120 ;
        RECT 805.020 -28.130 808.020 -28.120 ;
        RECT 895.020 -28.130 898.020 -28.120 ;
        RECT 985.020 -28.130 988.020 -28.120 ;
        RECT 1075.020 -28.130 1078.020 -28.120 ;
        RECT 1165.020 -28.130 1168.020 -28.120 ;
        RECT 1255.020 -28.130 1258.020 -28.120 ;
        RECT 1345.020 -28.130 1348.020 -28.120 ;
        RECT 1435.020 -28.130 1438.020 -28.120 ;
        RECT 1525.020 -28.130 1528.020 -28.120 ;
        RECT 1615.020 -28.130 1618.020 -28.120 ;
        RECT 1705.020 -28.130 1708.020 -28.120 ;
        RECT 1795.020 -28.130 1798.020 -28.120 ;
        RECT 1885.020 -28.130 1888.020 -28.120 ;
        RECT 1975.020 -28.130 1978.020 -28.120 ;
        RECT 2065.020 -28.130 2068.020 -28.120 ;
        RECT 2155.020 -28.130 2158.020 -28.120 ;
        RECT 2245.020 -28.130 2248.020 -28.120 ;
        RECT 2335.020 -28.130 2338.020 -28.120 ;
        RECT 2425.020 -28.130 2428.020 -28.120 ;
        RECT 2515.020 -28.130 2518.020 -28.120 ;
        RECT 2605.020 -28.130 2608.020 -28.120 ;
        RECT 2695.020 -28.130 2698.020 -28.120 ;
        RECT 2785.020 -28.130 2788.020 -28.120 ;
        RECT 2875.020 -28.130 2878.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 3519.700 61.020 3557.200 ;
        RECT 148.020 3519.700 151.020 3557.200 ;
        RECT 238.020 3519.700 241.020 3557.200 ;
        RECT 328.020 3519.700 331.020 3557.200 ;
        RECT 418.020 3519.700 421.020 3557.200 ;
        RECT 508.020 3519.700 511.020 3557.200 ;
        RECT 598.020 3519.700 601.020 3557.200 ;
        RECT 688.020 3519.700 691.020 3557.200 ;
        RECT 778.020 3519.700 781.020 3557.200 ;
        RECT 868.020 3519.700 871.020 3557.200 ;
        RECT 958.020 3519.700 961.020 3557.200 ;
        RECT 1048.020 3519.700 1051.020 3557.200 ;
        RECT 1138.020 3519.700 1141.020 3557.200 ;
        RECT 1228.020 3519.700 1231.020 3557.200 ;
        RECT 1318.020 3519.700 1321.020 3557.200 ;
        RECT 1408.020 3519.700 1411.020 3557.200 ;
        RECT 1498.020 3519.700 1501.020 3557.200 ;
        RECT 1588.020 3519.700 1591.020 3557.200 ;
        RECT 1678.020 3519.700 1681.020 3557.200 ;
        RECT 1768.020 3519.700 1771.020 3557.200 ;
        RECT 1858.020 3519.700 1861.020 3557.200 ;
        RECT 1948.020 3519.700 1951.020 3557.200 ;
        RECT 2038.020 3519.700 2041.020 3557.200 ;
        RECT 2128.020 3519.700 2131.020 3557.200 ;
        RECT 2218.020 3519.700 2221.020 3557.200 ;
        RECT 2308.020 3519.700 2311.020 3557.200 ;
        RECT 2398.020 3519.700 2401.020 3557.200 ;
        RECT 2488.020 3519.700 2491.020 3557.200 ;
        RECT 2578.020 3519.700 2581.020 3557.200 ;
        RECT 2668.020 3519.700 2671.020 3557.200 ;
        RECT 2758.020 3519.700 2761.020 3557.200 ;
        RECT 2848.020 3519.700 2851.020 3557.200 ;
        RECT 58.020 -37.520 61.020 0.300 ;
        RECT 148.020 -37.520 151.020 0.300 ;
        RECT 238.020 -37.520 241.020 0.300 ;
        RECT 328.020 -37.520 331.020 0.300 ;
        RECT 418.020 -37.520 421.020 0.300 ;
        RECT 508.020 -37.520 511.020 0.300 ;
        RECT 598.020 -37.520 601.020 0.300 ;
        RECT 688.020 -37.520 691.020 0.300 ;
        RECT 778.020 -37.520 781.020 0.300 ;
        RECT 868.020 -37.520 871.020 0.300 ;
        RECT 958.020 -37.520 961.020 0.300 ;
        RECT 1048.020 -37.520 1051.020 0.300 ;
        RECT 1138.020 -37.520 1141.020 0.300 ;
        RECT 1228.020 -37.520 1231.020 0.300 ;
        RECT 1318.020 -37.520 1321.020 0.300 ;
        RECT 1408.020 -37.520 1411.020 0.300 ;
        RECT 1498.020 -37.520 1501.020 0.300 ;
        RECT 1588.020 -37.520 1591.020 0.300 ;
        RECT 1678.020 -37.520 1681.020 0.300 ;
        RECT 1768.020 -37.520 1771.020 0.300 ;
        RECT 1858.020 -37.520 1861.020 0.300 ;
        RECT 1948.020 -37.520 1951.020 0.300 ;
        RECT 2038.020 -37.520 2041.020 0.300 ;
        RECT 2128.020 -37.520 2131.020 0.300 ;
        RECT 2218.020 -37.520 2221.020 0.300 ;
        RECT 2308.020 -37.520 2311.020 0.300 ;
        RECT 2398.020 -37.520 2401.020 0.300 ;
        RECT 2488.020 -37.520 2491.020 0.300 ;
        RECT 2578.020 -37.520 2581.020 0.300 ;
        RECT 2668.020 -37.520 2671.020 0.300 ;
        RECT 2758.020 -37.520 2761.020 0.300 ;
        RECT 2848.020 -37.520 2851.020 0.300 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 148.930 3551.210 150.110 3552.390 ;
        RECT 148.930 3549.610 150.110 3550.790 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 328.930 3551.210 330.110 3552.390 ;
        RECT 328.930 3549.610 330.110 3550.790 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 508.930 3551.210 510.110 3552.390 ;
        RECT 508.930 3549.610 510.110 3550.790 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 688.930 3551.210 690.110 3552.390 ;
        RECT 688.930 3549.610 690.110 3550.790 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 868.930 3551.210 870.110 3552.390 ;
        RECT 868.930 3549.610 870.110 3550.790 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 1048.930 3551.210 1050.110 3552.390 ;
        RECT 1048.930 3549.610 1050.110 3550.790 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1228.930 3551.210 1230.110 3552.390 ;
        RECT 1228.930 3549.610 1230.110 3550.790 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1408.930 3551.210 1410.110 3552.390 ;
        RECT 1408.930 3549.610 1410.110 3550.790 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1588.930 3551.210 1590.110 3552.390 ;
        RECT 1588.930 3549.610 1590.110 3550.790 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1768.930 3551.210 1770.110 3552.390 ;
        RECT 1768.930 3549.610 1770.110 3550.790 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1948.930 3551.210 1950.110 3552.390 ;
        RECT 1948.930 3549.610 1950.110 3550.790 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2128.930 3551.210 2130.110 3552.390 ;
        RECT 2128.930 3549.610 2130.110 3550.790 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2308.930 3551.210 2310.110 3552.390 ;
        RECT 2308.930 3549.610 2310.110 3550.790 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2488.930 3551.210 2490.110 3552.390 ;
        RECT 2488.930 3549.610 2490.110 3550.790 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2668.930 3551.210 2670.110 3552.390 ;
        RECT 2668.930 3549.610 2670.110 3550.790 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2848.930 3551.210 2850.110 3552.390 ;
        RECT 2848.930 3549.610 2850.110 3550.790 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3395.090 -36.090 3396.270 ;
        RECT -37.270 3393.490 -36.090 3394.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3215.090 -36.090 3216.270 ;
        RECT -37.270 3213.490 -36.090 3214.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 3035.090 -36.090 3036.270 ;
        RECT -37.270 3033.490 -36.090 3034.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2855.090 -36.090 2856.270 ;
        RECT -37.270 2853.490 -36.090 2854.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2675.090 -36.090 2676.270 ;
        RECT -37.270 2673.490 -36.090 2674.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2495.090 -36.090 2496.270 ;
        RECT -37.270 2493.490 -36.090 2494.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2315.090 -36.090 2316.270 ;
        RECT -37.270 2313.490 -36.090 2314.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2135.090 -36.090 2136.270 ;
        RECT -37.270 2133.490 -36.090 2134.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1955.090 -36.090 1956.270 ;
        RECT -37.270 1953.490 -36.090 1954.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1775.090 -36.090 1776.270 ;
        RECT -37.270 1773.490 -36.090 1774.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1595.090 -36.090 1596.270 ;
        RECT -37.270 1593.490 -36.090 1594.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1415.090 -36.090 1416.270 ;
        RECT -37.270 1413.490 -36.090 1414.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1235.090 -36.090 1236.270 ;
        RECT -37.270 1233.490 -36.090 1234.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 1055.090 -36.090 1056.270 ;
        RECT -37.270 1053.490 -36.090 1054.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 875.090 -36.090 876.270 ;
        RECT -37.270 873.490 -36.090 874.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 695.090 -36.090 696.270 ;
        RECT -37.270 693.490 -36.090 694.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 515.090 -36.090 516.270 ;
        RECT -37.270 513.490 -36.090 514.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 335.090 -36.090 336.270 ;
        RECT -37.270 333.490 -36.090 334.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 155.090 -36.090 156.270 ;
        RECT -37.270 153.490 -36.090 154.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3395.090 2956.890 3396.270 ;
        RECT 2955.710 3393.490 2956.890 3394.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3215.090 2956.890 3216.270 ;
        RECT 2955.710 3213.490 2956.890 3214.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 3035.090 2956.890 3036.270 ;
        RECT 2955.710 3033.490 2956.890 3034.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2855.090 2956.890 2856.270 ;
        RECT 2955.710 2853.490 2956.890 2854.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2675.090 2956.890 2676.270 ;
        RECT 2955.710 2673.490 2956.890 2674.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2495.090 2956.890 2496.270 ;
        RECT 2955.710 2493.490 2956.890 2494.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2315.090 2956.890 2316.270 ;
        RECT 2955.710 2313.490 2956.890 2314.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2135.090 2956.890 2136.270 ;
        RECT 2955.710 2133.490 2956.890 2134.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1955.090 2956.890 1956.270 ;
        RECT 2955.710 1953.490 2956.890 1954.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1775.090 2956.890 1776.270 ;
        RECT 2955.710 1773.490 2956.890 1774.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1595.090 2956.890 1596.270 ;
        RECT 2955.710 1593.490 2956.890 1594.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1415.090 2956.890 1416.270 ;
        RECT 2955.710 1413.490 2956.890 1414.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1235.090 2956.890 1236.270 ;
        RECT 2955.710 1233.490 2956.890 1234.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 1055.090 2956.890 1056.270 ;
        RECT 2955.710 1053.490 2956.890 1054.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 875.090 2956.890 876.270 ;
        RECT 2955.710 873.490 2956.890 874.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 695.090 2956.890 696.270 ;
        RECT 2955.710 693.490 2956.890 694.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 515.090 2956.890 516.270 ;
        RECT 2955.710 513.490 2956.890 514.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 335.090 2956.890 336.270 ;
        RECT 2955.710 333.490 2956.890 334.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 155.090 2956.890 156.270 ;
        RECT 2955.710 153.490 2956.890 154.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 148.930 -31.110 150.110 -29.930 ;
        RECT 148.930 -32.710 150.110 -31.530 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 328.930 -31.110 330.110 -29.930 ;
        RECT 328.930 -32.710 330.110 -31.530 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 508.930 -31.110 510.110 -29.930 ;
        RECT 508.930 -32.710 510.110 -31.530 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 688.930 -31.110 690.110 -29.930 ;
        RECT 688.930 -32.710 690.110 -31.530 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 868.930 -31.110 870.110 -29.930 ;
        RECT 868.930 -32.710 870.110 -31.530 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1048.930 -31.110 1050.110 -29.930 ;
        RECT 1048.930 -32.710 1050.110 -31.530 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1228.930 -31.110 1230.110 -29.930 ;
        RECT 1228.930 -32.710 1230.110 -31.530 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1408.930 -31.110 1410.110 -29.930 ;
        RECT 1408.930 -32.710 1410.110 -31.530 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1588.930 -31.110 1590.110 -29.930 ;
        RECT 1588.930 -32.710 1590.110 -31.530 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1768.930 -31.110 1770.110 -29.930 ;
        RECT 1768.930 -32.710 1770.110 -31.530 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 1948.930 -31.110 1950.110 -29.930 ;
        RECT 1948.930 -32.710 1950.110 -31.530 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2128.930 -31.110 2130.110 -29.930 ;
        RECT 2128.930 -32.710 2130.110 -31.530 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2308.930 -31.110 2310.110 -29.930 ;
        RECT 2308.930 -32.710 2310.110 -31.530 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2488.930 -31.110 2490.110 -29.930 ;
        RECT 2488.930 -32.710 2490.110 -31.530 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2668.930 -31.110 2670.110 -29.930 ;
        RECT 2668.930 -32.710 2670.110 -31.530 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2848.930 -31.110 2850.110 -29.930 ;
        RECT 2848.930 -32.710 2850.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 148.020 3552.500 151.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 328.020 3552.500 331.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 508.020 3552.500 511.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 688.020 3552.500 691.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 868.020 3552.500 871.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1048.020 3552.500 1051.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1228.020 3552.500 1231.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1408.020 3552.500 1411.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1588.020 3552.500 1591.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1768.020 3552.500 1771.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 1948.020 3552.500 1951.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2128.020 3552.500 2131.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2308.020 3552.500 2311.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2488.020 3552.500 2491.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2668.020 3552.500 2671.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2848.020 3552.500 2851.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 148.020 3549.490 151.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 328.020 3549.490 331.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 508.020 3549.490 511.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 688.020 3549.490 691.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 868.020 3549.490 871.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1048.020 3549.490 1051.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1228.020 3549.490 1231.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1408.020 3549.490 1411.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1588.020 3549.490 1591.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1768.020 3549.490 1771.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 1948.020 3549.490 1951.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2128.020 3549.490 2131.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2308.020 3549.490 2311.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2488.020 3549.490 2491.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2668.020 3549.490 2671.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2848.020 3549.490 2851.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 0.300 3486.380 ;
        RECT 2919.700 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3396.380 -35.180 3396.390 ;
        RECT 2954.800 3396.380 2957.800 3396.390 ;
        RECT -42.880 3393.380 0.300 3396.380 ;
        RECT 2919.700 3393.380 2962.500 3396.380 ;
        RECT -38.180 3393.370 -35.180 3393.380 ;
        RECT 2954.800 3393.370 2957.800 3393.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 0.300 3306.380 ;
        RECT 2919.700 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3216.380 -35.180 3216.390 ;
        RECT 2954.800 3216.380 2957.800 3216.390 ;
        RECT -42.880 3213.380 0.300 3216.380 ;
        RECT 2919.700 3213.380 2962.500 3216.380 ;
        RECT -38.180 3213.370 -35.180 3213.380 ;
        RECT 2954.800 3213.370 2957.800 3213.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 0.300 3126.380 ;
        RECT 2919.700 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 3036.380 -35.180 3036.390 ;
        RECT 2954.800 3036.380 2957.800 3036.390 ;
        RECT -42.880 3033.380 0.300 3036.380 ;
        RECT 2919.700 3033.380 2962.500 3036.380 ;
        RECT -38.180 3033.370 -35.180 3033.380 ;
        RECT 2954.800 3033.370 2957.800 3033.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 0.300 2946.380 ;
        RECT 2919.700 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2856.380 -35.180 2856.390 ;
        RECT 2954.800 2856.380 2957.800 2856.390 ;
        RECT -42.880 2853.380 0.300 2856.380 ;
        RECT 2919.700 2853.380 2962.500 2856.380 ;
        RECT -38.180 2853.370 -35.180 2853.380 ;
        RECT 2954.800 2853.370 2957.800 2853.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 0.300 2766.380 ;
        RECT 2919.700 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2676.380 -35.180 2676.390 ;
        RECT 2954.800 2676.380 2957.800 2676.390 ;
        RECT -42.880 2673.380 0.300 2676.380 ;
        RECT 2919.700 2673.380 2962.500 2676.380 ;
        RECT -38.180 2673.370 -35.180 2673.380 ;
        RECT 2954.800 2673.370 2957.800 2673.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 0.300 2586.380 ;
        RECT 2919.700 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2496.380 -35.180 2496.390 ;
        RECT 2954.800 2496.380 2957.800 2496.390 ;
        RECT -42.880 2493.380 0.300 2496.380 ;
        RECT 2919.700 2493.380 2962.500 2496.380 ;
        RECT -38.180 2493.370 -35.180 2493.380 ;
        RECT 2954.800 2493.370 2957.800 2493.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 0.300 2406.380 ;
        RECT 2919.700 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2316.380 -35.180 2316.390 ;
        RECT 2954.800 2316.380 2957.800 2316.390 ;
        RECT -42.880 2313.380 0.300 2316.380 ;
        RECT 2919.700 2313.380 2962.500 2316.380 ;
        RECT -38.180 2313.370 -35.180 2313.380 ;
        RECT 2954.800 2313.370 2957.800 2313.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 0.300 2226.380 ;
        RECT 2919.700 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2136.380 -35.180 2136.390 ;
        RECT 2954.800 2136.380 2957.800 2136.390 ;
        RECT -42.880 2133.380 0.300 2136.380 ;
        RECT 2919.700 2133.380 2962.500 2136.380 ;
        RECT -38.180 2133.370 -35.180 2133.380 ;
        RECT 2954.800 2133.370 2957.800 2133.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 0.300 2046.380 ;
        RECT 2919.700 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1956.380 -35.180 1956.390 ;
        RECT 2954.800 1956.380 2957.800 1956.390 ;
        RECT -42.880 1953.380 0.300 1956.380 ;
        RECT 2919.700 1953.380 2962.500 1956.380 ;
        RECT -38.180 1953.370 -35.180 1953.380 ;
        RECT 2954.800 1953.370 2957.800 1953.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 0.300 1866.380 ;
        RECT 2919.700 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1776.380 -35.180 1776.390 ;
        RECT 2954.800 1776.380 2957.800 1776.390 ;
        RECT -42.880 1773.380 0.300 1776.380 ;
        RECT 2919.700 1773.380 2962.500 1776.380 ;
        RECT -38.180 1773.370 -35.180 1773.380 ;
        RECT 2954.800 1773.370 2957.800 1773.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 0.300 1686.380 ;
        RECT 2919.700 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1596.380 -35.180 1596.390 ;
        RECT 2954.800 1596.380 2957.800 1596.390 ;
        RECT -42.880 1593.380 0.300 1596.380 ;
        RECT 2919.700 1593.380 2962.500 1596.380 ;
        RECT -38.180 1593.370 -35.180 1593.380 ;
        RECT 2954.800 1593.370 2957.800 1593.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 0.300 1506.380 ;
        RECT 2919.700 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1416.380 -35.180 1416.390 ;
        RECT 2954.800 1416.380 2957.800 1416.390 ;
        RECT -42.880 1413.380 0.300 1416.380 ;
        RECT 2919.700 1413.380 2962.500 1416.380 ;
        RECT -38.180 1413.370 -35.180 1413.380 ;
        RECT 2954.800 1413.370 2957.800 1413.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 0.300 1326.380 ;
        RECT 2919.700 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1236.380 -35.180 1236.390 ;
        RECT 2954.800 1236.380 2957.800 1236.390 ;
        RECT -42.880 1233.380 0.300 1236.380 ;
        RECT 2919.700 1233.380 2962.500 1236.380 ;
        RECT -38.180 1233.370 -35.180 1233.380 ;
        RECT 2954.800 1233.370 2957.800 1233.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 0.300 1146.380 ;
        RECT 2919.700 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 1056.380 -35.180 1056.390 ;
        RECT 2954.800 1056.380 2957.800 1056.390 ;
        RECT -42.880 1053.380 0.300 1056.380 ;
        RECT 2919.700 1053.380 2962.500 1056.380 ;
        RECT -38.180 1053.370 -35.180 1053.380 ;
        RECT 2954.800 1053.370 2957.800 1053.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 0.300 966.380 ;
        RECT 2919.700 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 876.380 -35.180 876.390 ;
        RECT 2954.800 876.380 2957.800 876.390 ;
        RECT -42.880 873.380 0.300 876.380 ;
        RECT 2919.700 873.380 2962.500 876.380 ;
        RECT -38.180 873.370 -35.180 873.380 ;
        RECT 2954.800 873.370 2957.800 873.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 0.300 786.380 ;
        RECT 2919.700 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 696.380 -35.180 696.390 ;
        RECT 2954.800 696.380 2957.800 696.390 ;
        RECT -42.880 693.380 0.300 696.380 ;
        RECT 2919.700 693.380 2962.500 696.380 ;
        RECT -38.180 693.370 -35.180 693.380 ;
        RECT 2954.800 693.370 2957.800 693.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 0.300 606.380 ;
        RECT 2919.700 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 516.380 -35.180 516.390 ;
        RECT 2954.800 516.380 2957.800 516.390 ;
        RECT -42.880 513.380 0.300 516.380 ;
        RECT 2919.700 513.380 2962.500 516.380 ;
        RECT -38.180 513.370 -35.180 513.380 ;
        RECT 2954.800 513.370 2957.800 513.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 0.300 426.380 ;
        RECT 2919.700 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 336.380 -35.180 336.390 ;
        RECT 2954.800 336.380 2957.800 336.390 ;
        RECT -42.880 333.380 0.300 336.380 ;
        RECT 2919.700 333.380 2962.500 336.380 ;
        RECT -38.180 333.370 -35.180 333.380 ;
        RECT 2954.800 333.370 2957.800 333.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 0.300 246.380 ;
        RECT 2919.700 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 156.380 -35.180 156.390 ;
        RECT 2954.800 156.380 2957.800 156.390 ;
        RECT -42.880 153.380 0.300 156.380 ;
        RECT 2919.700 153.380 2962.500 156.380 ;
        RECT -38.180 153.370 -35.180 153.380 ;
        RECT 2954.800 153.370 2957.800 153.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 0.300 66.380 ;
        RECT 2919.700 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 148.020 -29.820 151.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 328.020 -29.820 331.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 508.020 -29.820 511.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 688.020 -29.820 691.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 868.020 -29.820 871.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1048.020 -29.820 1051.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1228.020 -29.820 1231.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1408.020 -29.820 1411.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1588.020 -29.820 1591.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1768.020 -29.820 1771.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 1948.020 -29.820 1951.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2128.020 -29.820 2131.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2308.020 -29.820 2311.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2488.020 -29.820 2491.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2668.020 -29.820 2671.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2848.020 -29.820 2851.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 148.020 -32.830 151.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 328.020 -32.830 331.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 508.020 -32.830 511.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 688.020 -32.830 691.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 868.020 -32.830 871.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1048.020 -32.830 1051.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1228.020 -32.830 1231.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1408.020 -32.830 1411.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1588.020 -32.830 1591.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1768.020 -32.830 1771.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 1948.020 -32.830 1951.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2128.020 -32.830 2131.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2308.020 -32.830 2311.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2488.020 -32.830 2491.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2668.020 -32.830 2671.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2848.020 -32.830 2851.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 103.020 3519.700 106.020 3557.200 ;
        RECT 193.020 3519.700 196.020 3557.200 ;
        RECT 283.020 3519.700 286.020 3557.200 ;
        RECT 373.020 3519.700 376.020 3557.200 ;
        RECT 463.020 3519.700 466.020 3557.200 ;
        RECT 553.020 3519.700 556.020 3557.200 ;
        RECT 643.020 3519.700 646.020 3557.200 ;
        RECT 733.020 3519.700 736.020 3557.200 ;
        RECT 823.020 3519.700 826.020 3557.200 ;
        RECT 913.020 3519.700 916.020 3557.200 ;
        RECT 1003.020 3519.700 1006.020 3557.200 ;
        RECT 1093.020 3519.700 1096.020 3557.200 ;
        RECT 1183.020 3519.700 1186.020 3557.200 ;
        RECT 1273.020 3519.700 1276.020 3557.200 ;
        RECT 1363.020 3519.700 1366.020 3557.200 ;
        RECT 1453.020 3519.700 1456.020 3557.200 ;
        RECT 1543.020 3519.700 1546.020 3557.200 ;
        RECT 1633.020 3519.700 1636.020 3557.200 ;
        RECT 1723.020 3519.700 1726.020 3557.200 ;
        RECT 1813.020 3519.700 1816.020 3557.200 ;
        RECT 1903.020 3519.700 1906.020 3557.200 ;
        RECT 1993.020 3519.700 1996.020 3557.200 ;
        RECT 2083.020 3519.700 2086.020 3557.200 ;
        RECT 2173.020 3519.700 2176.020 3557.200 ;
        RECT 2263.020 3519.700 2266.020 3557.200 ;
        RECT 2353.020 3519.700 2356.020 3557.200 ;
        RECT 2443.020 3519.700 2446.020 3557.200 ;
        RECT 2533.020 3519.700 2536.020 3557.200 ;
        RECT 2623.020 3519.700 2626.020 3557.200 ;
        RECT 2713.020 3519.700 2716.020 3557.200 ;
        RECT 2803.020 3519.700 2806.020 3557.200 ;
        RECT 2893.020 3519.700 2896.020 3557.200 ;
        RECT 103.020 -37.520 106.020 0.300 ;
        RECT 193.020 -37.520 196.020 0.300 ;
        RECT 283.020 -37.520 286.020 0.300 ;
        RECT 373.020 -37.520 376.020 0.300 ;
        RECT 463.020 -37.520 466.020 0.300 ;
        RECT 553.020 -37.520 556.020 0.300 ;
        RECT 643.020 -37.520 646.020 0.300 ;
        RECT 733.020 -37.520 736.020 0.300 ;
        RECT 823.020 -37.520 826.020 0.300 ;
        RECT 913.020 -37.520 916.020 0.300 ;
        RECT 1003.020 -37.520 1006.020 0.300 ;
        RECT 1093.020 -37.520 1096.020 0.300 ;
        RECT 1183.020 -37.520 1186.020 0.300 ;
        RECT 1273.020 -37.520 1276.020 0.300 ;
        RECT 1363.020 -37.520 1366.020 0.300 ;
        RECT 1453.020 -37.520 1456.020 0.300 ;
        RECT 1543.020 -37.520 1546.020 0.300 ;
        RECT 1633.020 -37.520 1636.020 0.300 ;
        RECT 1723.020 -37.520 1726.020 0.300 ;
        RECT 1813.020 -37.520 1816.020 0.300 ;
        RECT 1903.020 -37.520 1906.020 0.300 ;
        RECT 1993.020 -37.520 1996.020 0.300 ;
        RECT 2083.020 -37.520 2086.020 0.300 ;
        RECT 2173.020 -37.520 2176.020 0.300 ;
        RECT 2263.020 -37.520 2266.020 0.300 ;
        RECT 2353.020 -37.520 2356.020 0.300 ;
        RECT 2443.020 -37.520 2446.020 0.300 ;
        RECT 2533.020 -37.520 2536.020 0.300 ;
        RECT 2623.020 -37.520 2626.020 0.300 ;
        RECT 2713.020 -37.520 2716.020 0.300 ;
        RECT 2803.020 -37.520 2806.020 0.300 ;
        RECT 2893.020 -37.520 2896.020 0.300 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 103.930 3555.910 105.110 3557.090 ;
        RECT 103.930 3554.310 105.110 3555.490 ;
        RECT 193.930 3555.910 195.110 3557.090 ;
        RECT 193.930 3554.310 195.110 3555.490 ;
        RECT 283.930 3555.910 285.110 3557.090 ;
        RECT 283.930 3554.310 285.110 3555.490 ;
        RECT 373.930 3555.910 375.110 3557.090 ;
        RECT 373.930 3554.310 375.110 3555.490 ;
        RECT 463.930 3555.910 465.110 3557.090 ;
        RECT 463.930 3554.310 465.110 3555.490 ;
        RECT 553.930 3555.910 555.110 3557.090 ;
        RECT 553.930 3554.310 555.110 3555.490 ;
        RECT 643.930 3555.910 645.110 3557.090 ;
        RECT 643.930 3554.310 645.110 3555.490 ;
        RECT 733.930 3555.910 735.110 3557.090 ;
        RECT 733.930 3554.310 735.110 3555.490 ;
        RECT 823.930 3555.910 825.110 3557.090 ;
        RECT 823.930 3554.310 825.110 3555.490 ;
        RECT 913.930 3555.910 915.110 3557.090 ;
        RECT 913.930 3554.310 915.110 3555.490 ;
        RECT 1003.930 3555.910 1005.110 3557.090 ;
        RECT 1003.930 3554.310 1005.110 3555.490 ;
        RECT 1093.930 3555.910 1095.110 3557.090 ;
        RECT 1093.930 3554.310 1095.110 3555.490 ;
        RECT 1183.930 3555.910 1185.110 3557.090 ;
        RECT 1183.930 3554.310 1185.110 3555.490 ;
        RECT 1273.930 3555.910 1275.110 3557.090 ;
        RECT 1273.930 3554.310 1275.110 3555.490 ;
        RECT 1363.930 3555.910 1365.110 3557.090 ;
        RECT 1363.930 3554.310 1365.110 3555.490 ;
        RECT 1453.930 3555.910 1455.110 3557.090 ;
        RECT 1453.930 3554.310 1455.110 3555.490 ;
        RECT 1543.930 3555.910 1545.110 3557.090 ;
        RECT 1543.930 3554.310 1545.110 3555.490 ;
        RECT 1633.930 3555.910 1635.110 3557.090 ;
        RECT 1633.930 3554.310 1635.110 3555.490 ;
        RECT 1723.930 3555.910 1725.110 3557.090 ;
        RECT 1723.930 3554.310 1725.110 3555.490 ;
        RECT 1813.930 3555.910 1815.110 3557.090 ;
        RECT 1813.930 3554.310 1815.110 3555.490 ;
        RECT 1903.930 3555.910 1905.110 3557.090 ;
        RECT 1903.930 3554.310 1905.110 3555.490 ;
        RECT 1993.930 3555.910 1995.110 3557.090 ;
        RECT 1993.930 3554.310 1995.110 3555.490 ;
        RECT 2083.930 3555.910 2085.110 3557.090 ;
        RECT 2083.930 3554.310 2085.110 3555.490 ;
        RECT 2173.930 3555.910 2175.110 3557.090 ;
        RECT 2173.930 3554.310 2175.110 3555.490 ;
        RECT 2263.930 3555.910 2265.110 3557.090 ;
        RECT 2263.930 3554.310 2265.110 3555.490 ;
        RECT 2353.930 3555.910 2355.110 3557.090 ;
        RECT 2353.930 3554.310 2355.110 3555.490 ;
        RECT 2443.930 3555.910 2445.110 3557.090 ;
        RECT 2443.930 3554.310 2445.110 3555.490 ;
        RECT 2533.930 3555.910 2535.110 3557.090 ;
        RECT 2533.930 3554.310 2535.110 3555.490 ;
        RECT 2623.930 3555.910 2625.110 3557.090 ;
        RECT 2623.930 3554.310 2625.110 3555.490 ;
        RECT 2713.930 3555.910 2715.110 3557.090 ;
        RECT 2713.930 3554.310 2715.110 3555.490 ;
        RECT 2803.930 3555.910 2805.110 3557.090 ;
        RECT 2803.930 3554.310 2805.110 3555.490 ;
        RECT 2893.930 3555.910 2895.110 3557.090 ;
        RECT 2893.930 3554.310 2895.110 3555.490 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT -41.970 3440.090 -40.790 3441.270 ;
        RECT -41.970 3438.490 -40.790 3439.670 ;
        RECT -41.970 3350.090 -40.790 3351.270 ;
        RECT -41.970 3348.490 -40.790 3349.670 ;
        RECT -41.970 3260.090 -40.790 3261.270 ;
        RECT -41.970 3258.490 -40.790 3259.670 ;
        RECT -41.970 3170.090 -40.790 3171.270 ;
        RECT -41.970 3168.490 -40.790 3169.670 ;
        RECT -41.970 3080.090 -40.790 3081.270 ;
        RECT -41.970 3078.490 -40.790 3079.670 ;
        RECT -41.970 2990.090 -40.790 2991.270 ;
        RECT -41.970 2988.490 -40.790 2989.670 ;
        RECT -41.970 2900.090 -40.790 2901.270 ;
        RECT -41.970 2898.490 -40.790 2899.670 ;
        RECT -41.970 2810.090 -40.790 2811.270 ;
        RECT -41.970 2808.490 -40.790 2809.670 ;
        RECT -41.970 2720.090 -40.790 2721.270 ;
        RECT -41.970 2718.490 -40.790 2719.670 ;
        RECT -41.970 2630.090 -40.790 2631.270 ;
        RECT -41.970 2628.490 -40.790 2629.670 ;
        RECT -41.970 2540.090 -40.790 2541.270 ;
        RECT -41.970 2538.490 -40.790 2539.670 ;
        RECT -41.970 2450.090 -40.790 2451.270 ;
        RECT -41.970 2448.490 -40.790 2449.670 ;
        RECT -41.970 2360.090 -40.790 2361.270 ;
        RECT -41.970 2358.490 -40.790 2359.670 ;
        RECT -41.970 2270.090 -40.790 2271.270 ;
        RECT -41.970 2268.490 -40.790 2269.670 ;
        RECT -41.970 2180.090 -40.790 2181.270 ;
        RECT -41.970 2178.490 -40.790 2179.670 ;
        RECT -41.970 2090.090 -40.790 2091.270 ;
        RECT -41.970 2088.490 -40.790 2089.670 ;
        RECT -41.970 2000.090 -40.790 2001.270 ;
        RECT -41.970 1998.490 -40.790 1999.670 ;
        RECT -41.970 1910.090 -40.790 1911.270 ;
        RECT -41.970 1908.490 -40.790 1909.670 ;
        RECT -41.970 1820.090 -40.790 1821.270 ;
        RECT -41.970 1818.490 -40.790 1819.670 ;
        RECT -41.970 1730.090 -40.790 1731.270 ;
        RECT -41.970 1728.490 -40.790 1729.670 ;
        RECT -41.970 1640.090 -40.790 1641.270 ;
        RECT -41.970 1638.490 -40.790 1639.670 ;
        RECT -41.970 1550.090 -40.790 1551.270 ;
        RECT -41.970 1548.490 -40.790 1549.670 ;
        RECT -41.970 1460.090 -40.790 1461.270 ;
        RECT -41.970 1458.490 -40.790 1459.670 ;
        RECT -41.970 1370.090 -40.790 1371.270 ;
        RECT -41.970 1368.490 -40.790 1369.670 ;
        RECT -41.970 1280.090 -40.790 1281.270 ;
        RECT -41.970 1278.490 -40.790 1279.670 ;
        RECT -41.970 1190.090 -40.790 1191.270 ;
        RECT -41.970 1188.490 -40.790 1189.670 ;
        RECT -41.970 1100.090 -40.790 1101.270 ;
        RECT -41.970 1098.490 -40.790 1099.670 ;
        RECT -41.970 1010.090 -40.790 1011.270 ;
        RECT -41.970 1008.490 -40.790 1009.670 ;
        RECT -41.970 920.090 -40.790 921.270 ;
        RECT -41.970 918.490 -40.790 919.670 ;
        RECT -41.970 830.090 -40.790 831.270 ;
        RECT -41.970 828.490 -40.790 829.670 ;
        RECT -41.970 740.090 -40.790 741.270 ;
        RECT -41.970 738.490 -40.790 739.670 ;
        RECT -41.970 650.090 -40.790 651.270 ;
        RECT -41.970 648.490 -40.790 649.670 ;
        RECT -41.970 560.090 -40.790 561.270 ;
        RECT -41.970 558.490 -40.790 559.670 ;
        RECT -41.970 470.090 -40.790 471.270 ;
        RECT -41.970 468.490 -40.790 469.670 ;
        RECT -41.970 380.090 -40.790 381.270 ;
        RECT -41.970 378.490 -40.790 379.670 ;
        RECT -41.970 290.090 -40.790 291.270 ;
        RECT -41.970 288.490 -40.790 289.670 ;
        RECT -41.970 200.090 -40.790 201.270 ;
        RECT -41.970 198.490 -40.790 199.670 ;
        RECT -41.970 110.090 -40.790 111.270 ;
        RECT -41.970 108.490 -40.790 109.670 ;
        RECT 2960.410 3440.090 2961.590 3441.270 ;
        RECT 2960.410 3438.490 2961.590 3439.670 ;
        RECT 2960.410 3350.090 2961.590 3351.270 ;
        RECT 2960.410 3348.490 2961.590 3349.670 ;
        RECT 2960.410 3260.090 2961.590 3261.270 ;
        RECT 2960.410 3258.490 2961.590 3259.670 ;
        RECT 2960.410 3170.090 2961.590 3171.270 ;
        RECT 2960.410 3168.490 2961.590 3169.670 ;
        RECT 2960.410 3080.090 2961.590 3081.270 ;
        RECT 2960.410 3078.490 2961.590 3079.670 ;
        RECT 2960.410 2990.090 2961.590 2991.270 ;
        RECT 2960.410 2988.490 2961.590 2989.670 ;
        RECT 2960.410 2900.090 2961.590 2901.270 ;
        RECT 2960.410 2898.490 2961.590 2899.670 ;
        RECT 2960.410 2810.090 2961.590 2811.270 ;
        RECT 2960.410 2808.490 2961.590 2809.670 ;
        RECT 2960.410 2720.090 2961.590 2721.270 ;
        RECT 2960.410 2718.490 2961.590 2719.670 ;
        RECT 2960.410 2630.090 2961.590 2631.270 ;
        RECT 2960.410 2628.490 2961.590 2629.670 ;
        RECT 2960.410 2540.090 2961.590 2541.270 ;
        RECT 2960.410 2538.490 2961.590 2539.670 ;
        RECT 2960.410 2450.090 2961.590 2451.270 ;
        RECT 2960.410 2448.490 2961.590 2449.670 ;
        RECT 2960.410 2360.090 2961.590 2361.270 ;
        RECT 2960.410 2358.490 2961.590 2359.670 ;
        RECT 2960.410 2270.090 2961.590 2271.270 ;
        RECT 2960.410 2268.490 2961.590 2269.670 ;
        RECT 2960.410 2180.090 2961.590 2181.270 ;
        RECT 2960.410 2178.490 2961.590 2179.670 ;
        RECT 2960.410 2090.090 2961.590 2091.270 ;
        RECT 2960.410 2088.490 2961.590 2089.670 ;
        RECT 2960.410 2000.090 2961.590 2001.270 ;
        RECT 2960.410 1998.490 2961.590 1999.670 ;
        RECT 2960.410 1910.090 2961.590 1911.270 ;
        RECT 2960.410 1908.490 2961.590 1909.670 ;
        RECT 2960.410 1820.090 2961.590 1821.270 ;
        RECT 2960.410 1818.490 2961.590 1819.670 ;
        RECT 2960.410 1730.090 2961.590 1731.270 ;
        RECT 2960.410 1728.490 2961.590 1729.670 ;
        RECT 2960.410 1640.090 2961.590 1641.270 ;
        RECT 2960.410 1638.490 2961.590 1639.670 ;
        RECT 2960.410 1550.090 2961.590 1551.270 ;
        RECT 2960.410 1548.490 2961.590 1549.670 ;
        RECT 2960.410 1460.090 2961.590 1461.270 ;
        RECT 2960.410 1458.490 2961.590 1459.670 ;
        RECT 2960.410 1370.090 2961.590 1371.270 ;
        RECT 2960.410 1368.490 2961.590 1369.670 ;
        RECT 2960.410 1280.090 2961.590 1281.270 ;
        RECT 2960.410 1278.490 2961.590 1279.670 ;
        RECT 2960.410 1190.090 2961.590 1191.270 ;
        RECT 2960.410 1188.490 2961.590 1189.670 ;
        RECT 2960.410 1100.090 2961.590 1101.270 ;
        RECT 2960.410 1098.490 2961.590 1099.670 ;
        RECT 2960.410 1010.090 2961.590 1011.270 ;
        RECT 2960.410 1008.490 2961.590 1009.670 ;
        RECT 2960.410 920.090 2961.590 921.270 ;
        RECT 2960.410 918.490 2961.590 919.670 ;
        RECT 2960.410 830.090 2961.590 831.270 ;
        RECT 2960.410 828.490 2961.590 829.670 ;
        RECT 2960.410 740.090 2961.590 741.270 ;
        RECT 2960.410 738.490 2961.590 739.670 ;
        RECT 2960.410 650.090 2961.590 651.270 ;
        RECT 2960.410 648.490 2961.590 649.670 ;
        RECT 2960.410 560.090 2961.590 561.270 ;
        RECT 2960.410 558.490 2961.590 559.670 ;
        RECT 2960.410 470.090 2961.590 471.270 ;
        RECT 2960.410 468.490 2961.590 469.670 ;
        RECT 2960.410 380.090 2961.590 381.270 ;
        RECT 2960.410 378.490 2961.590 379.670 ;
        RECT 2960.410 290.090 2961.590 291.270 ;
        RECT 2960.410 288.490 2961.590 289.670 ;
        RECT 2960.410 200.090 2961.590 201.270 ;
        RECT 2960.410 198.490 2961.590 199.670 ;
        RECT 2960.410 110.090 2961.590 111.270 ;
        RECT 2960.410 108.490 2961.590 109.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 103.930 -35.810 105.110 -34.630 ;
        RECT 103.930 -37.410 105.110 -36.230 ;
        RECT 193.930 -35.810 195.110 -34.630 ;
        RECT 193.930 -37.410 195.110 -36.230 ;
        RECT 283.930 -35.810 285.110 -34.630 ;
        RECT 283.930 -37.410 285.110 -36.230 ;
        RECT 373.930 -35.810 375.110 -34.630 ;
        RECT 373.930 -37.410 375.110 -36.230 ;
        RECT 463.930 -35.810 465.110 -34.630 ;
        RECT 463.930 -37.410 465.110 -36.230 ;
        RECT 553.930 -35.810 555.110 -34.630 ;
        RECT 553.930 -37.410 555.110 -36.230 ;
        RECT 643.930 -35.810 645.110 -34.630 ;
        RECT 643.930 -37.410 645.110 -36.230 ;
        RECT 733.930 -35.810 735.110 -34.630 ;
        RECT 733.930 -37.410 735.110 -36.230 ;
        RECT 823.930 -35.810 825.110 -34.630 ;
        RECT 823.930 -37.410 825.110 -36.230 ;
        RECT 913.930 -35.810 915.110 -34.630 ;
        RECT 913.930 -37.410 915.110 -36.230 ;
        RECT 1003.930 -35.810 1005.110 -34.630 ;
        RECT 1003.930 -37.410 1005.110 -36.230 ;
        RECT 1093.930 -35.810 1095.110 -34.630 ;
        RECT 1093.930 -37.410 1095.110 -36.230 ;
        RECT 1183.930 -35.810 1185.110 -34.630 ;
        RECT 1183.930 -37.410 1185.110 -36.230 ;
        RECT 1273.930 -35.810 1275.110 -34.630 ;
        RECT 1273.930 -37.410 1275.110 -36.230 ;
        RECT 1363.930 -35.810 1365.110 -34.630 ;
        RECT 1363.930 -37.410 1365.110 -36.230 ;
        RECT 1453.930 -35.810 1455.110 -34.630 ;
        RECT 1453.930 -37.410 1455.110 -36.230 ;
        RECT 1543.930 -35.810 1545.110 -34.630 ;
        RECT 1543.930 -37.410 1545.110 -36.230 ;
        RECT 1633.930 -35.810 1635.110 -34.630 ;
        RECT 1633.930 -37.410 1635.110 -36.230 ;
        RECT 1723.930 -35.810 1725.110 -34.630 ;
        RECT 1723.930 -37.410 1725.110 -36.230 ;
        RECT 1813.930 -35.810 1815.110 -34.630 ;
        RECT 1813.930 -37.410 1815.110 -36.230 ;
        RECT 1903.930 -35.810 1905.110 -34.630 ;
        RECT 1903.930 -37.410 1905.110 -36.230 ;
        RECT 1993.930 -35.810 1995.110 -34.630 ;
        RECT 1993.930 -37.410 1995.110 -36.230 ;
        RECT 2083.930 -35.810 2085.110 -34.630 ;
        RECT 2083.930 -37.410 2085.110 -36.230 ;
        RECT 2173.930 -35.810 2175.110 -34.630 ;
        RECT 2173.930 -37.410 2175.110 -36.230 ;
        RECT 2263.930 -35.810 2265.110 -34.630 ;
        RECT 2263.930 -37.410 2265.110 -36.230 ;
        RECT 2353.930 -35.810 2355.110 -34.630 ;
        RECT 2353.930 -37.410 2355.110 -36.230 ;
        RECT 2443.930 -35.810 2445.110 -34.630 ;
        RECT 2443.930 -37.410 2445.110 -36.230 ;
        RECT 2533.930 -35.810 2535.110 -34.630 ;
        RECT 2533.930 -37.410 2535.110 -36.230 ;
        RECT 2623.930 -35.810 2625.110 -34.630 ;
        RECT 2623.930 -37.410 2625.110 -36.230 ;
        RECT 2713.930 -35.810 2715.110 -34.630 ;
        RECT 2713.930 -37.410 2715.110 -36.230 ;
        RECT 2803.930 -35.810 2805.110 -34.630 ;
        RECT 2803.930 -37.410 2805.110 -36.230 ;
        RECT 2893.930 -35.810 2895.110 -34.630 ;
        RECT 2893.930 -37.410 2895.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 103.020 3557.200 106.020 3557.210 ;
        RECT 193.020 3557.200 196.020 3557.210 ;
        RECT 283.020 3557.200 286.020 3557.210 ;
        RECT 373.020 3557.200 376.020 3557.210 ;
        RECT 463.020 3557.200 466.020 3557.210 ;
        RECT 553.020 3557.200 556.020 3557.210 ;
        RECT 643.020 3557.200 646.020 3557.210 ;
        RECT 733.020 3557.200 736.020 3557.210 ;
        RECT 823.020 3557.200 826.020 3557.210 ;
        RECT 913.020 3557.200 916.020 3557.210 ;
        RECT 1003.020 3557.200 1006.020 3557.210 ;
        RECT 1093.020 3557.200 1096.020 3557.210 ;
        RECT 1183.020 3557.200 1186.020 3557.210 ;
        RECT 1273.020 3557.200 1276.020 3557.210 ;
        RECT 1363.020 3557.200 1366.020 3557.210 ;
        RECT 1453.020 3557.200 1456.020 3557.210 ;
        RECT 1543.020 3557.200 1546.020 3557.210 ;
        RECT 1633.020 3557.200 1636.020 3557.210 ;
        RECT 1723.020 3557.200 1726.020 3557.210 ;
        RECT 1813.020 3557.200 1816.020 3557.210 ;
        RECT 1903.020 3557.200 1906.020 3557.210 ;
        RECT 1993.020 3557.200 1996.020 3557.210 ;
        RECT 2083.020 3557.200 2086.020 3557.210 ;
        RECT 2173.020 3557.200 2176.020 3557.210 ;
        RECT 2263.020 3557.200 2266.020 3557.210 ;
        RECT 2353.020 3557.200 2356.020 3557.210 ;
        RECT 2443.020 3557.200 2446.020 3557.210 ;
        RECT 2533.020 3557.200 2536.020 3557.210 ;
        RECT 2623.020 3557.200 2626.020 3557.210 ;
        RECT 2713.020 3557.200 2716.020 3557.210 ;
        RECT 2803.020 3557.200 2806.020 3557.210 ;
        RECT 2893.020 3557.200 2896.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 103.020 3554.190 106.020 3554.200 ;
        RECT 193.020 3554.190 196.020 3554.200 ;
        RECT 283.020 3554.190 286.020 3554.200 ;
        RECT 373.020 3554.190 376.020 3554.200 ;
        RECT 463.020 3554.190 466.020 3554.200 ;
        RECT 553.020 3554.190 556.020 3554.200 ;
        RECT 643.020 3554.190 646.020 3554.200 ;
        RECT 733.020 3554.190 736.020 3554.200 ;
        RECT 823.020 3554.190 826.020 3554.200 ;
        RECT 913.020 3554.190 916.020 3554.200 ;
        RECT 1003.020 3554.190 1006.020 3554.200 ;
        RECT 1093.020 3554.190 1096.020 3554.200 ;
        RECT 1183.020 3554.190 1186.020 3554.200 ;
        RECT 1273.020 3554.190 1276.020 3554.200 ;
        RECT 1363.020 3554.190 1366.020 3554.200 ;
        RECT 1453.020 3554.190 1456.020 3554.200 ;
        RECT 1543.020 3554.190 1546.020 3554.200 ;
        RECT 1633.020 3554.190 1636.020 3554.200 ;
        RECT 1723.020 3554.190 1726.020 3554.200 ;
        RECT 1813.020 3554.190 1816.020 3554.200 ;
        RECT 1903.020 3554.190 1906.020 3554.200 ;
        RECT 1993.020 3554.190 1996.020 3554.200 ;
        RECT 2083.020 3554.190 2086.020 3554.200 ;
        RECT 2173.020 3554.190 2176.020 3554.200 ;
        RECT 2263.020 3554.190 2266.020 3554.200 ;
        RECT 2353.020 3554.190 2356.020 3554.200 ;
        RECT 2443.020 3554.190 2446.020 3554.200 ;
        RECT 2533.020 3554.190 2536.020 3554.200 ;
        RECT 2623.020 3554.190 2626.020 3554.200 ;
        RECT 2713.020 3554.190 2716.020 3554.200 ;
        RECT 2803.020 3554.190 2806.020 3554.200 ;
        RECT 2893.020 3554.190 2896.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3441.380 -39.880 3441.390 ;
        RECT 2959.500 3441.380 2962.500 3441.390 ;
        RECT -42.880 3438.380 0.300 3441.380 ;
        RECT 2919.700 3438.380 2962.500 3441.380 ;
        RECT -42.880 3438.370 -39.880 3438.380 ;
        RECT 2959.500 3438.370 2962.500 3438.380 ;
        RECT -42.880 3351.380 -39.880 3351.390 ;
        RECT 2959.500 3351.380 2962.500 3351.390 ;
        RECT -42.880 3348.380 0.300 3351.380 ;
        RECT 2919.700 3348.380 2962.500 3351.380 ;
        RECT -42.880 3348.370 -39.880 3348.380 ;
        RECT 2959.500 3348.370 2962.500 3348.380 ;
        RECT -42.880 3261.380 -39.880 3261.390 ;
        RECT 2959.500 3261.380 2962.500 3261.390 ;
        RECT -42.880 3258.380 0.300 3261.380 ;
        RECT 2919.700 3258.380 2962.500 3261.380 ;
        RECT -42.880 3258.370 -39.880 3258.380 ;
        RECT 2959.500 3258.370 2962.500 3258.380 ;
        RECT -42.880 3171.380 -39.880 3171.390 ;
        RECT 2959.500 3171.380 2962.500 3171.390 ;
        RECT -42.880 3168.380 0.300 3171.380 ;
        RECT 2919.700 3168.380 2962.500 3171.380 ;
        RECT -42.880 3168.370 -39.880 3168.380 ;
        RECT 2959.500 3168.370 2962.500 3168.380 ;
        RECT -42.880 3081.380 -39.880 3081.390 ;
        RECT 2959.500 3081.380 2962.500 3081.390 ;
        RECT -42.880 3078.380 0.300 3081.380 ;
        RECT 2919.700 3078.380 2962.500 3081.380 ;
        RECT -42.880 3078.370 -39.880 3078.380 ;
        RECT 2959.500 3078.370 2962.500 3078.380 ;
        RECT -42.880 2991.380 -39.880 2991.390 ;
        RECT 2959.500 2991.380 2962.500 2991.390 ;
        RECT -42.880 2988.380 0.300 2991.380 ;
        RECT 2919.700 2988.380 2962.500 2991.380 ;
        RECT -42.880 2988.370 -39.880 2988.380 ;
        RECT 2959.500 2988.370 2962.500 2988.380 ;
        RECT -42.880 2901.380 -39.880 2901.390 ;
        RECT 2959.500 2901.380 2962.500 2901.390 ;
        RECT -42.880 2898.380 0.300 2901.380 ;
        RECT 2919.700 2898.380 2962.500 2901.380 ;
        RECT -42.880 2898.370 -39.880 2898.380 ;
        RECT 2959.500 2898.370 2962.500 2898.380 ;
        RECT -42.880 2811.380 -39.880 2811.390 ;
        RECT 2959.500 2811.380 2962.500 2811.390 ;
        RECT -42.880 2808.380 0.300 2811.380 ;
        RECT 2919.700 2808.380 2962.500 2811.380 ;
        RECT -42.880 2808.370 -39.880 2808.380 ;
        RECT 2959.500 2808.370 2962.500 2808.380 ;
        RECT -42.880 2721.380 -39.880 2721.390 ;
        RECT 2959.500 2721.380 2962.500 2721.390 ;
        RECT -42.880 2718.380 0.300 2721.380 ;
        RECT 2919.700 2718.380 2962.500 2721.380 ;
        RECT -42.880 2718.370 -39.880 2718.380 ;
        RECT 2959.500 2718.370 2962.500 2718.380 ;
        RECT -42.880 2631.380 -39.880 2631.390 ;
        RECT 2959.500 2631.380 2962.500 2631.390 ;
        RECT -42.880 2628.380 0.300 2631.380 ;
        RECT 2919.700 2628.380 2962.500 2631.380 ;
        RECT -42.880 2628.370 -39.880 2628.380 ;
        RECT 2959.500 2628.370 2962.500 2628.380 ;
        RECT -42.880 2541.380 -39.880 2541.390 ;
        RECT 2959.500 2541.380 2962.500 2541.390 ;
        RECT -42.880 2538.380 0.300 2541.380 ;
        RECT 2919.700 2538.380 2962.500 2541.380 ;
        RECT -42.880 2538.370 -39.880 2538.380 ;
        RECT 2959.500 2538.370 2962.500 2538.380 ;
        RECT -42.880 2451.380 -39.880 2451.390 ;
        RECT 2959.500 2451.380 2962.500 2451.390 ;
        RECT -42.880 2448.380 0.300 2451.380 ;
        RECT 2919.700 2448.380 2962.500 2451.380 ;
        RECT -42.880 2448.370 -39.880 2448.380 ;
        RECT 2959.500 2448.370 2962.500 2448.380 ;
        RECT -42.880 2361.380 -39.880 2361.390 ;
        RECT 2959.500 2361.380 2962.500 2361.390 ;
        RECT -42.880 2358.380 0.300 2361.380 ;
        RECT 2919.700 2358.380 2962.500 2361.380 ;
        RECT -42.880 2358.370 -39.880 2358.380 ;
        RECT 2959.500 2358.370 2962.500 2358.380 ;
        RECT -42.880 2271.380 -39.880 2271.390 ;
        RECT 2959.500 2271.380 2962.500 2271.390 ;
        RECT -42.880 2268.380 0.300 2271.380 ;
        RECT 2919.700 2268.380 2962.500 2271.380 ;
        RECT -42.880 2268.370 -39.880 2268.380 ;
        RECT 2959.500 2268.370 2962.500 2268.380 ;
        RECT -42.880 2181.380 -39.880 2181.390 ;
        RECT 2959.500 2181.380 2962.500 2181.390 ;
        RECT -42.880 2178.380 0.300 2181.380 ;
        RECT 2919.700 2178.380 2962.500 2181.380 ;
        RECT -42.880 2178.370 -39.880 2178.380 ;
        RECT 2959.500 2178.370 2962.500 2178.380 ;
        RECT -42.880 2091.380 -39.880 2091.390 ;
        RECT 2959.500 2091.380 2962.500 2091.390 ;
        RECT -42.880 2088.380 0.300 2091.380 ;
        RECT 2919.700 2088.380 2962.500 2091.380 ;
        RECT -42.880 2088.370 -39.880 2088.380 ;
        RECT 2959.500 2088.370 2962.500 2088.380 ;
        RECT -42.880 2001.380 -39.880 2001.390 ;
        RECT 2959.500 2001.380 2962.500 2001.390 ;
        RECT -42.880 1998.380 0.300 2001.380 ;
        RECT 2919.700 1998.380 2962.500 2001.380 ;
        RECT -42.880 1998.370 -39.880 1998.380 ;
        RECT 2959.500 1998.370 2962.500 1998.380 ;
        RECT -42.880 1911.380 -39.880 1911.390 ;
        RECT 2959.500 1911.380 2962.500 1911.390 ;
        RECT -42.880 1908.380 0.300 1911.380 ;
        RECT 2919.700 1908.380 2962.500 1911.380 ;
        RECT -42.880 1908.370 -39.880 1908.380 ;
        RECT 2959.500 1908.370 2962.500 1908.380 ;
        RECT -42.880 1821.380 -39.880 1821.390 ;
        RECT 2959.500 1821.380 2962.500 1821.390 ;
        RECT -42.880 1818.380 0.300 1821.380 ;
        RECT 2919.700 1818.380 2962.500 1821.380 ;
        RECT -42.880 1818.370 -39.880 1818.380 ;
        RECT 2959.500 1818.370 2962.500 1818.380 ;
        RECT -42.880 1731.380 -39.880 1731.390 ;
        RECT 2959.500 1731.380 2962.500 1731.390 ;
        RECT -42.880 1728.380 0.300 1731.380 ;
        RECT 2919.700 1728.380 2962.500 1731.380 ;
        RECT -42.880 1728.370 -39.880 1728.380 ;
        RECT 2959.500 1728.370 2962.500 1728.380 ;
        RECT -42.880 1641.380 -39.880 1641.390 ;
        RECT 2959.500 1641.380 2962.500 1641.390 ;
        RECT -42.880 1638.380 0.300 1641.380 ;
        RECT 2919.700 1638.380 2962.500 1641.380 ;
        RECT -42.880 1638.370 -39.880 1638.380 ;
        RECT 2959.500 1638.370 2962.500 1638.380 ;
        RECT -42.880 1551.380 -39.880 1551.390 ;
        RECT 2959.500 1551.380 2962.500 1551.390 ;
        RECT -42.880 1548.380 0.300 1551.380 ;
        RECT 2919.700 1548.380 2962.500 1551.380 ;
        RECT -42.880 1548.370 -39.880 1548.380 ;
        RECT 2959.500 1548.370 2962.500 1548.380 ;
        RECT -42.880 1461.380 -39.880 1461.390 ;
        RECT 2959.500 1461.380 2962.500 1461.390 ;
        RECT -42.880 1458.380 0.300 1461.380 ;
        RECT 2919.700 1458.380 2962.500 1461.380 ;
        RECT -42.880 1458.370 -39.880 1458.380 ;
        RECT 2959.500 1458.370 2962.500 1458.380 ;
        RECT -42.880 1371.380 -39.880 1371.390 ;
        RECT 2959.500 1371.380 2962.500 1371.390 ;
        RECT -42.880 1368.380 0.300 1371.380 ;
        RECT 2919.700 1368.380 2962.500 1371.380 ;
        RECT -42.880 1368.370 -39.880 1368.380 ;
        RECT 2959.500 1368.370 2962.500 1368.380 ;
        RECT -42.880 1281.380 -39.880 1281.390 ;
        RECT 2959.500 1281.380 2962.500 1281.390 ;
        RECT -42.880 1278.380 0.300 1281.380 ;
        RECT 2919.700 1278.380 2962.500 1281.380 ;
        RECT -42.880 1278.370 -39.880 1278.380 ;
        RECT 2959.500 1278.370 2962.500 1278.380 ;
        RECT -42.880 1191.380 -39.880 1191.390 ;
        RECT 2959.500 1191.380 2962.500 1191.390 ;
        RECT -42.880 1188.380 0.300 1191.380 ;
        RECT 2919.700 1188.380 2962.500 1191.380 ;
        RECT -42.880 1188.370 -39.880 1188.380 ;
        RECT 2959.500 1188.370 2962.500 1188.380 ;
        RECT -42.880 1101.380 -39.880 1101.390 ;
        RECT 2959.500 1101.380 2962.500 1101.390 ;
        RECT -42.880 1098.380 0.300 1101.380 ;
        RECT 2919.700 1098.380 2962.500 1101.380 ;
        RECT -42.880 1098.370 -39.880 1098.380 ;
        RECT 2959.500 1098.370 2962.500 1098.380 ;
        RECT -42.880 1011.380 -39.880 1011.390 ;
        RECT 2959.500 1011.380 2962.500 1011.390 ;
        RECT -42.880 1008.380 0.300 1011.380 ;
        RECT 2919.700 1008.380 2962.500 1011.380 ;
        RECT -42.880 1008.370 -39.880 1008.380 ;
        RECT 2959.500 1008.370 2962.500 1008.380 ;
        RECT -42.880 921.380 -39.880 921.390 ;
        RECT 2959.500 921.380 2962.500 921.390 ;
        RECT -42.880 918.380 0.300 921.380 ;
        RECT 2919.700 918.380 2962.500 921.380 ;
        RECT -42.880 918.370 -39.880 918.380 ;
        RECT 2959.500 918.370 2962.500 918.380 ;
        RECT -42.880 831.380 -39.880 831.390 ;
        RECT 2959.500 831.380 2962.500 831.390 ;
        RECT -42.880 828.380 0.300 831.380 ;
        RECT 2919.700 828.380 2962.500 831.380 ;
        RECT -42.880 828.370 -39.880 828.380 ;
        RECT 2959.500 828.370 2962.500 828.380 ;
        RECT -42.880 741.380 -39.880 741.390 ;
        RECT 2959.500 741.380 2962.500 741.390 ;
        RECT -42.880 738.380 0.300 741.380 ;
        RECT 2919.700 738.380 2962.500 741.380 ;
        RECT -42.880 738.370 -39.880 738.380 ;
        RECT 2959.500 738.370 2962.500 738.380 ;
        RECT -42.880 651.380 -39.880 651.390 ;
        RECT 2959.500 651.380 2962.500 651.390 ;
        RECT -42.880 648.380 0.300 651.380 ;
        RECT 2919.700 648.380 2962.500 651.380 ;
        RECT -42.880 648.370 -39.880 648.380 ;
        RECT 2959.500 648.370 2962.500 648.380 ;
        RECT -42.880 561.380 -39.880 561.390 ;
        RECT 2959.500 561.380 2962.500 561.390 ;
        RECT -42.880 558.380 0.300 561.380 ;
        RECT 2919.700 558.380 2962.500 561.380 ;
        RECT -42.880 558.370 -39.880 558.380 ;
        RECT 2959.500 558.370 2962.500 558.380 ;
        RECT -42.880 471.380 -39.880 471.390 ;
        RECT 2959.500 471.380 2962.500 471.390 ;
        RECT -42.880 468.380 0.300 471.380 ;
        RECT 2919.700 468.380 2962.500 471.380 ;
        RECT -42.880 468.370 -39.880 468.380 ;
        RECT 2959.500 468.370 2962.500 468.380 ;
        RECT -42.880 381.380 -39.880 381.390 ;
        RECT 2959.500 381.380 2962.500 381.390 ;
        RECT -42.880 378.380 0.300 381.380 ;
        RECT 2919.700 378.380 2962.500 381.380 ;
        RECT -42.880 378.370 -39.880 378.380 ;
        RECT 2959.500 378.370 2962.500 378.380 ;
        RECT -42.880 291.380 -39.880 291.390 ;
        RECT 2959.500 291.380 2962.500 291.390 ;
        RECT -42.880 288.380 0.300 291.380 ;
        RECT 2919.700 288.380 2962.500 291.380 ;
        RECT -42.880 288.370 -39.880 288.380 ;
        RECT 2959.500 288.370 2962.500 288.380 ;
        RECT -42.880 201.380 -39.880 201.390 ;
        RECT 2959.500 201.380 2962.500 201.390 ;
        RECT -42.880 198.380 0.300 201.380 ;
        RECT 2919.700 198.380 2962.500 201.380 ;
        RECT -42.880 198.370 -39.880 198.380 ;
        RECT 2959.500 198.370 2962.500 198.380 ;
        RECT -42.880 111.380 -39.880 111.390 ;
        RECT 2959.500 111.380 2962.500 111.390 ;
        RECT -42.880 108.380 0.300 111.380 ;
        RECT 2919.700 108.380 2962.500 111.380 ;
        RECT -42.880 108.370 -39.880 108.380 ;
        RECT 2959.500 108.370 2962.500 108.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 103.020 -34.520 106.020 -34.510 ;
        RECT 193.020 -34.520 196.020 -34.510 ;
        RECT 283.020 -34.520 286.020 -34.510 ;
        RECT 373.020 -34.520 376.020 -34.510 ;
        RECT 463.020 -34.520 466.020 -34.510 ;
        RECT 553.020 -34.520 556.020 -34.510 ;
        RECT 643.020 -34.520 646.020 -34.510 ;
        RECT 733.020 -34.520 736.020 -34.510 ;
        RECT 823.020 -34.520 826.020 -34.510 ;
        RECT 913.020 -34.520 916.020 -34.510 ;
        RECT 1003.020 -34.520 1006.020 -34.510 ;
        RECT 1093.020 -34.520 1096.020 -34.510 ;
        RECT 1183.020 -34.520 1186.020 -34.510 ;
        RECT 1273.020 -34.520 1276.020 -34.510 ;
        RECT 1363.020 -34.520 1366.020 -34.510 ;
        RECT 1453.020 -34.520 1456.020 -34.510 ;
        RECT 1543.020 -34.520 1546.020 -34.510 ;
        RECT 1633.020 -34.520 1636.020 -34.510 ;
        RECT 1723.020 -34.520 1726.020 -34.510 ;
        RECT 1813.020 -34.520 1816.020 -34.510 ;
        RECT 1903.020 -34.520 1906.020 -34.510 ;
        RECT 1993.020 -34.520 1996.020 -34.510 ;
        RECT 2083.020 -34.520 2086.020 -34.510 ;
        RECT 2173.020 -34.520 2176.020 -34.510 ;
        RECT 2263.020 -34.520 2266.020 -34.510 ;
        RECT 2353.020 -34.520 2356.020 -34.510 ;
        RECT 2443.020 -34.520 2446.020 -34.510 ;
        RECT 2533.020 -34.520 2536.020 -34.510 ;
        RECT 2623.020 -34.520 2626.020 -34.510 ;
        RECT 2713.020 -34.520 2716.020 -34.510 ;
        RECT 2803.020 -34.520 2806.020 -34.510 ;
        RECT 2893.020 -34.520 2896.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 103.020 -37.530 106.020 -37.520 ;
        RECT 193.020 -37.530 196.020 -37.520 ;
        RECT 283.020 -37.530 286.020 -37.520 ;
        RECT 373.020 -37.530 376.020 -37.520 ;
        RECT 463.020 -37.530 466.020 -37.520 ;
        RECT 553.020 -37.530 556.020 -37.520 ;
        RECT 643.020 -37.530 646.020 -37.520 ;
        RECT 733.020 -37.530 736.020 -37.520 ;
        RECT 823.020 -37.530 826.020 -37.520 ;
        RECT 913.020 -37.530 916.020 -37.520 ;
        RECT 1003.020 -37.530 1006.020 -37.520 ;
        RECT 1093.020 -37.530 1096.020 -37.520 ;
        RECT 1183.020 -37.530 1186.020 -37.520 ;
        RECT 1273.020 -37.530 1276.020 -37.520 ;
        RECT 1363.020 -37.530 1366.020 -37.520 ;
        RECT 1453.020 -37.530 1456.020 -37.520 ;
        RECT 1543.020 -37.530 1546.020 -37.520 ;
        RECT 1633.020 -37.530 1636.020 -37.520 ;
        RECT 1723.020 -37.530 1726.020 -37.520 ;
        RECT 1813.020 -37.530 1816.020 -37.520 ;
        RECT 1903.020 -37.530 1906.020 -37.520 ;
        RECT 1993.020 -37.530 1996.020 -37.520 ;
        RECT 2083.020 -37.530 2086.020 -37.520 ;
        RECT 2173.020 -37.530 2176.020 -37.520 ;
        RECT 2263.020 -37.530 2266.020 -37.520 ;
        RECT 2353.020 -37.530 2356.020 -37.520 ;
        RECT 2443.020 -37.530 2446.020 -37.520 ;
        RECT 2533.020 -37.530 2536.020 -37.520 ;
        RECT 2623.020 -37.530 2626.020 -37.520 ;
        RECT 2713.020 -37.530 2716.020 -37.520 ;
        RECT 2803.020 -37.530 2806.020 -37.520 ;
        RECT 2893.020 -37.530 2896.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 2.805 2910.420 3506.165 ;
      LAYER met1 ;
        RECT 2.830 2.760 2914.100 3509.040 ;
      LAYER met2 ;
        RECT 2.710 0.300 2917.370 3519.700 ;
      LAYER met3 ;
        RECT 0.300 10.715 2919.700 3508.965 ;
      LAYER met4 ;
        RECT 4.020 0.300 2905.020 3519.700 ;
      LAYER met5 ;
        RECT 0.300 9.130 2919.700 3495.390 ;
  END
END user_project_wrapper
END LIBRARY

