*---------------------------------------------------------------------------
* SPDX-FileCopyrightText: 2020 Efabless Corporation
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*---------------------------------------------------------------------------
* NGSPICE file created from ycell.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

.subckt ycell cbitin cbitout confclk confclko dempty din[0] din[1] dout[0] dout[1]
+ hempty hempty2 lempty lin[0] lin[1] lout[0] lout[1] rempty reset reseto rin[0] rin[1]
+ rout[0] rout[1] uempty uin[0] uin[1] uout[0] uout[1] vempty vempty2 vccd1 vssd1
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_131_ _068_/A _133_/X _121_/Y _121_/A _155_/D vssd1 vssd1 vccd1 vccd1 rout[1] sky130_fd_sc_hd__a32o_4
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_114_ _070_/A _155_/C _108_/Y vssd1 vssd1 vccd1 vccd1 _070_/A sky130_fd_sc_hd__o21a_4
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_130_ _129_/X vssd1 vssd1 vccd1 vccd1 _155_/D sky130_fd_sc_hd__inv_4
XFILLER_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_113_ lin[0] _113_/B vssd1 vssd1 vccd1 vccd1 _155_/C sky130_fd_sc_hd__and2_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_112_ lempty vssd1 vssd1 vccd1 vccd1 _113_/B sky130_fd_sc_hd__inv_2
XFILLER_13_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_111_ _068_/A _110_/Y _108_/Y vssd1 vssd1 vccd1 vccd1 _068_/A sky130_fd_sc_hd__o21a_4
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_110_ _106_/Y _082_/A vssd1 vssd1 vccd1 vccd1 _110_/Y sky130_fd_sc_hd__nor2_4
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_099_ _137_/B vssd1 vssd1 vccd1 vccd1 _099_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_098_ _137_/A _152_/X vssd1 vssd1 vccd1 vccd1 _098_/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_097_ _087_/Y dout[1] din[1] _087_/A vssd1 vssd1 vccd1 vccd1 uout[1] sky130_fd_sc_hd__o22a_4
XFILLER_19_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_149_ _137_/B _147_/Y _148_/Y vssd1 vssd1 vccd1 vccd1 _137_/B sky130_fd_sc_hd__o21a_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_148_ _136_/X vssd1 vssd1 vccd1 vccd1 _148_/Y sky130_fd_sc_hd__inv_2
X_096_ _137_/A _153_/X _090_/Y _090_/A _134_/D vssd1 vssd1 vccd1 vccd1 dout[1] sky130_fd_sc_hd__a32o_4
XFILLER_1_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_079_ _073_/X _163_/Q _138_/C vssd1 vssd1 vccd1 vccd1 _079_/X sky130_fd_sc_hd__or3_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_095_ _091_/Y _085_/A _094_/Y _092_/Y uin[1] vssd1 vssd1 vccd1 vccd1 _134_/D sky130_fd_sc_hd__a32o_4
X_164_ confclk _163_/Q vssd1 vssd1 vccd1 vccd1 cbitout sky130_fd_sc_hd__dfxtp_4
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_078_ uout[1] vssd1 vssd1 vccd1 vccd1 _078_/Y sky130_fd_sc_hd__inv_2
X_147_ _150_/A _142_/X vssd1 vssd1 vccd1 vccd1 _147_/Y sky130_fd_sc_hd__nor2_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_094_ _093_/X vssd1 vssd1 vccd1 vccd1 _094_/Y sky130_fd_sc_hd__inv_2
X_163_ confclk _162_/Q vssd1 vssd1 vccd1 vccd1 _163_/Q sky130_fd_sc_hd__dfxtp_4
X_129_ lempty _122_/Y lout[0] _128_/X vssd1 vssd1 vccd1 vccd1 _129_/X sky130_fd_sc_hd__o22a_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_146_ _146_/A vssd1 vssd1 vccd1 vccd1 _134_/A sky130_fd_sc_hd__inv_2
X_077_ _138_/A _163_/Q _138_/C vssd1 vssd1 vccd1 vccd1 _077_/X sky130_fd_sc_hd__or3_4
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_162_ confclk cbitin vssd1 vssd1 vccd1 vccd1 _162_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_13_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_093_ _092_/Y dempty uout[1] uout[0] vssd1 vssd1 vccd1 vccd1 _093_/X sky130_fd_sc_hd__or4_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_076_ _076_/A vssd1 vssd1 vccd1 vccd1 _138_/C sky130_fd_sc_hd__buf_2
X_145_ _137_/X _141_/X _142_/X _150_/A _144_/X vssd1 vssd1 vccd1 vccd1 _146_/A sky130_fd_sc_hd__a32o_4
XFILLER_16_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_128_ _113_/B rempty lout[1] _157_/A vssd1 vssd1 vccd1 vccd1 _128_/X sky130_fd_sc_hd__or4_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_092_ uempty vssd1 vssd1 vccd1 vccd1 _092_/Y sky130_fd_sc_hd__inv_2
X_161_ vempty vssd1 vssd1 vccd1 vccd1 vempty2 sky130_fd_sc_hd__buf_2
XFILLER_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_144_ _152_/X _153_/X _137_/A _137_/B vssd1 vssd1 vccd1 vccd1 _144_/X sky130_fd_sc_hd__or4_4
X_127_ reset hempty vssd1 vssd1 vccd1 vccd1 _157_/A sky130_fd_sc_hd__or2_4
X_075_ cbitout vssd1 vssd1 vccd1 vccd1 _076_/A sky130_fd_sc_hd__inv_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_091_ reset vssd1 vssd1 vccd1 vccd1 _091_/Y sky130_fd_sc_hd__inv_2
X_074_ _073_/X vssd1 vssd1 vccd1 vccd1 _138_/A sky130_fd_sc_hd__inv_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_160_ reset vssd1 vssd1 vccd1 vccd1 reseto sky130_fd_sc_hd__buf_2
X_143_ _134_/A vssd1 vssd1 vccd1 vccd1 _150_/A sky130_fd_sc_hd__inv_2
XFILLER_16_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_126_ _125_/Y vssd1 vssd1 vccd1 vccd1 lout[0] sky130_fd_sc_hd__inv_4
X_109_ _069_/A _107_/Y _108_/Y vssd1 vssd1 vccd1 vccd1 _069_/A sky130_fd_sc_hd__o21a_4
XFILLER_13_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_090_ _090_/A vssd1 vssd1 vccd1 vccd1 _090_/Y sky130_fd_sc_hd__inv_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_073_ _162_/Q vssd1 vssd1 vccd1 vccd1 _073_/X sky130_fd_sc_hd__buf_4
X_125_ _117_/X rout[0] rin[0] _118_/Y vssd1 vssd1 vccd1 vccd1 _125_/Y sky130_fd_sc_hd__a22oi_4
X_142_ _125_/Y _140_/X _139_/Y _138_/X vssd1 vssd1 vccd1 vccd1 _142_/X sky130_fd_sc_hd__o22a_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_108_ _157_/X vssd1 vssd1 vccd1 vccd1 _108_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_072_ uout[0] vssd1 vssd1 vccd1 vccd1 _072_/Y sky130_fd_sc_hd__inv_2
X_141_ _125_/Y _138_/X _139_/Y _140_/X vssd1 vssd1 vccd1 vccd1 _141_/X sky130_fd_sc_hd__o22a_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_124_ _155_/C _121_/Y _121_/A _123_/X vssd1 vssd1 vccd1 vccd1 rout[0] sky130_fd_sc_hd__o22a_4
XFILLER_2_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_107_ _106_/Y _107_/B vssd1 vssd1 vccd1 vccd1 _107_/Y sky130_fd_sc_hd__nor2_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_071_ _106_/A _155_/B vssd1 vssd1 vccd1 vccd1 _071_/X sky130_fd_sc_hd__or2_4
X_140_ _073_/X _138_/B _138_/C vssd1 vssd1 vccd1 vccd1 _140_/X sky130_fd_sc_hd__or3_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_106_ _106_/A vssd1 vssd1 vccd1 vccd1 _106_/Y sky130_fd_sc_hd__inv_2
X_123_ _069_/Y _155_/B _068_/A _070_/A vssd1 vssd1 vccd1 vccd1 _123_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_070_ _070_/A _133_/X vssd1 vssd1 vccd1 vccd1 _155_/B sky130_fd_sc_hd__nor2_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_122_ lin[1] vssd1 vssd1 vccd1 vccd1 _122_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_105_ _087_/Y _104_/X din[0] _087_/Y vssd1 vssd1 vccd1 vccd1 uout[0] sky130_fd_sc_hd__a2bb2o_4
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_121_ _121_/A vssd1 vssd1 vccd1 vccd1 _121_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_104_ _090_/Y _098_/Y _101_/X _090_/A _103_/Y vssd1 vssd1 vccd1 vccd1 _104_/X sky130_fd_sc_hd__a32o_4
XFILLER_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_120_ _073_/X _138_/B _138_/C _090_/Y _119_/X vssd1 vssd1 vccd1 vccd1 _121_/A sky130_fd_sc_hd__a32o_4
X_103_ _102_/X vssd1 vssd1 vccd1 vccd1 _103_/Y sky130_fd_sc_hd__inv_2
XPHY_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_102_ uin[0] _092_/Y vssd1 vssd1 vccd1 vccd1 _102_/X sky130_fd_sc_hd__and2_4
XFILLER_17_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_101_ _099_/Y _134_/C vssd1 vssd1 vccd1 vccd1 _101_/X sky130_fd_sc_hd__or2_4
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_100_ _152_/X _153_/X vssd1 vssd1 vccd1 vccd1 _134_/C sky130_fd_sc_hd__nor2_4
XFILLER_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_159_ hempty vssd1 vssd1 vccd1 vccd1 hempty2 sky130_fd_sc_hd__buf_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_089_ _138_/B _076_/A _085_/A vssd1 vssd1 vccd1 vccd1 _090_/A sky130_fd_sc_hd__o21a_4
X_158_ confclk vssd1 vssd1 vccd1 vccd1 confclko sky130_fd_sc_hd__buf_2
XFILLER_0_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_157_ _157_/A _156_/Y vssd1 vssd1 vccd1 vccd1 _157_/X sky130_fd_sc_hd__or2_4
X_088_ _163_/Q vssd1 vssd1 vccd1 vccd1 _138_/B sky130_fd_sc_hd__inv_2
XFILLER_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_156_ _156_/A vssd1 vssd1 vccd1 vccd1 _156_/Y sky130_fd_sc_hd__inv_2
X_087_ _087_/A vssd1 vssd1 vccd1 vccd1 _087_/Y sky130_fd_sc_hd__inv_2
X_139_ lout[1] vssd1 vssd1 vccd1 vccd1 _139_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_155_ _106_/A _155_/B _155_/C _155_/D vssd1 vssd1 vccd1 vccd1 _156_/A sky130_fd_sc_hd__or4_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_086_ dempty vempty vssd1 vssd1 vccd1 vccd1 _087_/A sky130_fd_sc_hd__or2_4
X_069_ _069_/A vssd1 vssd1 vccd1 vccd1 _069_/Y sky130_fd_sc_hd__inv_2
X_138_ _138_/A _138_/B _138_/C vssd1 vssd1 vccd1 vccd1 _138_/X sky130_fd_sc_hd__or3_4
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_47 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_085_ _085_/A vssd1 vssd1 vccd1 vccd1 vempty sky130_fd_sc_hd__inv_2
X_154_ _104_/X vssd1 vssd1 vccd1 vccd1 dout[0] sky130_fd_sc_hd__inv_2
XFILLER_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_068_ _068_/A vssd1 vssd1 vccd1 vccd1 _068_/Y sky130_fd_sc_hd__inv_2
X_137_ _137_/A _137_/B vssd1 vssd1 vccd1 vccd1 _137_/X sky130_fd_sc_hd__or2_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_084_ _162_/Q cbitout vssd1 vssd1 vccd1 vccd1 _085_/A sky130_fd_sc_hd__or2_4
X_153_ _153_/X _134_/D _148_/Y vssd1 vssd1 vccd1 vccd1 _153_/X sky130_fd_sc_hd__o21a_4
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_136_ reset vempty _135_/Y vssd1 vssd1 vccd1 vccd1 _136_/X sky130_fd_sc_hd__or3_4
X_119_ _163_/Q cbitout vssd1 vssd1 vccd1 vccd1 _119_/X sky130_fd_sc_hd__or2_4
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_152_ _152_/X _102_/X _148_/Y vssd1 vssd1 vccd1 vccd1 _152_/X sky130_fd_sc_hd__o21a_4
X_083_ _068_/Y _069_/Y _071_/X _106_/A _082_/Y vssd1 vssd1 vccd1 vccd1 _106_/A sky130_fd_sc_hd__a32o_4
XFILLER_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_118_ _117_/X vssd1 vssd1 vccd1 vccd1 _118_/Y sky130_fd_sc_hd__inv_2
X_135_ _135_/A vssd1 vssd1 vccd1 vccd1 _135_/Y sky130_fd_sc_hd__inv_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_134_ _134_/A _102_/X _134_/C _134_/D vssd1 vssd1 vccd1 vccd1 _135_/A sky130_fd_sc_hd__or4_4
X_082_ _082_/A _107_/B vssd1 vssd1 vccd1 vccd1 _082_/Y sky130_fd_sc_hd__nand2_4
X_151_ _137_/A _150_/Y _148_/Y vssd1 vssd1 vccd1 vccd1 _137_/A sky130_fd_sc_hd__o21a_4
XFILLER_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_117_ rempty hempty vssd1 vssd1 vccd1 vccd1 _117_/X sky130_fd_sc_hd__or2_4
XFILLER_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_081_ _072_/Y _079_/X _078_/Y _077_/X vssd1 vssd1 vccd1 vccd1 _107_/B sky130_fd_sc_hd__o22a_4
X_150_ _150_/A _141_/X vssd1 vssd1 vccd1 vccd1 _150_/Y sky130_fd_sc_hd__nor2_4
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_133_ _133_/X _155_/D _108_/Y vssd1 vssd1 vccd1 vccd1 _133_/X sky130_fd_sc_hd__o21a_4
XFILLER_0_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_116_ cbitout _116_/B vssd1 vssd1 vccd1 vccd1 hempty sky130_fd_sc_hd__nor2_4
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_080_ _072_/Y _077_/X _078_/Y _079_/X vssd1 vssd1 vccd1 vccd1 _082_/A sky130_fd_sc_hd__o22a_4
X_132_ _118_/Y rout[1] rin[1] _117_/X vssd1 vssd1 vccd1 vccd1 lout[1] sky130_fd_sc_hd__o22a_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_115_ _073_/X _163_/Q _138_/A _138_/B vssd1 vssd1 vccd1 vccd1 _116_/B sky130_fd_sc_hd__o22a_4
XFILLER_0_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
.ends

