// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module mprj2_logic_high(HI, vccd2, vssd2);
  output HI;
  input vccd2;
  input vssd2;
  sky130_fd_sc_hd__decap_12 FILLER_0_106 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_118 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_125 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_137 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_149 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_15 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_156 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_168 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_180 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_187 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_199 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_211 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_218 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_230 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_242 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_0_249 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_27 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_3 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_32 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_44 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_56 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_63 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_75 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_0_87 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_0_94 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_110 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_123 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_135 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_14 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_147 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_159 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_171 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_184 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_196 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_208 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_220 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_232 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_245 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_26 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_3 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_38 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_50 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_58 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_62 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_74 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_86 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_98 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_106 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_118 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_125 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_137 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_149 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_15 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_156 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_168 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_180 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_187 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_199 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_211 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_218 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_230 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_242 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_249 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_27 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_3 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_32 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_44 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_56 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_63 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_75 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_87 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_94 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_18 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_19 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_20 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_21 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_22 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_23 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_24 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_25 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9 (
    .VGND(vssd2),
    .VPWR(vccd2)
  );
  sky130_fd_sc_hd__conb_1 inst (
    .HI(HI),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2)
  );
endmodule
