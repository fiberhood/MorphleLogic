magic
tech sky130A
magscale 1 2
timestamp 1608069679
<< locali >>
rect 299857 666587 299891 684437
rect 364349 666587 364383 676141
rect 429577 666587 429611 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 299673 601715 299707 608549
rect 429393 601715 429427 608549
rect 559113 601715 559147 608549
rect 299857 589339 299891 598893
rect 429577 589339 429611 598893
rect 559297 589339 559331 598893
rect 299581 550647 299615 560201
rect 429209 550647 429243 553401
rect 559021 550647 559055 560201
rect 19349 542963 19383 543065
rect 12449 542827 12483 542929
rect 28917 542895 28951 543065
rect 38669 542963 38703 543065
rect 31769 542827 31803 542929
rect 48237 542895 48271 543065
rect 57989 542963 58023 543065
rect 51089 542827 51123 542929
rect 67557 542895 67591 543065
rect 77309 542963 77343 543065
rect 70409 542827 70443 542929
rect 86877 542895 86911 543065
rect 96629 542963 96663 543065
rect 89729 542827 89763 542929
rect 106197 542895 106231 543065
rect 115949 542963 115983 543065
rect 109049 542827 109083 542929
rect 125517 542895 125551 543065
rect 144929 543031 144963 543133
rect 137971 542929 138029 542963
rect 128369 542827 128403 542929
rect 154497 542895 154531 543133
rect 154681 542895 154715 542929
rect 154623 542861 154715 542895
rect 161857 542895 161891 544697
rect 164065 543983 164099 544697
rect 169585 544119 169619 544697
rect 172161 544187 172195 544697
rect 174921 544323 174955 544697
rect 180073 544391 180107 544697
rect 182649 544459 182683 544697
rect 195529 544527 195563 544697
rect 200681 544595 200715 544697
rect 412189 544255 412223 544629
rect 417341 544051 417375 544629
rect 427829 543915 427863 544629
rect 432797 543847 432831 544629
rect 438225 543711 438259 544629
rect 443101 543779 443135 544629
rect 164249 542963 164283 543201
rect 168849 542895 168883 542997
rect 168941 542895 168975 543201
rect 173817 542895 173851 542997
rect 173909 542895 173943 543065
rect 176485 542895 176519 543133
rect 178693 542895 178727 543065
rect 183477 542963 183511 543133
rect 183569 542963 183603 543201
rect 188169 542895 188203 542997
rect 188261 542895 188295 543201
rect 193137 542895 193171 542997
rect 193229 542895 193263 543065
rect 193321 542895 193355 543133
rect 198013 542895 198047 543065
rect 202797 542963 202831 543133
rect 202889 542963 202923 543201
rect 207489 542895 207523 542997
rect 207581 542895 207615 543201
rect 211169 542895 211203 543133
rect 215769 542895 215803 542997
rect 220737 542963 220771 543133
rect 249809 543099 249843 543201
rect 259377 543031 259411 543201
rect 263701 542895 263735 542929
rect 241563 542861 241713 542895
rect 263551 542861 263735 542895
rect 265173 542895 265207 542997
rect 270509 542895 270543 543065
rect 273085 542895 273119 543133
rect 275293 542895 275327 543065
rect 280077 542963 280111 543133
rect 280169 542963 280203 543201
rect 284769 542895 284803 542997
rect 284861 542895 284895 543201
rect 289737 542895 289771 542997
rect 289829 542895 289863 543065
rect 292405 542895 292439 543133
rect 294613 542895 294647 543065
rect 299397 542963 299431 543133
rect 299489 542895 299523 543133
rect 308873 542895 308907 543133
rect 309149 542895 309183 543065
rect 308873 542861 309057 542895
rect 311725 542895 311759 543133
rect 313933 542895 313967 543065
rect 318717 542963 318751 543133
rect 318809 542963 318843 543201
rect 323409 542895 323443 542997
rect 323501 542895 323535 543201
rect 327089 542895 327123 543065
rect 328503 542997 328595 543031
rect 328561 542963 328595 542997
rect 346593 542963 346627 543133
rect 355977 543031 356011 543133
rect 424977 543099 425011 543201
rect 365821 542895 365855 542997
rect 369777 542997 370053 543031
rect 389131 542997 389189 543031
rect 398791 542997 398941 543031
rect 369777 542895 369811 542997
rect 48329 242811 48363 242913
rect 57897 242743 57931 242913
rect 67649 242811 67683 242913
rect 77217 242743 77251 242913
rect 60691 242709 60749 242743
rect 82093 242743 82127 242913
rect 86877 242539 86911 242913
rect 132509 242811 132543 242913
rect 89637 242539 89671 242777
rect 94513 242539 94547 242777
rect 103529 241791 103563 242505
rect 113097 241791 113131 242505
rect 113189 241723 113223 242777
rect 122757 241723 122791 242777
rect 142261 242539 142295 242913
rect 122699 241689 122791 241723
rect 152473 242539 152507 242777
rect 142169 241519 142203 242505
rect 152565 241519 152599 242505
rect 162133 242335 162167 242777
rect 171793 242335 171827 242845
rect 178785 242675 178819 242845
rect 183293 242845 183511 242879
rect 183293 242743 183327 242845
rect 183477 242811 183511 242845
rect 183569 242675 183603 243049
rect 184213 242743 184247 242981
rect 190653 242879 190687 243049
rect 200773 242675 200807 242845
rect 273177 242811 273211 242913
rect 220093 242131 220127 242777
rect 238493 242199 238527 242301
rect 238401 241587 238435 242165
rect 261493 241927 261527 242777
rect 267657 242607 267691 242777
rect 238677 241519 238711 241757
rect 268301 241519 268335 242573
rect 268393 241519 268427 242029
rect 271337 241655 271371 242709
rect 276765 242267 276799 242709
rect 341993 242471 342027 242641
rect 342913 242539 342947 242913
rect 345673 242199 345707 242505
rect 345949 241995 345983 242845
rect 347697 242607 347731 242913
rect 350215 242845 350365 242879
rect 350365 242777 350457 242811
rect 350365 242743 350399 242777
rect 350583 242641 350767 242675
rect 274373 241587 274407 241825
rect 344017 241655 344051 241893
rect 344109 241723 344143 241893
rect 350549 241723 350583 242505
rect 344201 241655 344235 241689
rect 344017 241621 344235 241655
rect 350641 241519 350675 242505
rect 350733 241927 350767 242641
rect 350825 242607 350859 242913
rect 355241 241927 355275 242437
rect 355425 242267 355459 243185
rect 364625 242471 364659 242777
rect 367235 242709 367327 242743
rect 367293 242675 367327 242709
rect 367235 242573 367385 242607
rect 350733 241893 350917 241927
rect 350583 241485 350675 241519
rect 353309 241519 353343 241689
rect 355149 241451 355183 241893
rect 355333 241791 355367 242233
rect 367201 241587 367235 242437
rect 369225 242335 369259 242437
rect 369961 241519 369995 242913
rect 370053 242335 370087 242777
rect 379529 242743 379563 242845
rect 379529 242641 379621 242675
rect 379529 242199 379563 242641
rect 412775 242437 412925 242471
rect 379621 241791 379655 242165
rect 379563 241757 379655 241791
rect 393973 241655 394007 242097
rect 394249 241791 394283 242369
rect 414029 242335 414063 242505
rect 418169 242335 418203 242913
rect 431911 242573 432003 242607
rect 422953 242471 422987 242573
rect 431969 242471 432003 242573
rect 395537 241859 395571 242165
rect 412833 242131 412867 242233
rect 418261 242131 418295 242233
rect 418353 241519 418387 242233
rect 450001 242131 450035 242777
rect 419549 241519 419583 242097
rect 442641 242097 443101 242131
rect 442641 242063 442675 242097
rect 154865 222207 154899 224961
rect 156153 222207 156187 224961
rect 169953 222207 169987 227001
rect 194977 226355 195011 235909
rect 198289 231863 198323 241417
rect 237665 231863 237699 239377
rect 303813 231863 303847 241417
rect 423229 239275 423263 241417
rect 191941 222207 191975 224961
rect 278881 222207 278915 225029
rect 223865 220847 223899 222173
rect 403541 222207 403575 231761
rect 423229 222207 423263 224961
rect 225153 220847 225187 222173
rect 178233 212551 178267 215237
rect 179521 212551 179555 215373
rect 216965 211123 216999 219385
rect 214021 202895 214055 209797
rect 218253 205615 218287 219385
rect 263793 212551 263827 215237
rect 265081 212551 265115 215373
rect 270601 212551 270635 215373
rect 272073 212551 272107 215237
rect 424701 212551 424735 222105
rect 384681 205615 384715 211089
rect 423229 202895 423263 205649
rect 150725 183583 150759 201433
rect 218253 193171 218287 201433
rect 248153 191879 248187 201433
rect 423229 193307 423263 202725
rect 150725 173723 150759 182121
rect 190745 173927 190779 183481
rect 192033 173927 192067 183413
rect 196265 179435 196299 188989
rect 423137 183583 423171 186337
rect 218253 180047 218287 183413
rect 219541 180047 219575 183481
rect 194793 169779 194827 179333
rect 238493 172567 238527 182121
rect 384589 176647 384623 182121
rect 424517 173859 424551 182121
rect 156153 154615 156187 164169
rect 174001 157335 174035 164169
rect 194793 158763 194827 168317
rect 150817 131155 150851 140709
rect 152197 131155 152231 140709
rect 162961 137955 162995 143497
rect 174001 137955 174035 144857
rect 189273 133943 189307 143497
rect 194701 140811 194735 150365
rect 198289 149107 198323 158661
rect 206017 157335 206051 162809
rect 219541 162435 219575 171037
rect 216781 151827 216815 161381
rect 219541 150467 219575 160021
rect 236285 157267 236319 164169
rect 237573 157267 237607 164169
rect 248337 153255 248371 162809
rect 252753 157335 252787 164169
rect 284401 157335 284435 164169
rect 307953 157335 307987 164169
rect 346225 157335 346259 164169
rect 357265 157335 357299 164169
rect 423229 162911 423263 172465
rect 263793 148359 263827 154513
rect 374285 153255 374319 162809
rect 379069 157335 379103 162809
rect 384589 153255 384623 162809
rect 424701 157335 424735 162809
rect 153393 124219 153427 133841
rect 156153 124219 156187 133841
rect 168849 124219 168883 133841
rect 150725 103547 150759 116297
rect 152013 111843 152047 121397
rect 162961 114563 162995 124117
rect 174001 118643 174035 125545
rect 178233 115991 178267 125545
rect 192033 124151 192067 132413
rect 216781 129727 216815 135201
rect 234813 124287 234847 133841
rect 238677 125647 238711 143497
rect 248337 133943 248371 143497
rect 252753 137955 252787 144857
rect 245761 124219 245795 133841
rect 263793 132515 263827 142069
rect 284401 137955 284435 144857
rect 307953 137955 307987 144857
rect 346225 137955 346259 144857
rect 357265 137955 357299 144857
rect 423229 143599 423263 153153
rect 374285 133943 374319 143497
rect 379161 132515 379195 142069
rect 424701 137955 424735 143497
rect 189273 114563 189307 124117
rect 234813 114563 234847 124117
rect 238585 114563 238619 124117
rect 248337 114563 248371 124117
rect 252753 118643 252787 125545
rect 153301 104907 153335 114393
rect 168849 106267 168883 114461
rect 191941 111843 191975 113237
rect 152013 92531 152047 102085
rect 154773 96747 154807 106165
rect 168849 95251 168883 104805
rect 174001 99331 174035 106233
rect 178233 96679 178267 106233
rect 190653 101371 190687 106233
rect 207029 104907 207063 114461
rect 263793 114291 263827 122757
rect 264989 113203 265023 122757
rect 284401 118643 284435 125545
rect 307953 118643 307987 125545
rect 346225 118643 346259 125545
rect 357265 118643 357299 125545
rect 374285 114563 374319 124117
rect 379161 122859 379195 132345
rect 384681 127823 384715 133841
rect 424701 124287 424735 133841
rect 208409 104907 208443 106301
rect 245761 104907 245795 109701
rect 152013 73219 152047 82773
rect 150725 64855 150759 70261
rect 154773 67643 154807 77197
rect 162961 75939 162995 85493
rect 169769 77299 169803 86921
rect 174001 77299 174035 86921
rect 178233 77299 178267 86921
rect 188997 85595 189031 95149
rect 206017 93891 206051 103445
rect 208409 95115 208443 103445
rect 223773 95251 223807 104805
rect 238677 95251 238711 104805
rect 248337 95251 248371 104805
rect 252753 99331 252787 106233
rect 263793 96883 263827 104805
rect 190653 80699 190687 86921
rect 191941 75939 191975 86921
rect 206017 85595 206051 86989
rect 211353 85595 211387 95149
rect 216873 85595 216907 95149
rect 218345 85595 218379 95149
rect 219633 85595 219667 95149
rect 270509 93891 270543 103445
rect 272073 93891 272107 103445
rect 284401 99331 284435 106233
rect 307953 99331 307987 106233
rect 346225 99331 346259 106233
rect 357265 99331 357299 106233
rect 384589 104907 384623 114393
rect 423229 113203 423263 122757
rect 424701 114563 424735 124117
rect 423045 104907 423079 109701
rect 374285 95251 374319 104805
rect 226625 92531 226659 93789
rect 194885 74579 194919 84133
rect 190653 66283 190687 70465
rect 207029 66283 207063 84133
rect 208501 66351 208535 84133
rect 223773 74579 223807 85493
rect 154773 48399 154807 57885
rect 162869 56627 162903 66181
rect 168481 56627 168515 66181
rect 211261 64991 211295 74477
rect 174001 48331 174035 57885
rect 178233 48331 178267 57885
rect 154773 43707 154807 48229
rect 189181 46971 189215 64821
rect 190653 56627 190687 64617
rect 192033 53839 192067 55301
rect 194701 53839 194735 55233
rect 198197 53839 198231 63461
rect 207121 56355 207155 64821
rect 208501 55267 208535 64821
rect 211353 55267 211387 64821
rect 168573 37315 168607 46869
rect 169861 37315 169895 46869
rect 207121 37315 207155 46869
rect 211261 45611 211295 47277
rect 174001 29019 174035 33813
rect 190653 27727 190687 37213
rect 207213 27727 207247 37145
rect 208593 29019 208627 42041
rect 214113 32419 214147 46869
rect 216965 45611 216999 55165
rect 218253 46971 218287 64821
rect 219541 46971 219575 66181
rect 223681 55267 223715 64821
rect 226533 55267 226567 82773
rect 238677 75939 238711 85493
rect 245761 83215 245795 90389
rect 379161 89403 379195 100045
rect 424701 99331 424735 107049
rect 247049 77299 247083 86921
rect 248337 75939 248371 85493
rect 252753 77299 252787 86921
rect 258089 77299 258123 86921
rect 270509 75939 270543 85493
rect 272073 75939 272107 85493
rect 284401 77299 284435 86921
rect 307953 77299 307987 86921
rect 346225 77299 346259 86921
rect 357265 77299 357299 86921
rect 238677 48331 238711 66181
rect 246037 64923 246071 74477
rect 303905 70227 303939 77197
rect 252753 66283 252787 67677
rect 357265 67643 357299 77129
rect 374285 75939 374319 85493
rect 424701 77299 424735 86921
rect 384681 66283 384715 75837
rect 248337 56627 248371 66181
rect 258181 48331 258215 57885
rect 263701 48331 263735 66181
rect 265081 60707 265115 66181
rect 270601 48331 270635 51153
rect 271889 48331 271923 51085
rect 307861 48331 307895 57885
rect 357265 48331 357299 57885
rect 374285 56627 374319 66181
rect 379161 56695 379195 66181
rect 424701 57987 424735 67541
rect 219449 37247 219483 45509
rect 222485 29019 222519 42041
rect 223773 29019 223807 42041
rect 234813 38675 234847 48229
rect 238585 37315 238619 46869
rect 238677 27727 238711 28985
rect 245761 27659 245795 45509
rect 247417 37247 247451 45509
rect 248337 37315 248371 46869
rect 284493 41395 284527 48229
rect 379161 46971 379195 56525
rect 247417 27659 247451 31297
rect 270601 27659 270635 31841
rect 273361 27659 273395 31841
rect 284401 29019 284435 38573
rect 307953 29019 307987 38573
rect 357265 31739 357299 38573
rect 374285 37315 374319 46869
rect 424701 38675 424735 48229
rect 403817 29019 403851 38573
rect 174001 22083 174035 27557
rect 179521 18003 179555 27557
rect 191941 26299 191975 27625
rect 154865 12427 154899 17901
rect 189181 16643 189215 26197
rect 191941 9707 191975 21369
rect 194701 16643 194735 26197
rect 207121 18003 207155 27557
rect 211353 19363 211387 27557
rect 223681 9707 223715 27557
rect 238585 9707 238619 27557
rect 245853 19363 245887 27217
rect 247969 9707 248003 19261
rect 252753 18003 252787 27557
rect 264989 18003 265023 27557
rect 346225 22083 346259 27557
rect 270509 9707 270543 19329
rect 374285 18003 374319 27557
rect 379253 22083 379287 27489
rect 384589 18003 384623 27557
rect 394065 19363 394099 28917
rect 374193 9707 374227 12529
rect 55263 5321 55355 5355
rect 55229 4607 55263 5185
rect 55321 4471 55355 5321
rect 64705 5321 64797 5355
rect 74583 5321 74675 5355
rect 64705 4471 64739 5321
rect 64797 4607 64831 5185
rect 74549 4199 74583 5185
rect 74641 4267 74675 5321
rect 80161 4267 80195 5525
rect 84117 5355 84151 5525
rect 93869 5219 93903 5525
rect 83749 5185 84117 5219
rect 103437 5219 103471 5525
rect 113189 5219 113223 5661
rect 122757 5219 122791 5661
rect 132509 5219 132543 5661
rect 142077 5219 142111 5661
rect 422861 5525 423079 5559
rect 422861 5491 422895 5525
rect 152105 5321 152289 5355
rect 152105 5287 152139 5321
rect 83749 4199 83783 5185
rect 148977 5015 149011 5117
rect 160845 5083 160879 5253
rect 162225 5219 162259 5321
rect 181453 5287 181487 5389
rect 183569 4743 183603 5457
rect 188353 4403 188387 4709
rect 191113 4675 191147 5389
rect 400229 4743 400263 4777
rect 400229 4709 400413 4743
rect 403541 4539 403575 5049
rect 388361 4199 388395 4301
rect 393881 4267 393915 4369
rect 403633 4267 403667 4573
rect 412465 4267 412499 4573
rect 412557 4539 412591 5049
rect 422217 4539 422251 5117
rect 422953 4879 422987 5457
rect 423045 5083 423079 5525
rect 423321 5151 423355 8109
rect 432463 5389 432647 5423
rect 423045 5049 423355 5083
rect 423137 4811 423171 4981
rect 422769 4777 422987 4811
rect 422769 4675 422803 4777
rect 422953 4743 422987 4777
rect 423229 4743 423263 4981
rect 423321 4811 423355 5049
rect 422953 4709 423263 4743
rect 422861 4607 422895 4709
rect 422861 4573 423045 4607
rect 424057 4471 424091 5389
rect 432613 5219 432647 5389
rect 432613 5185 432889 5219
rect 426449 4539 426483 5117
rect 427829 4403 427863 4777
rect 432521 4743 432555 5185
rect 437121 5015 437155 5185
rect 438317 4879 438351 4981
rect 440709 4947 440743 5117
rect 432613 4845 432797 4879
rect 441537 4879 441571 5321
rect 441663 5049 441939 5083
rect 441905 4879 441939 5049
rect 446505 4947 446539 5185
rect 432613 4811 432647 4845
rect 446597 4811 446631 4913
rect 432521 4709 432705 4743
rect 181361 3315 181395 3621
rect 186237 3315 186271 3553
rect 191021 3383 191055 3757
rect 191205 3655 191239 4097
rect 196725 3655 196759 4097
rect 209329 3655 209363 3961
rect 216505 3655 216539 3961
rect 191113 3247 191147 3553
rect 200773 3247 200807 3553
rect 208777 3315 208811 3553
rect 220093 3315 220127 3553
rect 225245 3383 225279 3621
rect 226349 3519 226383 3621
rect 231869 3519 231903 3621
rect 235825 3519 235859 3689
rect 239505 3519 239539 3757
rect 231961 3383 231995 3485
rect 235917 3485 236469 3519
rect 235733 3451 235767 3485
rect 235917 3451 235951 3485
rect 235733 3417 235951 3451
rect 220185 3179 220219 3281
rect 232053 3111 232087 3349
rect 244289 3247 244323 3621
rect 256893 3315 256927 3825
rect 263609 3587 263643 3757
rect 268393 3655 268427 4029
rect 268485 3655 268519 3757
rect 342729 3383 342763 4029
rect 345765 3655 345799 4029
rect 253799 3281 254777 3315
rect 232145 2907 232179 3077
rect 127449 2873 127633 2907
rect 127449 2839 127483 2873
rect 249073 2839 249107 3281
rect 250545 2771 250579 3213
rect 345581 3111 345615 3553
rect 350457 3111 350491 3485
rect 290749 595 290783 2805
rect 386429 2771 386463 2941
rect 395997 2771 396031 2873
rect 374009 595 374043 2669
<< viali >>
rect 299857 684437 299891 684471
rect 429577 684437 429611 684471
rect 299857 666553 299891 666587
rect 364349 676141 364383 676175
rect 364349 666553 364383 666587
rect 559297 684437 559331 684471
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 299673 608549 299707 608583
rect 299673 601681 299707 601715
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 299857 598893 299891 598927
rect 299857 589305 299891 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 299581 560201 299615 560235
rect 559021 560201 559055 560235
rect 299581 550613 299615 550647
rect 429209 553401 429243 553435
rect 429209 550613 429243 550647
rect 559021 550613 559055 550647
rect 161857 544697 161891 544731
rect 144929 543133 144963 543167
rect 19349 543065 19383 543099
rect 12449 542929 12483 542963
rect 19349 542929 19383 542963
rect 28917 543065 28951 543099
rect 38669 543065 38703 543099
rect 28917 542861 28951 542895
rect 31769 542929 31803 542963
rect 38669 542929 38703 542963
rect 48237 543065 48271 543099
rect 12449 542793 12483 542827
rect 57989 543065 58023 543099
rect 48237 542861 48271 542895
rect 51089 542929 51123 542963
rect 57989 542929 58023 542963
rect 67557 543065 67591 543099
rect 31769 542793 31803 542827
rect 77309 543065 77343 543099
rect 67557 542861 67591 542895
rect 70409 542929 70443 542963
rect 77309 542929 77343 542963
rect 86877 543065 86911 543099
rect 51089 542793 51123 542827
rect 96629 543065 96663 543099
rect 86877 542861 86911 542895
rect 89729 542929 89763 542963
rect 96629 542929 96663 542963
rect 106197 543065 106231 543099
rect 70409 542793 70443 542827
rect 115949 543065 115983 543099
rect 106197 542861 106231 542895
rect 109049 542929 109083 542963
rect 115949 542929 115983 542963
rect 125517 543065 125551 543099
rect 89729 542793 89763 542827
rect 144929 542997 144963 543031
rect 154497 543133 154531 543167
rect 125517 542861 125551 542895
rect 128369 542929 128403 542963
rect 137937 542929 137971 542963
rect 138029 542929 138063 542963
rect 109049 542793 109083 542827
rect 154681 542929 154715 542963
rect 154497 542861 154531 542895
rect 154589 542861 154623 542895
rect 164065 544697 164099 544731
rect 169585 544697 169619 544731
rect 172161 544697 172195 544731
rect 174921 544697 174955 544731
rect 180073 544697 180107 544731
rect 182649 544697 182683 544731
rect 195529 544697 195563 544731
rect 200681 544697 200715 544731
rect 200681 544561 200715 544595
rect 412189 544629 412223 544663
rect 195529 544493 195563 544527
rect 182649 544425 182683 544459
rect 180073 544357 180107 544391
rect 174921 544289 174955 544323
rect 412189 544221 412223 544255
rect 417341 544629 417375 544663
rect 172161 544153 172195 544187
rect 169585 544085 169619 544119
rect 417341 544017 417375 544051
rect 427829 544629 427863 544663
rect 164065 543949 164099 543983
rect 427829 543881 427863 543915
rect 432797 544629 432831 544663
rect 432797 543813 432831 543847
rect 438225 544629 438259 544663
rect 443101 544629 443135 544663
rect 443101 543745 443135 543779
rect 438225 543677 438259 543711
rect 164249 543201 164283 543235
rect 168941 543201 168975 543235
rect 164249 542929 164283 542963
rect 168849 542997 168883 543031
rect 161857 542861 161891 542895
rect 168849 542861 168883 542895
rect 183569 543201 183603 543235
rect 176485 543133 176519 543167
rect 173909 543065 173943 543099
rect 168941 542861 168975 542895
rect 173817 542997 173851 543031
rect 173817 542861 173851 542895
rect 173909 542861 173943 542895
rect 183477 543133 183511 543167
rect 176485 542861 176519 542895
rect 178693 543065 178727 543099
rect 183477 542929 183511 542963
rect 188261 543201 188295 543235
rect 183569 542929 183603 542963
rect 188169 542997 188203 543031
rect 178693 542861 178727 542895
rect 188169 542861 188203 542895
rect 202889 543201 202923 543235
rect 193321 543133 193355 543167
rect 193229 543065 193263 543099
rect 188261 542861 188295 542895
rect 193137 542997 193171 543031
rect 193137 542861 193171 542895
rect 193229 542861 193263 542895
rect 202797 543133 202831 543167
rect 193321 542861 193355 542895
rect 198013 543065 198047 543099
rect 202797 542929 202831 542963
rect 207581 543201 207615 543235
rect 202889 542929 202923 542963
rect 207489 542997 207523 543031
rect 198013 542861 198047 542895
rect 207489 542861 207523 542895
rect 249809 543201 249843 543235
rect 207581 542861 207615 542895
rect 211169 543133 211203 543167
rect 220737 543133 220771 543167
rect 211169 542861 211203 542895
rect 215769 542997 215803 543031
rect 249809 543065 249843 543099
rect 259377 543201 259411 543235
rect 280169 543201 280203 543235
rect 273085 543133 273119 543167
rect 270509 543065 270543 543099
rect 259377 542997 259411 543031
rect 265173 542997 265207 543031
rect 220737 542929 220771 542963
rect 263701 542929 263735 542963
rect 215769 542861 215803 542895
rect 241529 542861 241563 542895
rect 241713 542861 241747 542895
rect 263517 542861 263551 542895
rect 265173 542861 265207 542895
rect 270509 542861 270543 542895
rect 280077 543133 280111 543167
rect 273085 542861 273119 542895
rect 275293 543065 275327 543099
rect 280077 542929 280111 542963
rect 284861 543201 284895 543235
rect 280169 542929 280203 542963
rect 284769 542997 284803 543031
rect 275293 542861 275327 542895
rect 284769 542861 284803 542895
rect 318809 543201 318843 543235
rect 292405 543133 292439 543167
rect 289829 543065 289863 543099
rect 284861 542861 284895 542895
rect 289737 542997 289771 543031
rect 289737 542861 289771 542895
rect 289829 542861 289863 542895
rect 299397 543133 299431 543167
rect 292405 542861 292439 542895
rect 294613 543065 294647 543099
rect 299397 542929 299431 542963
rect 299489 543133 299523 543167
rect 294613 542861 294647 542895
rect 299489 542861 299523 542895
rect 308873 543133 308907 543167
rect 311725 543133 311759 543167
rect 309149 543065 309183 543099
rect 309057 542861 309091 542895
rect 309149 542861 309183 542895
rect 318717 543133 318751 543167
rect 311725 542861 311759 542895
rect 313933 543065 313967 543099
rect 318717 542929 318751 542963
rect 323501 543201 323535 543235
rect 318809 542929 318843 542963
rect 323409 542997 323443 543031
rect 313933 542861 313967 542895
rect 323409 542861 323443 542895
rect 424977 543201 425011 543235
rect 346593 543133 346627 543167
rect 323501 542861 323535 542895
rect 327089 543065 327123 543099
rect 328469 542997 328503 543031
rect 328561 542929 328595 542963
rect 355977 543133 356011 543167
rect 424977 543065 425011 543099
rect 355977 542997 356011 543031
rect 365821 542997 365855 543031
rect 346593 542929 346627 542963
rect 327089 542861 327123 542895
rect 365821 542861 365855 542895
rect 370053 542997 370087 543031
rect 389097 542997 389131 543031
rect 389189 542997 389223 543031
rect 398757 542997 398791 543031
rect 398941 542997 398975 543031
rect 369777 542861 369811 542895
rect 128369 542793 128403 542827
rect 355425 243185 355459 243219
rect 183569 243049 183603 243083
rect 48329 242913 48363 242947
rect 48329 242777 48363 242811
rect 57897 242913 57931 242947
rect 67649 242913 67683 242947
rect 67649 242777 67683 242811
rect 77217 242913 77251 242947
rect 57897 242709 57931 242743
rect 60657 242709 60691 242743
rect 60749 242709 60783 242743
rect 77217 242709 77251 242743
rect 82093 242913 82127 242947
rect 82093 242709 82127 242743
rect 86877 242913 86911 242947
rect 132509 242913 132543 242947
rect 86877 242505 86911 242539
rect 89637 242777 89671 242811
rect 89637 242505 89671 242539
rect 94513 242777 94547 242811
rect 113189 242777 113223 242811
rect 94513 242505 94547 242539
rect 103529 242505 103563 242539
rect 103529 241757 103563 241791
rect 113097 242505 113131 242539
rect 113097 241757 113131 241791
rect 122757 242777 122791 242811
rect 132509 242777 132543 242811
rect 142261 242913 142295 242947
rect 171793 242845 171827 242879
rect 113189 241689 113223 241723
rect 122665 241689 122699 241723
rect 142169 242505 142203 242539
rect 142261 242505 142295 242539
rect 152473 242777 152507 242811
rect 162133 242777 162167 242811
rect 152473 242505 152507 242539
rect 152565 242505 152599 242539
rect 142169 241485 142203 241519
rect 162133 242301 162167 242335
rect 178785 242845 178819 242879
rect 183477 242777 183511 242811
rect 183293 242709 183327 242743
rect 178785 242641 178819 242675
rect 190653 243049 190687 243083
rect 184213 242981 184247 243015
rect 273177 242913 273211 242947
rect 190653 242845 190687 242879
rect 200773 242845 200807 242879
rect 184213 242709 184247 242743
rect 183569 242641 183603 242675
rect 200773 242641 200807 242675
rect 220093 242777 220127 242811
rect 171793 242301 171827 242335
rect 261493 242777 261527 242811
rect 238493 242301 238527 242335
rect 220093 242097 220127 242131
rect 238401 242165 238435 242199
rect 238493 242165 238527 242199
rect 267657 242777 267691 242811
rect 273177 242777 273211 242811
rect 342913 242913 342947 242947
rect 271337 242709 271371 242743
rect 267657 242573 267691 242607
rect 268301 242573 268335 242607
rect 261493 241893 261527 241927
rect 238401 241553 238435 241587
rect 238677 241757 238711 241791
rect 152565 241485 152599 241519
rect 238677 241485 238711 241519
rect 268301 241485 268335 241519
rect 268393 242029 268427 242063
rect 276765 242709 276799 242743
rect 341993 242641 342027 242675
rect 347697 242913 347731 242947
rect 345949 242845 345983 242879
rect 342913 242505 342947 242539
rect 345673 242505 345707 242539
rect 341993 242437 342027 242471
rect 276765 242233 276799 242267
rect 345673 242165 345707 242199
rect 350825 242913 350859 242947
rect 350181 242845 350215 242879
rect 350365 242845 350399 242879
rect 350457 242777 350491 242811
rect 350365 242709 350399 242743
rect 350549 242641 350583 242675
rect 347697 242573 347731 242607
rect 345949 241961 345983 241995
rect 350549 242505 350583 242539
rect 344017 241893 344051 241927
rect 271337 241621 271371 241655
rect 274373 241825 274407 241859
rect 344109 241893 344143 241927
rect 344109 241689 344143 241723
rect 344201 241689 344235 241723
rect 350549 241689 350583 241723
rect 350641 242505 350675 242539
rect 274373 241553 274407 241587
rect 350825 242573 350859 242607
rect 355241 242437 355275 242471
rect 369961 242913 369995 242947
rect 364625 242777 364659 242811
rect 367201 242709 367235 242743
rect 367293 242641 367327 242675
rect 367201 242573 367235 242607
rect 367385 242573 367419 242607
rect 364625 242437 364659 242471
rect 367201 242437 367235 242471
rect 350917 241893 350951 241927
rect 355149 241893 355183 241927
rect 355241 241893 355275 241927
rect 355333 242233 355367 242267
rect 355425 242233 355459 242267
rect 268393 241485 268427 241519
rect 350549 241485 350583 241519
rect 353309 241689 353343 241723
rect 353309 241485 353343 241519
rect 355333 241757 355367 241791
rect 369225 242437 369259 242471
rect 369225 242301 369259 242335
rect 367201 241553 367235 241587
rect 418169 242913 418203 242947
rect 379529 242845 379563 242879
rect 370053 242777 370087 242811
rect 379529 242709 379563 242743
rect 370053 242301 370087 242335
rect 379621 242641 379655 242675
rect 414029 242505 414063 242539
rect 412741 242437 412775 242471
rect 412925 242437 412959 242471
rect 394249 242369 394283 242403
rect 379529 242165 379563 242199
rect 379621 242165 379655 242199
rect 379529 241757 379563 241791
rect 393973 242097 394007 242131
rect 414029 242301 414063 242335
rect 450001 242777 450035 242811
rect 422953 242573 422987 242607
rect 431877 242573 431911 242607
rect 422953 242437 422987 242471
rect 431969 242437 432003 242471
rect 418169 242301 418203 242335
rect 412833 242233 412867 242267
rect 395537 242165 395571 242199
rect 412833 242097 412867 242131
rect 418261 242233 418295 242267
rect 418261 242097 418295 242131
rect 418353 242233 418387 242267
rect 395537 241825 395571 241859
rect 394249 241757 394283 241791
rect 393973 241621 394007 241655
rect 369961 241485 369995 241519
rect 418353 241485 418387 241519
rect 419549 242097 419583 242131
rect 443101 242097 443135 242131
rect 450001 242097 450035 242131
rect 442641 242029 442675 242063
rect 419549 241485 419583 241519
rect 198289 241417 198323 241451
rect 194977 235909 195011 235943
rect 169953 227001 169987 227035
rect 154865 224961 154899 224995
rect 154865 222173 154899 222207
rect 156153 224961 156187 224995
rect 156153 222173 156187 222207
rect 303813 241417 303847 241451
rect 355149 241417 355183 241451
rect 423229 241417 423263 241451
rect 198289 231829 198323 231863
rect 237665 239377 237699 239411
rect 237665 231829 237699 231863
rect 423229 239241 423263 239275
rect 303813 231829 303847 231863
rect 194977 226321 195011 226355
rect 403541 231761 403575 231795
rect 278881 225029 278915 225063
rect 169953 222173 169987 222207
rect 191941 224961 191975 224995
rect 191941 222173 191975 222207
rect 223865 222173 223899 222207
rect 223865 220813 223899 220847
rect 225153 222173 225187 222207
rect 278881 222173 278915 222207
rect 403541 222173 403575 222207
rect 423229 224961 423263 224995
rect 423229 222173 423263 222207
rect 225153 220813 225187 220847
rect 424701 222105 424735 222139
rect 216965 219385 216999 219419
rect 179521 215373 179555 215407
rect 178233 215237 178267 215271
rect 178233 212517 178267 212551
rect 179521 212517 179555 212551
rect 216965 211089 216999 211123
rect 218253 219385 218287 219419
rect 214021 209797 214055 209831
rect 265081 215373 265115 215407
rect 263793 215237 263827 215271
rect 263793 212517 263827 212551
rect 265081 212517 265115 212551
rect 270601 215373 270635 215407
rect 270601 212517 270635 212551
rect 272073 215237 272107 215271
rect 272073 212517 272107 212551
rect 424701 212517 424735 212551
rect 218253 205581 218287 205615
rect 384681 211089 384715 211123
rect 384681 205581 384715 205615
rect 423229 205649 423263 205683
rect 214021 202861 214055 202895
rect 423229 202861 423263 202895
rect 423229 202725 423263 202759
rect 150725 201433 150759 201467
rect 218253 201433 218287 201467
rect 218253 193137 218287 193171
rect 248153 201433 248187 201467
rect 423229 193273 423263 193307
rect 248153 191845 248187 191879
rect 150725 183549 150759 183583
rect 196265 188989 196299 189023
rect 190745 183481 190779 183515
rect 150725 182121 150759 182155
rect 190745 173893 190779 173927
rect 192033 183413 192067 183447
rect 423137 186337 423171 186371
rect 423137 183549 423171 183583
rect 219541 183481 219575 183515
rect 218253 183413 218287 183447
rect 218253 180013 218287 180047
rect 219541 180013 219575 180047
rect 238493 182121 238527 182155
rect 196265 179401 196299 179435
rect 192033 173893 192067 173927
rect 194793 179333 194827 179367
rect 150725 173689 150759 173723
rect 384589 182121 384623 182155
rect 384589 176613 384623 176647
rect 424517 182121 424551 182155
rect 424517 173825 424551 173859
rect 238493 172533 238527 172567
rect 423229 172465 423263 172499
rect 194793 169745 194827 169779
rect 219541 171037 219575 171071
rect 194793 168317 194827 168351
rect 156153 164169 156187 164203
rect 174001 164169 174035 164203
rect 194793 158729 194827 158763
rect 206017 162809 206051 162843
rect 174001 157301 174035 157335
rect 198289 158661 198323 158695
rect 156153 154581 156187 154615
rect 194701 150365 194735 150399
rect 174001 144857 174035 144891
rect 162961 143497 162995 143531
rect 150817 140709 150851 140743
rect 150817 131121 150851 131155
rect 152197 140709 152231 140743
rect 162961 137921 162995 137955
rect 174001 137921 174035 137955
rect 189273 143497 189307 143531
rect 219541 162401 219575 162435
rect 236285 164169 236319 164203
rect 206017 157301 206051 157335
rect 216781 161381 216815 161415
rect 216781 151793 216815 151827
rect 219541 160021 219575 160055
rect 236285 157233 236319 157267
rect 237573 164169 237607 164203
rect 252753 164169 252787 164203
rect 237573 157233 237607 157267
rect 248337 162809 248371 162843
rect 252753 157301 252787 157335
rect 284401 164169 284435 164203
rect 284401 157301 284435 157335
rect 307953 164169 307987 164203
rect 307953 157301 307987 157335
rect 346225 164169 346259 164203
rect 346225 157301 346259 157335
rect 357265 164169 357299 164203
rect 423229 162877 423263 162911
rect 357265 157301 357299 157335
rect 374285 162809 374319 162843
rect 248337 153221 248371 153255
rect 263793 154513 263827 154547
rect 219541 150433 219575 150467
rect 198289 149073 198323 149107
rect 379069 162809 379103 162843
rect 379069 157301 379103 157335
rect 384589 162809 384623 162843
rect 374285 153221 374319 153255
rect 424701 162809 424735 162843
rect 424701 157301 424735 157335
rect 384589 153221 384623 153255
rect 263793 148325 263827 148359
rect 423229 153153 423263 153187
rect 252753 144857 252787 144891
rect 194701 140777 194735 140811
rect 238677 143497 238711 143531
rect 189273 133909 189307 133943
rect 216781 135201 216815 135235
rect 152197 131121 152231 131155
rect 153393 133841 153427 133875
rect 153393 124185 153427 124219
rect 156153 133841 156187 133875
rect 156153 124185 156187 124219
rect 168849 133841 168883 133875
rect 192033 132413 192067 132447
rect 168849 124185 168883 124219
rect 174001 125545 174035 125579
rect 162961 124117 162995 124151
rect 152013 121397 152047 121431
rect 150725 116297 150759 116331
rect 174001 118609 174035 118643
rect 178233 125545 178267 125579
rect 216781 129693 216815 129727
rect 234813 133841 234847 133875
rect 248337 143497 248371 143531
rect 284401 144857 284435 144891
rect 252753 137921 252787 137955
rect 263793 142069 263827 142103
rect 248337 133909 248371 133943
rect 238677 125613 238711 125647
rect 245761 133841 245795 133875
rect 234813 124253 234847 124287
rect 284401 137921 284435 137955
rect 307953 144857 307987 144891
rect 307953 137921 307987 137955
rect 346225 144857 346259 144891
rect 346225 137921 346259 137955
rect 357265 144857 357299 144891
rect 423229 143565 423263 143599
rect 357265 137921 357299 137955
rect 374285 143497 374319 143531
rect 424701 143497 424735 143531
rect 374285 133909 374319 133943
rect 379161 142069 379195 142103
rect 263793 132481 263827 132515
rect 424701 137921 424735 137955
rect 379161 132481 379195 132515
rect 384681 133841 384715 133875
rect 379161 132345 379195 132379
rect 245761 124185 245795 124219
rect 252753 125545 252787 125579
rect 178233 115957 178267 115991
rect 189273 124117 189307 124151
rect 192033 124117 192067 124151
rect 234813 124117 234847 124151
rect 162961 114529 162995 114563
rect 189273 114529 189307 114563
rect 234813 114529 234847 114563
rect 238585 124117 238619 124151
rect 238585 114529 238619 114563
rect 248337 124117 248371 124151
rect 284401 125545 284435 125579
rect 252753 118609 252787 118643
rect 263793 122757 263827 122791
rect 248337 114529 248371 114563
rect 168849 114461 168883 114495
rect 152013 111809 152047 111843
rect 153301 114393 153335 114427
rect 207029 114461 207063 114495
rect 191941 113237 191975 113271
rect 191941 111809 191975 111843
rect 168849 106233 168883 106267
rect 174001 106233 174035 106267
rect 153301 104873 153335 104907
rect 154773 106165 154807 106199
rect 150725 103513 150759 103547
rect 152013 102085 152047 102119
rect 154773 96713 154807 96747
rect 168849 104805 168883 104839
rect 174001 99297 174035 99331
rect 178233 106233 178267 106267
rect 190653 106233 190687 106267
rect 263793 114257 263827 114291
rect 264989 122757 265023 122791
rect 284401 118609 284435 118643
rect 307953 125545 307987 125579
rect 307953 118609 307987 118643
rect 346225 125545 346259 125579
rect 346225 118609 346259 118643
rect 357265 125545 357299 125579
rect 357265 118609 357299 118643
rect 374285 124117 374319 124151
rect 384681 127789 384715 127823
rect 424701 133841 424735 133875
rect 424701 124253 424735 124287
rect 379161 122825 379195 122859
rect 424701 124117 424735 124151
rect 374285 114529 374319 114563
rect 423229 122757 423263 122791
rect 264989 113169 265023 113203
rect 384589 114393 384623 114427
rect 245761 109701 245795 109735
rect 207029 104873 207063 104907
rect 208409 106301 208443 106335
rect 208409 104873 208443 104907
rect 245761 104873 245795 104907
rect 252753 106233 252787 106267
rect 223773 104805 223807 104839
rect 190653 101337 190687 101371
rect 206017 103445 206051 103479
rect 178233 96645 178267 96679
rect 168849 95217 168883 95251
rect 152013 92497 152047 92531
rect 188997 95149 189031 95183
rect 169769 86921 169803 86955
rect 162961 85493 162995 85527
rect 152013 82773 152047 82807
rect 152013 73185 152047 73219
rect 154773 77197 154807 77231
rect 150725 70261 150759 70295
rect 169769 77265 169803 77299
rect 174001 86921 174035 86955
rect 174001 77265 174035 77299
rect 178233 86921 178267 86955
rect 208409 103445 208443 103479
rect 223773 95217 223807 95251
rect 238677 104805 238711 104839
rect 238677 95217 238711 95251
rect 248337 104805 248371 104839
rect 284401 106233 284435 106267
rect 252753 99297 252787 99331
rect 263793 104805 263827 104839
rect 263793 96849 263827 96883
rect 270509 103445 270543 103479
rect 248337 95217 248371 95251
rect 208409 95081 208443 95115
rect 211353 95149 211387 95183
rect 206017 93857 206051 93891
rect 206017 86989 206051 87023
rect 188997 85561 189031 85595
rect 190653 86921 190687 86955
rect 190653 80665 190687 80699
rect 191941 86921 191975 86955
rect 178233 77265 178267 77299
rect 162961 75905 162995 75939
rect 206017 85561 206051 85595
rect 211353 85561 211387 85595
rect 216873 95149 216907 95183
rect 216873 85561 216907 85595
rect 218345 95149 218379 95183
rect 218345 85561 218379 85595
rect 219633 95149 219667 95183
rect 270509 93857 270543 93891
rect 272073 103445 272107 103479
rect 284401 99297 284435 99331
rect 307953 106233 307987 106267
rect 307953 99297 307987 99331
rect 346225 106233 346259 106267
rect 346225 99297 346259 99331
rect 357265 106233 357299 106267
rect 424701 114529 424735 114563
rect 423229 113169 423263 113203
rect 384589 104873 384623 104907
rect 423045 109701 423079 109735
rect 423045 104873 423079 104907
rect 424701 107049 424735 107083
rect 357265 99297 357299 99331
rect 374285 104805 374319 104839
rect 374285 95217 374319 95251
rect 379161 100045 379195 100079
rect 272073 93857 272107 93891
rect 226625 93789 226659 93823
rect 226625 92497 226659 92531
rect 219633 85561 219667 85595
rect 245761 90389 245795 90423
rect 223773 85493 223807 85527
rect 191941 75905 191975 75939
rect 194885 84133 194919 84167
rect 194885 74545 194919 74579
rect 207029 84133 207063 84167
rect 154773 67609 154807 67643
rect 190653 70465 190687 70499
rect 190653 66249 190687 66283
rect 208501 84133 208535 84167
rect 238677 85493 238711 85527
rect 223773 74545 223807 74579
rect 226533 82773 226567 82807
rect 208501 66317 208535 66351
rect 211261 74477 211295 74511
rect 207029 66249 207063 66283
rect 150725 64821 150759 64855
rect 162869 66181 162903 66215
rect 154773 57885 154807 57919
rect 162869 56593 162903 56627
rect 168481 66181 168515 66215
rect 211261 64957 211295 64991
rect 219541 66181 219575 66215
rect 189181 64821 189215 64855
rect 168481 56593 168515 56627
rect 174001 57885 174035 57919
rect 154773 48365 154807 48399
rect 174001 48297 174035 48331
rect 178233 57885 178267 57919
rect 178233 48297 178267 48331
rect 154773 48229 154807 48263
rect 207121 64821 207155 64855
rect 190653 64617 190687 64651
rect 190653 56593 190687 56627
rect 198197 63461 198231 63495
rect 192033 55301 192067 55335
rect 192033 53805 192067 53839
rect 194701 55233 194735 55267
rect 194701 53805 194735 53839
rect 207121 56321 207155 56355
rect 208501 64821 208535 64855
rect 208501 55233 208535 55267
rect 211353 64821 211387 64855
rect 211353 55233 211387 55267
rect 218253 64821 218287 64855
rect 198197 53805 198231 53839
rect 216965 55165 216999 55199
rect 189181 46937 189215 46971
rect 211261 47277 211295 47311
rect 154773 43673 154807 43707
rect 168573 46869 168607 46903
rect 168573 37281 168607 37315
rect 169861 46869 169895 46903
rect 169861 37281 169895 37315
rect 207121 46869 207155 46903
rect 211261 45577 211295 45611
rect 214113 46869 214147 46903
rect 207121 37281 207155 37315
rect 208593 42041 208627 42075
rect 190653 37213 190687 37247
rect 174001 33813 174035 33847
rect 174001 28985 174035 29019
rect 190653 27693 190687 27727
rect 207213 37145 207247 37179
rect 218253 46937 218287 46971
rect 223681 64821 223715 64855
rect 223681 55233 223715 55267
rect 424701 99297 424735 99331
rect 379161 89369 379195 89403
rect 245761 83181 245795 83215
rect 247049 86921 247083 86955
rect 252753 86921 252787 86955
rect 247049 77265 247083 77299
rect 248337 85493 248371 85527
rect 238677 75905 238711 75939
rect 252753 77265 252787 77299
rect 258089 86921 258123 86955
rect 284401 86921 284435 86955
rect 258089 77265 258123 77299
rect 270509 85493 270543 85527
rect 248337 75905 248371 75939
rect 270509 75905 270543 75939
rect 272073 85493 272107 85527
rect 284401 77265 284435 77299
rect 307953 86921 307987 86955
rect 307953 77265 307987 77299
rect 346225 86921 346259 86955
rect 346225 77265 346259 77299
rect 357265 86921 357299 86955
rect 424701 86921 424735 86955
rect 357265 77265 357299 77299
rect 374285 85493 374319 85527
rect 272073 75905 272107 75939
rect 303905 77197 303939 77231
rect 246037 74477 246071 74511
rect 226533 55233 226567 55267
rect 238677 66181 238711 66215
rect 303905 70193 303939 70227
rect 357265 77129 357299 77163
rect 252753 67677 252787 67711
rect 424701 77265 424735 77299
rect 374285 75905 374319 75939
rect 357265 67609 357299 67643
rect 384681 75837 384715 75871
rect 252753 66249 252787 66283
rect 384681 66249 384715 66283
rect 424701 67541 424735 67575
rect 246037 64889 246071 64923
rect 248337 66181 248371 66215
rect 263701 66181 263735 66215
rect 248337 56593 248371 56627
rect 258181 57885 258215 57919
rect 238677 48297 238711 48331
rect 258181 48297 258215 48331
rect 265081 66181 265115 66215
rect 265081 60673 265115 60707
rect 374285 66181 374319 66215
rect 307861 57885 307895 57919
rect 263701 48297 263735 48331
rect 270601 51153 270635 51187
rect 270601 48297 270635 48331
rect 271889 51085 271923 51119
rect 271889 48297 271923 48331
rect 307861 48297 307895 48331
rect 357265 57885 357299 57919
rect 379161 66181 379195 66215
rect 424701 57953 424735 57987
rect 379161 56661 379195 56695
rect 374285 56593 374319 56627
rect 357265 48297 357299 48331
rect 379161 56525 379195 56559
rect 219541 46937 219575 46971
rect 234813 48229 234847 48263
rect 216965 45577 216999 45611
rect 219449 45509 219483 45543
rect 219449 37213 219483 37247
rect 222485 42041 222519 42075
rect 214113 32385 214147 32419
rect 208593 28985 208627 29019
rect 222485 28985 222519 29019
rect 223773 42041 223807 42075
rect 284493 48229 284527 48263
rect 234813 38641 234847 38675
rect 238585 46869 238619 46903
rect 248337 46869 248371 46903
rect 238585 37281 238619 37315
rect 245761 45509 245795 45543
rect 223773 28985 223807 29019
rect 238677 28985 238711 29019
rect 207213 27693 207247 27727
rect 238677 27693 238711 27727
rect 247417 45509 247451 45543
rect 379161 46937 379195 46971
rect 424701 48229 424735 48263
rect 284493 41361 284527 41395
rect 374285 46869 374319 46903
rect 248337 37281 248371 37315
rect 284401 38573 284435 38607
rect 247417 37213 247451 37247
rect 270601 31841 270635 31875
rect 191941 27625 191975 27659
rect 245761 27625 245795 27659
rect 247417 31297 247451 31331
rect 247417 27625 247451 27659
rect 270601 27625 270635 27659
rect 273361 31841 273395 31875
rect 284401 28985 284435 29019
rect 307953 38573 307987 38607
rect 357265 38573 357299 38607
rect 424701 38641 424735 38675
rect 374285 37281 374319 37315
rect 403817 38573 403851 38607
rect 357265 31705 357299 31739
rect 307953 28985 307987 29019
rect 403817 28985 403851 29019
rect 273361 27625 273395 27659
rect 394065 28917 394099 28951
rect 174001 27557 174035 27591
rect 174001 22049 174035 22083
rect 179521 27557 179555 27591
rect 191941 26265 191975 26299
rect 207121 27557 207155 27591
rect 179521 17969 179555 18003
rect 189181 26197 189215 26231
rect 154865 17901 154899 17935
rect 194701 26197 194735 26231
rect 189181 16609 189215 16643
rect 191941 21369 191975 21403
rect 154865 12393 154899 12427
rect 211353 27557 211387 27591
rect 211353 19329 211387 19363
rect 223681 27557 223715 27591
rect 207121 17969 207155 18003
rect 194701 16609 194735 16643
rect 191941 9673 191975 9707
rect 223681 9673 223715 9707
rect 238585 27557 238619 27591
rect 252753 27557 252787 27591
rect 245853 27217 245887 27251
rect 245853 19329 245887 19363
rect 238585 9673 238619 9707
rect 247969 19261 248003 19295
rect 252753 17969 252787 18003
rect 264989 27557 265023 27591
rect 346225 27557 346259 27591
rect 346225 22049 346259 22083
rect 374285 27557 374319 27591
rect 264989 17969 265023 18003
rect 270509 19329 270543 19363
rect 247969 9673 248003 9707
rect 384589 27557 384623 27591
rect 379253 27489 379287 27523
rect 379253 22049 379287 22083
rect 374285 17969 374319 18003
rect 394065 19329 394099 19363
rect 384589 17969 384623 18003
rect 270509 9673 270543 9707
rect 374193 12529 374227 12563
rect 374193 9673 374227 9707
rect 423321 8109 423355 8143
rect 113189 5661 113223 5695
rect 80161 5525 80195 5559
rect 55229 5321 55263 5355
rect 55229 5185 55263 5219
rect 55229 4573 55263 4607
rect 55321 4437 55355 4471
rect 64797 5321 64831 5355
rect 74549 5321 74583 5355
rect 64797 5185 64831 5219
rect 64797 4573 64831 4607
rect 74549 5185 74583 5219
rect 64705 4437 64739 4471
rect 74641 4233 74675 4267
rect 84117 5525 84151 5559
rect 84117 5321 84151 5355
rect 93869 5525 93903 5559
rect 80161 4233 80195 4267
rect 84117 5185 84151 5219
rect 93869 5185 93903 5219
rect 103437 5525 103471 5559
rect 103437 5185 103471 5219
rect 113189 5185 113223 5219
rect 122757 5661 122791 5695
rect 122757 5185 122791 5219
rect 132509 5661 132543 5695
rect 132509 5185 132543 5219
rect 142077 5661 142111 5695
rect 183569 5457 183603 5491
rect 422861 5457 422895 5491
rect 422953 5457 422987 5491
rect 181453 5389 181487 5423
rect 152289 5321 152323 5355
rect 162225 5321 162259 5355
rect 152105 5253 152139 5287
rect 160845 5253 160879 5287
rect 142077 5185 142111 5219
rect 74549 4165 74583 4199
rect 148977 5117 149011 5151
rect 181453 5253 181487 5287
rect 162225 5185 162259 5219
rect 160845 5049 160879 5083
rect 148977 4981 149011 5015
rect 191113 5389 191147 5423
rect 183569 4709 183603 4743
rect 188353 4709 188387 4743
rect 422217 5117 422251 5151
rect 403541 5049 403575 5083
rect 400229 4777 400263 4811
rect 400413 4709 400447 4743
rect 191113 4641 191147 4675
rect 412557 5049 412591 5083
rect 403541 4505 403575 4539
rect 403633 4573 403667 4607
rect 188353 4369 188387 4403
rect 393881 4369 393915 4403
rect 83749 4165 83783 4199
rect 388361 4301 388395 4335
rect 393881 4233 393915 4267
rect 403633 4233 403667 4267
rect 412465 4573 412499 4607
rect 412557 4505 412591 4539
rect 423321 5117 423355 5151
rect 424057 5389 424091 5423
rect 432429 5389 432463 5423
rect 422953 4845 422987 4879
rect 423137 4981 423171 5015
rect 423137 4777 423171 4811
rect 423229 4981 423263 5015
rect 423321 4777 423355 4811
rect 422769 4641 422803 4675
rect 422861 4709 422895 4743
rect 423045 4573 423079 4607
rect 422217 4505 422251 4539
rect 441537 5321 441571 5355
rect 432521 5185 432555 5219
rect 432889 5185 432923 5219
rect 437121 5185 437155 5219
rect 426449 5117 426483 5151
rect 426449 4505 426483 4539
rect 427829 4777 427863 4811
rect 424057 4437 424091 4471
rect 440709 5117 440743 5151
rect 437121 4981 437155 5015
rect 438317 4981 438351 5015
rect 440709 4913 440743 4947
rect 432797 4845 432831 4879
rect 438317 4845 438351 4879
rect 446505 5185 446539 5219
rect 441629 5049 441663 5083
rect 441537 4845 441571 4879
rect 446505 4913 446539 4947
rect 446597 4913 446631 4947
rect 441905 4845 441939 4879
rect 432613 4777 432647 4811
rect 446597 4777 446631 4811
rect 432705 4709 432739 4743
rect 427829 4369 427863 4403
rect 412465 4233 412499 4267
rect 388361 4165 388395 4199
rect 191205 4097 191239 4131
rect 191021 3757 191055 3791
rect 181361 3621 181395 3655
rect 181361 3281 181395 3315
rect 186237 3553 186271 3587
rect 191205 3621 191239 3655
rect 196725 4097 196759 4131
rect 268393 4029 268427 4063
rect 196725 3621 196759 3655
rect 209329 3961 209363 3995
rect 209329 3621 209363 3655
rect 216505 3961 216539 3995
rect 256893 3825 256927 3859
rect 239505 3757 239539 3791
rect 235825 3689 235859 3723
rect 216505 3621 216539 3655
rect 225245 3621 225279 3655
rect 191021 3349 191055 3383
rect 191113 3553 191147 3587
rect 186237 3281 186271 3315
rect 191113 3213 191147 3247
rect 200773 3553 200807 3587
rect 208777 3553 208811 3587
rect 208777 3281 208811 3315
rect 220093 3553 220127 3587
rect 226349 3621 226383 3655
rect 226349 3485 226383 3519
rect 231869 3621 231903 3655
rect 231869 3485 231903 3519
rect 231961 3485 231995 3519
rect 225245 3349 225279 3383
rect 235733 3485 235767 3519
rect 235825 3485 235859 3519
rect 236469 3485 236503 3519
rect 239505 3485 239539 3519
rect 244289 3621 244323 3655
rect 231961 3349 231995 3383
rect 232053 3349 232087 3383
rect 220093 3281 220127 3315
rect 220185 3281 220219 3315
rect 200773 3213 200807 3247
rect 220185 3145 220219 3179
rect 263609 3757 263643 3791
rect 342729 4029 342763 4063
rect 268393 3621 268427 3655
rect 268485 3757 268519 3791
rect 268485 3621 268519 3655
rect 263609 3553 263643 3587
rect 345765 4029 345799 4063
rect 345765 3621 345799 3655
rect 342729 3349 342763 3383
rect 345581 3553 345615 3587
rect 244289 3213 244323 3247
rect 249073 3281 249107 3315
rect 253765 3281 253799 3315
rect 254777 3281 254811 3315
rect 256893 3281 256927 3315
rect 232053 3077 232087 3111
rect 232145 3077 232179 3111
rect 127633 2873 127667 2907
rect 232145 2873 232179 2907
rect 127449 2805 127483 2839
rect 249073 2805 249107 2839
rect 250545 3213 250579 3247
rect 345581 3077 345615 3111
rect 350457 3485 350491 3519
rect 350457 3077 350491 3111
rect 386429 2941 386463 2975
rect 250545 2737 250579 2771
rect 290749 2805 290783 2839
rect 386429 2737 386463 2771
rect 395997 2873 396031 2907
rect 395997 2737 396031 2771
rect 290749 561 290783 595
rect 374009 2669 374043 2703
rect 374009 561 374043 595
<< metal1 >>
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 318794 700992 318800 701004
rect 154172 700964 318800 700992
rect 154172 700952 154178 700964
rect 318794 700952 318800 700964
rect 318852 700952 318858 701004
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 316034 700924 316040 700936
rect 137888 700896 316040 700924
rect 137888 700884 137894 700896
rect 316034 700884 316040 700896
rect 316092 700884 316098 700936
rect 278682 700816 278688 700868
rect 278740 700856 278746 700868
rect 462314 700856 462320 700868
rect 278740 700828 462320 700856
rect 278740 700816 278746 700828
rect 462314 700816 462320 700828
rect 462372 700816 462378 700868
rect 281442 700748 281448 700800
rect 281500 700788 281506 700800
rect 478506 700788 478512 700800
rect 281500 700760 478512 700788
rect 281500 700748 281506 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 105446 700680 105452 700732
rect 105504 700720 105510 700732
rect 321554 700720 321560 700732
rect 105504 700692 321560 700720
rect 105504 700680 105510 700692
rect 321554 700680 321560 700692
rect 321612 700680 321618 700732
rect 89162 700612 89168 700664
rect 89220 700652 89226 700664
rect 327074 700652 327080 700664
rect 89220 700624 327080 700652
rect 89220 700612 89226 700624
rect 327074 700612 327080 700624
rect 327132 700612 327138 700664
rect 72970 700544 72976 700596
rect 73028 700584 73034 700596
rect 324314 700584 324320 700596
rect 73028 700556 324320 700584
rect 73028 700544 73034 700556
rect 324314 700544 324320 700556
rect 324372 700544 324378 700596
rect 270402 700476 270408 700528
rect 270460 700516 270466 700528
rect 527174 700516 527180 700528
rect 270460 700488 527180 700516
rect 270460 700476 270466 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 273162 700408 273168 700460
rect 273220 700448 273226 700460
rect 543458 700448 543464 700460
rect 273220 700420 543464 700448
rect 273220 700408 273226 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 328454 700380 328460 700392
rect 40552 700352 328460 700380
rect 40552 700340 40558 700352
rect 328454 700340 328460 700352
rect 328512 700340 328518 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 333974 700312 333980 700324
rect 24360 700284 333980 700312
rect 24360 700272 24366 700284
rect 333974 700272 333980 700284
rect 334032 700272 334038 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 313274 700244 313280 700256
rect 170364 700216 313280 700244
rect 170364 700204 170370 700216
rect 313274 700204 313280 700216
rect 313332 700204 313338 700256
rect 288342 700136 288348 700188
rect 288400 700176 288406 700188
rect 413646 700176 413652 700188
rect 288400 700148 413652 700176
rect 288400 700136 288406 700148
rect 413646 700136 413652 700148
rect 413704 700136 413710 700188
rect 286962 700068 286968 700120
rect 287020 700108 287026 700120
rect 397454 700108 397460 700120
rect 287020 700080 397460 700108
rect 287020 700068 287026 700080
rect 397454 700068 397460 700080
rect 397512 700068 397518 700120
rect 202782 700000 202788 700052
rect 202840 700040 202846 700052
rect 307754 700040 307760 700052
rect 202840 700012 307760 700040
rect 202840 700000 202846 700012
rect 307754 700000 307760 700012
rect 307812 700000 307818 700052
rect 218974 699932 218980 699984
rect 219032 699972 219038 699984
rect 310514 699972 310520 699984
rect 219032 699944 310520 699972
rect 219032 699932 219038 699944
rect 310514 699932 310520 699944
rect 310572 699932 310578 699984
rect 296622 699864 296628 699916
rect 296680 699904 296686 699916
rect 348786 699904 348792 699916
rect 296680 699876 348792 699904
rect 296680 699864 296686 699876
rect 348786 699864 348792 699876
rect 348844 699864 348850 699916
rect 293862 699796 293868 699848
rect 293920 699836 293926 699848
rect 332502 699836 332508 699848
rect 293920 699808 332508 699836
rect 293920 699796 293926 699808
rect 332502 699796 332508 699808
rect 332560 699796 332566 699848
rect 267642 699728 267648 699780
rect 267700 699768 267706 699780
rect 300854 699768 300860 699780
rect 267700 699740 300860 699768
rect 267700 699728 267706 699740
rect 300854 699728 300860 699740
rect 300912 699728 300918 699780
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 283834 699660 283840 699712
rect 283892 699700 283898 699712
rect 303614 699700 303620 699712
rect 283892 699672 303620 699700
rect 283892 699660 283898 699672
rect 303614 699660 303620 699672
rect 303672 699660 303678 699712
rect 263502 696940 263508 696992
rect 263560 696980 263566 696992
rect 580166 696980 580172 696992
rect 263560 696952 580172 696980
rect 263560 696940 263566 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 299658 688576 299664 688628
rect 299716 688616 299722 688628
rect 300118 688616 300124 688628
rect 299716 688588 300124 688616
rect 299716 688576 299722 688588
rect 300118 688576 300124 688588
rect 300176 688576 300182 688628
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 299492 685936 301268 685964
rect 266262 685856 266268 685908
rect 266320 685896 266326 685908
rect 299492 685896 299520 685936
rect 266320 685868 299520 685896
rect 301240 685896 301268 685936
rect 429212 685936 429976 685964
rect 429212 685896 429240 685936
rect 301240 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 266320 685856 266326 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299845 684471 299903 684477
rect 299845 684468 299857 684471
rect 299624 684440 299857 684468
rect 299624 684428 299630 684440
rect 299845 684437 299857 684440
rect 299891 684437 299903 684471
rect 299845 684431 299903 684437
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429565 684471 429623 684477
rect 429565 684468 429577 684471
rect 429344 684440 429577 684468
rect 429344 684428 429350 684440
rect 429565 684437 429577 684440
rect 429611 684437 429623 684471
rect 429565 684431 429623 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 336734 681748 336740 681760
rect 3568 681720 336740 681748
rect 3568 681708 3574 681720
rect 336734 681708 336740 681720
rect 336792 681708 336798 681760
rect 364334 676172 364340 676184
rect 364295 676144 364340 676172
rect 364334 676132 364340 676144
rect 364392 676132 364398 676184
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 260742 673480 260748 673532
rect 260800 673520 260806 673532
rect 580166 673520 580172 673532
rect 260800 673492 580172 673520
rect 260800 673480 260806 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 342254 667944 342260 667956
rect 3476 667916 342260 667944
rect 3476 667904 3482 667916
rect 342254 667904 342260 667916
rect 342312 667904 342318 667956
rect 299845 666587 299903 666593
rect 299845 666553 299857 666587
rect 299891 666584 299903 666587
rect 299934 666584 299940 666596
rect 299891 666556 299940 666584
rect 299891 666553 299903 666556
rect 299845 666547 299903 666553
rect 299934 666544 299940 666556
rect 299992 666544 299998 666596
rect 364337 666587 364395 666593
rect 364337 666553 364349 666587
rect 364383 666584 364395 666587
rect 364426 666584 364432 666596
rect 364383 666556 364432 666584
rect 364383 666553 364395 666556
rect 364337 666547 364395 666553
rect 364426 666544 364432 666556
rect 364484 666544 364490 666596
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 339494 652780 339500 652792
rect 3108 652752 339500 652780
rect 3108 652740 3114 652752
rect 339494 652740 339500 652752
rect 339552 652740 339558 652792
rect 255222 650020 255228 650072
rect 255280 650060 255286 650072
rect 580166 650060 580172 650072
rect 255280 650032 580172 650060
rect 255280 650020 255286 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 299658 647232 299664 647284
rect 299716 647272 299722 647284
rect 299750 647272 299756 647284
rect 299716 647244 299756 647272
rect 299716 647232 299722 647244
rect 299750 647232 299756 647244
rect 299808 647232 299814 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 299658 640364 299664 640416
rect 299716 640404 299722 640416
rect 299750 640404 299756 640416
rect 299716 640376 299756 640404
rect 299716 640364 299722 640376
rect 299750 640364 299756 640376
rect 299808 640364 299814 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 257982 638936 257988 638988
rect 258040 638976 258046 638988
rect 580166 638976 580172 638988
rect 258040 638948 580172 638976
rect 258040 638936 258046 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 364334 634788 364340 634840
rect 364392 634828 364398 634840
rect 364518 634828 364524 634840
rect 364392 634800 364524 634828
rect 364392 634788 364398 634800
rect 364518 634788 364524 634800
rect 364576 634788 364582 634840
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 299750 630680 299756 630692
rect 299624 630652 299756 630680
rect 299624 630640 299630 630652
rect 299750 630640 299756 630652
rect 299808 630640 299814 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 252462 626560 252468 626612
rect 252520 626600 252526 626612
rect 580166 626600 580172 626612
rect 252520 626572 580172 626600
rect 252520 626560 252526 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 345014 623812 345020 623824
rect 3476 623784 345020 623812
rect 3476 623772 3482 623784
rect 345014 623772 345020 623784
rect 345072 623772 345078 623824
rect 364334 615476 364340 615528
rect 364392 615516 364398 615528
rect 364518 615516 364524 615528
rect 364392 615488 364524 615516
rect 364392 615476 364398 615488
rect 364518 615476 364524 615488
rect 364576 615476 364582 615528
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 349154 610008 349160 610020
rect 3476 609980 349160 610008
rect 3476 609968 3482 609980
rect 349154 609968 349160 609980
rect 349212 609968 349218 610020
rect 299658 608580 299664 608592
rect 299619 608552 299664 608580
rect 299658 608540 299664 608552
rect 299716 608540 299722 608592
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 246942 603100 246948 603152
rect 247000 603140 247006 603152
rect 580166 603140 580172 603152
rect 247000 603112 580172 603140
rect 247000 603100 247006 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 299661 601715 299719 601721
rect 299661 601681 299673 601715
rect 299707 601712 299719 601715
rect 299842 601712 299848 601724
rect 299707 601684 299848 601712
rect 299707 601681 299719 601684
rect 299661 601675 299719 601681
rect 299842 601672 299848 601684
rect 299900 601672 299906 601724
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 299842 598924 299848 598936
rect 299803 598896 299848 598924
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 364334 596164 364340 596216
rect 364392 596204 364398 596216
rect 364518 596204 364524 596216
rect 364392 596176 364524 596204
rect 364392 596164 364398 596176
rect 364518 596164 364524 596176
rect 364576 596164 364582 596216
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 347774 594844 347780 594856
rect 3292 594816 347780 594844
rect 3292 594804 3298 594816
rect 347774 594804 347780 594816
rect 347832 594804 347838 594856
rect 249702 592016 249708 592068
rect 249760 592056 249766 592068
rect 580166 592056 580172 592068
rect 249760 592028 580172 592056
rect 249760 592016 249766 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 299845 589339 299903 589345
rect 299845 589305 299857 589339
rect 299891 589336 299903 589339
rect 299934 589336 299940 589348
rect 299891 589308 299940 589336
rect 299891 589305 299903 589308
rect 299845 589299 299903 589305
rect 299934 589296 299940 589308
rect 299992 589296 299998 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 364150 589228 364156 589280
rect 364208 589268 364214 589280
rect 364426 589268 364432 589280
rect 364208 589240 364432 589268
rect 364208 589228 364214 589240
rect 364426 589228 364432 589240
rect 364484 589228 364490 589280
rect 493870 589228 493876 589280
rect 493928 589268 493934 589280
rect 494146 589268 494152 589280
rect 493928 589240 494152 589268
rect 493928 589228 493934 589240
rect 494146 589228 494152 589240
rect 494204 589228 494210 589280
rect 299934 582468 299940 582480
rect 299860 582440 299940 582468
rect 299860 582344 299888 582440
rect 299934 582428 299940 582440
rect 299992 582428 299998 582480
rect 429654 582468 429660 582480
rect 429580 582440 429660 582468
rect 429580 582344 429608 582440
rect 429654 582428 429660 582440
rect 429712 582428 429718 582480
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 299842 582292 299848 582344
rect 299900 582292 299906 582344
rect 429562 582292 429568 582344
rect 429620 582292 429626 582344
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 245562 579640 245568 579692
rect 245620 579680 245626 579692
rect 580166 579680 580172 579692
rect 245620 579652 580172 579680
rect 245620 579640 245626 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 3418 567196 3424 567248
rect 3476 567236 3482 567248
rect 351914 567236 351920 567248
rect 3476 567208 351920 567236
rect 3476 567196 3482 567208
rect 351914 567196 351920 567208
rect 351972 567196 351978 567248
rect 299566 563116 299572 563168
rect 299624 563116 299630 563168
rect 429286 563116 429292 563168
rect 429344 563116 429350 563168
rect 559006 563116 559012 563168
rect 559064 563116 559070 563168
rect 299584 563032 299612 563116
rect 429304 563032 429332 563116
rect 559024 563032 559052 563116
rect 299566 562980 299572 563032
rect 299624 562980 299630 563032
rect 429286 562980 429292 563032
rect 429344 562980 429350 563032
rect 559006 562980 559012 563032
rect 559064 562980 559070 563032
rect 299566 560232 299572 560244
rect 299527 560204 299572 560232
rect 299566 560192 299572 560204
rect 299624 560192 299630 560244
rect 559006 560232 559012 560244
rect 558967 560204 559012 560232
rect 559006 560192 559012 560204
rect 559064 560192 559070 560244
rect 240042 556180 240048 556232
rect 240100 556220 240106 556232
rect 580166 556220 580172 556232
rect 240100 556192 580172 556220
rect 240100 556180 240106 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 429194 553432 429200 553444
rect 429155 553404 429200 553432
rect 429194 553392 429200 553404
rect 429252 553392 429258 553444
rect 3418 552100 3424 552152
rect 3476 552140 3482 552152
rect 357434 552140 357440 552152
rect 3476 552112 357440 552140
rect 3476 552100 3482 552112
rect 357434 552100 357440 552112
rect 357492 552100 357498 552152
rect 156414 552032 156420 552084
rect 156472 552072 156478 552084
rect 577498 552072 577504 552084
rect 156472 552044 577504 552072
rect 156472 552032 156478 552044
rect 577498 552032 577504 552044
rect 577556 552032 577562 552084
rect 299569 550647 299627 550653
rect 299569 550613 299581 550647
rect 299615 550644 299627 550647
rect 299658 550644 299664 550656
rect 299615 550616 299664 550644
rect 299615 550613 299627 550616
rect 299569 550607 299627 550613
rect 299658 550604 299664 550616
rect 299716 550604 299722 550656
rect 429194 550644 429200 550656
rect 429155 550616 429200 550644
rect 429194 550604 429200 550616
rect 429252 550604 429258 550656
rect 559009 550647 559067 550653
rect 559009 550613 559021 550647
rect 559055 550644 559067 550647
rect 559098 550644 559104 550656
rect 559055 550616 559104 550644
rect 559055 550613 559067 550616
rect 559009 550607 559067 550613
rect 559098 550604 559104 550616
rect 559156 550604 559162 550656
rect 235902 550128 235908 550180
rect 235960 550168 235966 550180
rect 306374 550168 306380 550180
rect 235960 550140 306380 550168
rect 235960 550128 235966 550140
rect 306374 550128 306380 550140
rect 306432 550128 306438 550180
rect 290918 550060 290924 550112
rect 290976 550100 290982 550112
rect 364334 550100 364340 550112
rect 290976 550072 364340 550100
rect 290976 550060 290982 550072
rect 364334 550060 364340 550072
rect 364392 550060 364398 550112
rect 283098 549992 283104 550044
rect 283156 550032 283162 550044
rect 429194 550032 429200 550044
rect 283156 550004 429200 550032
rect 283156 549992 283162 550004
rect 429194 549992 429200 550004
rect 429252 549992 429258 550044
rect 275370 549924 275376 549976
rect 275428 549964 275434 549976
rect 494054 549964 494060 549976
rect 275428 549936 494060 549964
rect 275428 549924 275434 549936
rect 494054 549924 494060 549936
rect 494112 549924 494118 549976
rect 267642 549856 267648 549908
rect 267700 549896 267706 549908
rect 559098 549896 559104 549908
rect 267700 549868 559104 549896
rect 267700 549856 267706 549868
rect 559098 549856 559104 549868
rect 559156 549856 559162 549908
rect 298646 549244 298652 549296
rect 298704 549284 298710 549296
rect 299566 549284 299572 549296
rect 298704 549256 299572 549284
rect 298704 549244 298710 549256
rect 299566 549244 299572 549256
rect 299624 549244 299630 549296
rect 226242 549176 226248 549228
rect 226300 549216 226306 549228
rect 449526 549216 449532 549228
rect 226300 549188 449532 549216
rect 226300 549176 226306 549188
rect 449526 549176 449532 549188
rect 449584 549176 449590 549228
rect 223666 549108 223672 549160
rect 223724 549148 223730 549160
rect 449618 549148 449624 549160
rect 223724 549120 449624 549148
rect 223724 549108 223730 549120
rect 449618 549108 449624 549120
rect 449676 549108 449682 549160
rect 218422 549040 218428 549092
rect 218480 549080 218486 549092
rect 449342 549080 449348 549092
rect 218480 549052 449348 549080
rect 218480 549040 218486 549052
rect 449342 549040 449348 549052
rect 449400 549040 449406 549092
rect 2958 548972 2964 549024
rect 3016 549012 3022 549024
rect 355502 549012 355508 549024
rect 3016 548984 355508 549012
rect 3016 548972 3022 548984
rect 355502 548972 355508 548984
rect 355560 548972 355566 549024
rect 4706 548904 4712 548956
rect 4764 548944 4770 548956
rect 365898 548944 365904 548956
rect 4764 548916 365904 548944
rect 4764 548904 4770 548916
rect 365898 548904 365904 548916
rect 365956 548904 365962 548956
rect 5258 548836 5264 548888
rect 5316 548876 5322 548888
rect 371050 548876 371056 548888
rect 5316 548848 371056 548876
rect 5316 548836 5322 548848
rect 371050 548836 371056 548848
rect 371108 548836 371114 548888
rect 3050 548768 3056 548820
rect 3108 548808 3114 548820
rect 368474 548808 368480 548820
rect 3108 548780 368480 548808
rect 3108 548768 3114 548780
rect 368474 548768 368480 548780
rect 368532 548768 368538 548820
rect 5350 548700 5356 548752
rect 5408 548740 5414 548752
rect 373626 548740 373632 548752
rect 5408 548712 373632 548740
rect 5408 548700 5414 548712
rect 373626 548700 373632 548712
rect 373684 548700 373690 548752
rect 3142 548632 3148 548684
rect 3200 548672 3206 548684
rect 376202 548672 376208 548684
rect 3200 548644 376208 548672
rect 3200 548632 3206 548644
rect 376202 548632 376208 548644
rect 376260 548632 376266 548684
rect 5166 548564 5172 548616
rect 5224 548604 5230 548616
rect 378778 548604 378784 548616
rect 5224 548576 378784 548604
rect 5224 548564 5230 548576
rect 378778 548564 378784 548576
rect 378836 548564 378842 548616
rect 6362 548496 6368 548548
rect 6420 548536 6426 548548
rect 381354 548536 381360 548548
rect 6420 548508 381360 548536
rect 6420 548496 6426 548508
rect 381354 548496 381360 548508
rect 381412 548496 381418 548548
rect 3234 548428 3240 548480
rect 3292 548468 3298 548480
rect 384022 548468 384028 548480
rect 3292 548440 384028 548468
rect 3292 548428 3298 548440
rect 384022 548428 384028 548440
rect 384080 548428 384086 548480
rect 6270 548360 6276 548412
rect 6328 548400 6334 548412
rect 389174 548400 389180 548412
rect 6328 548372 389180 548400
rect 6328 548360 6334 548372
rect 389174 548360 389180 548372
rect 389232 548360 389238 548412
rect 4062 548292 4068 548344
rect 4120 548332 4126 548344
rect 391750 548332 391756 548344
rect 4120 548304 391756 548332
rect 4120 548292 4126 548304
rect 391750 548292 391756 548304
rect 391808 548292 391814 548344
rect 5074 548224 5080 548276
rect 5132 548264 5138 548276
rect 394326 548264 394332 548276
rect 5132 548236 394332 548264
rect 5132 548224 5138 548236
rect 394326 548224 394332 548236
rect 394384 548224 394390 548276
rect 6178 548156 6184 548208
rect 6236 548196 6242 548208
rect 396902 548196 396908 548208
rect 6236 548168 396908 548196
rect 6236 548156 6242 548168
rect 396902 548156 396908 548168
rect 396960 548156 396966 548208
rect 10318 548088 10324 548140
rect 10376 548128 10382 548140
rect 404630 548128 404636 548140
rect 10376 548100 404636 548128
rect 10376 548088 10382 548100
rect 404630 548088 404636 548100
rect 404688 548088 404694 548140
rect 3970 548020 3976 548072
rect 4028 548060 4034 548072
rect 399478 548060 399484 548072
rect 4028 548032 399484 548060
rect 4028 548020 4034 548032
rect 399478 548020 399484 548032
rect 399536 548020 399542 548072
rect 19978 547952 19984 548004
rect 20036 547992 20042 548004
rect 420178 547992 420184 548004
rect 20036 547964 420184 547992
rect 20036 547952 20042 547964
rect 420178 547952 420184 547964
rect 420236 547952 420242 548004
rect 4890 547884 4896 547936
rect 4948 547924 4954 547936
rect 409874 547924 409880 547936
rect 4948 547896 409880 547924
rect 4948 547884 4954 547896
rect 409874 547884 409880 547896
rect 409932 547884 409938 547936
rect 149698 545504 149704 545556
rect 149756 545544 149762 545556
rect 401686 545544 401692 545556
rect 149756 545516 401692 545544
rect 149756 545504 149762 545516
rect 401686 545504 401692 545516
rect 401744 545504 401750 545556
rect 184750 545436 184756 545488
rect 184808 545476 184814 545488
rect 449250 545476 449256 545488
rect 184808 545448 449256 545476
rect 184808 545436 184814 545448
rect 449250 545436 449256 545448
rect 449308 545436 449314 545488
rect 177482 545368 177488 545420
rect 177540 545408 177546 545420
rect 449158 545408 449164 545420
rect 177540 545380 449164 545408
rect 177540 545368 177546 545380
rect 449158 545368 449164 545380
rect 449216 545368 449222 545420
rect 242066 545300 242072 545352
rect 242124 545340 242130 545352
rect 580166 545340 580172 545352
rect 242124 545312 580172 545340
rect 242124 545300 242130 545312
rect 580166 545300 580172 545312
rect 580224 545300 580230 545352
rect 5442 545232 5448 545284
rect 5500 545272 5506 545284
rect 363046 545272 363052 545284
rect 5500 545244 363052 545272
rect 5500 545232 5506 545244
rect 363046 545232 363052 545244
rect 363104 545232 363110 545284
rect 192846 545164 192852 545216
rect 192904 545204 192910 545216
rect 580718 545204 580724 545216
rect 192904 545176 580724 545204
rect 192904 545164 192910 545176
rect 580718 545164 580724 545176
rect 580776 545164 580782 545216
rect 187602 545096 187608 545148
rect 187660 545136 187666 545148
rect 580534 545136 580540 545148
rect 187660 545108 580540 545136
rect 187660 545096 187666 545108
rect 580534 545096 580540 545108
rect 580592 545096 580598 545148
rect 236914 544892 236920 544944
rect 236972 544932 236978 544944
rect 449066 544932 449072 544944
rect 236972 544904 449072 544932
rect 236972 544892 236978 544904
rect 449066 544892 449072 544904
rect 449124 544892 449130 544944
rect 229002 544824 229008 544876
rect 229060 544864 229066 544876
rect 449710 544864 449716 544876
rect 229060 544836 449716 544864
rect 229060 544824 229066 544836
rect 449710 544824 449716 544836
rect 449768 544824 449774 544876
rect 216122 544756 216128 544808
rect 216180 544796 216186 544808
rect 449434 544796 449440 544808
rect 216180 544768 449440 544796
rect 216180 544756 216186 544768
rect 449434 544756 449440 544768
rect 449492 544756 449498 544808
rect 161842 544728 161848 544740
rect 161803 544700 161848 544728
rect 161842 544688 161848 544700
rect 161900 544688 161906 544740
rect 164050 544728 164056 544740
rect 164011 544700 164056 544728
rect 164050 544688 164056 544700
rect 164108 544688 164114 544740
rect 169570 544728 169576 544740
rect 169531 544700 169576 544728
rect 169570 544688 169576 544700
rect 169628 544688 169634 544740
rect 172146 544728 172152 544740
rect 172107 544700 172152 544728
rect 172146 544688 172152 544700
rect 172204 544688 172210 544740
rect 174906 544728 174912 544740
rect 174867 544700 174912 544728
rect 174906 544688 174912 544700
rect 174964 544688 174970 544740
rect 180058 544728 180064 544740
rect 180019 544700 180064 544728
rect 180058 544688 180064 544700
rect 180116 544688 180122 544740
rect 182634 544728 182640 544740
rect 182595 544700 182640 544728
rect 182634 544688 182640 544700
rect 182692 544688 182698 544740
rect 195514 544728 195520 544740
rect 195475 544700 195520 544728
rect 195514 544688 195520 544700
rect 195572 544688 195578 544740
rect 200666 544728 200672 544740
rect 200627 544700 200672 544728
rect 200666 544688 200672 544700
rect 200724 544688 200730 544740
rect 234338 544688 234344 544740
rect 234396 544728 234402 544740
rect 580074 544728 580080 544740
rect 234396 544700 580080 544728
rect 234396 544688 234402 544700
rect 580074 544688 580080 544700
rect 580132 544688 580138 544740
rect 6454 544620 6460 544672
rect 6512 544660 6518 544672
rect 360470 544660 360476 544672
rect 6512 544632 360476 544660
rect 6512 544620 6518 544632
rect 360470 544620 360476 544632
rect 360528 544620 360534 544672
rect 412174 544660 412180 544672
rect 412135 544632 412180 544660
rect 412174 544620 412180 544632
rect 412232 544620 412238 544672
rect 417326 544660 417332 544672
rect 417287 544632 417332 544660
rect 417326 544620 417332 544632
rect 417384 544620 417390 544672
rect 427814 544620 427820 544672
rect 427872 544660 427878 544672
rect 432782 544660 432788 544672
rect 427872 544632 427917 544660
rect 432743 544632 432788 544660
rect 427872 544620 427878 544632
rect 432782 544620 432788 544632
rect 432840 544620 432846 544672
rect 438210 544660 438216 544672
rect 438171 544632 438216 544660
rect 438210 544620 438216 544632
rect 438268 544620 438274 544672
rect 443086 544660 443092 544672
rect 443047 544632 443092 544660
rect 443086 544620 443092 544632
rect 443144 544620 443150 544672
rect 200669 544595 200727 544601
rect 200669 544561 200681 544595
rect 200715 544592 200727 544595
rect 580902 544592 580908 544604
rect 200715 544564 580908 544592
rect 200715 544561 200727 544564
rect 200669 544555 200727 544561
rect 580902 544552 580908 544564
rect 580960 544552 580966 544604
rect 195517 544527 195575 544533
rect 195517 544493 195529 544527
rect 195563 544524 195575 544527
rect 580626 544524 580632 544536
rect 195563 544496 580632 544524
rect 195563 544493 195575 544496
rect 195517 544487 195575 544493
rect 580626 544484 580632 544496
rect 580684 544484 580690 544536
rect 182637 544459 182695 544465
rect 182637 544425 182649 544459
rect 182683 544456 182695 544459
rect 578050 544456 578056 544468
rect 182683 544428 578056 544456
rect 182683 544425 182695 544428
rect 182637 544419 182695 544425
rect 578050 544416 578056 544428
rect 578108 544416 578114 544468
rect 180061 544391 180119 544397
rect 180061 544357 180073 544391
rect 180107 544388 180119 544391
rect 580442 544388 580448 544400
rect 180107 544360 580448 544388
rect 180107 544357 180119 544360
rect 180061 544351 180119 544357
rect 580442 544348 580448 544360
rect 580500 544348 580506 544400
rect 174909 544323 174967 544329
rect 174909 544289 174921 544323
rect 174955 544320 174967 544323
rect 577958 544320 577964 544332
rect 174955 544292 577964 544320
rect 174955 544289 174967 544292
rect 174909 544283 174967 544289
rect 577958 544280 577964 544292
rect 578016 544280 578022 544332
rect 4982 544212 4988 544264
rect 5040 544252 5046 544264
rect 412177 544255 412235 544261
rect 412177 544252 412189 544255
rect 5040 544224 412189 544252
rect 5040 544212 5046 544224
rect 412177 544221 412189 544224
rect 412223 544221 412235 544255
rect 412177 544215 412235 544221
rect 172149 544187 172207 544193
rect 172149 544153 172161 544187
rect 172195 544184 172207 544187
rect 580350 544184 580356 544196
rect 172195 544156 580356 544184
rect 172195 544153 172207 544156
rect 172149 544147 172207 544153
rect 580350 544144 580356 544156
rect 580408 544144 580414 544196
rect 169573 544119 169631 544125
rect 169573 544085 169585 544119
rect 169619 544116 169631 544119
rect 577866 544116 577872 544128
rect 169619 544088 577872 544116
rect 169619 544085 169631 544088
rect 169573 544079 169631 544085
rect 577866 544076 577872 544088
rect 577924 544076 577930 544128
rect 3878 544008 3884 544060
rect 3936 544048 3942 544060
rect 417329 544051 417387 544057
rect 417329 544048 417341 544051
rect 3936 544020 417341 544048
rect 3936 544008 3942 544020
rect 417329 544017 417341 544020
rect 417375 544017 417387 544051
rect 417329 544011 417387 544017
rect 164053 543983 164111 543989
rect 164053 543949 164065 543983
rect 164099 543980 164111 543983
rect 577682 543980 577688 543992
rect 164099 543952 577688 543980
rect 164099 543949 164111 543952
rect 164053 543943 164111 543949
rect 577682 543940 577688 543952
rect 577740 543940 577746 543992
rect 3786 543872 3792 543924
rect 3844 543912 3850 543924
rect 427817 543915 427875 543921
rect 427817 543912 427829 543915
rect 3844 543884 427829 543912
rect 3844 543872 3850 543884
rect 427817 543881 427829 543884
rect 427863 543881 427875 543915
rect 427817 543875 427875 543881
rect 3602 543804 3608 543856
rect 3660 543844 3666 543856
rect 432785 543847 432843 543853
rect 432785 543844 432797 543847
rect 3660 543816 432797 543844
rect 3660 543804 3666 543816
rect 432785 543813 432797 543816
rect 432831 543813 432843 543847
rect 432785 543807 432843 543813
rect 3418 543736 3424 543788
rect 3476 543776 3482 543788
rect 443089 543779 443147 543785
rect 443089 543776 443101 543779
rect 3476 543748 443101 543776
rect 3476 543736 3482 543748
rect 443089 543745 443101 543748
rect 443135 543745 443147 543779
rect 443089 543739 443147 543745
rect 438213 543711 438271 543717
rect 438213 543708 438225 543711
rect 437400 543680 438225 543708
rect 164237 543235 164295 543241
rect 164237 543201 164249 543235
rect 164283 543232 164295 543235
rect 168929 543235 168987 543241
rect 168929 543232 168941 543235
rect 164283 543204 168941 543232
rect 164283 543201 164295 543204
rect 164237 543195 164295 543201
rect 168929 543201 168941 543204
rect 168975 543201 168987 543235
rect 168929 543195 168987 543201
rect 183557 543235 183615 543241
rect 183557 543201 183569 543235
rect 183603 543232 183615 543235
rect 188249 543235 188307 543241
rect 188249 543232 188261 543235
rect 183603 543204 188261 543232
rect 183603 543201 183615 543204
rect 183557 543195 183615 543201
rect 188249 543201 188261 543204
rect 188295 543201 188307 543235
rect 188249 543195 188307 543201
rect 202877 543235 202935 543241
rect 202877 543201 202889 543235
rect 202923 543232 202935 543235
rect 207569 543235 207627 543241
rect 207569 543232 207581 543235
rect 202923 543204 207581 543232
rect 202923 543201 202935 543204
rect 202877 543195 202935 543201
rect 207569 543201 207581 543204
rect 207615 543201 207627 543235
rect 207569 543195 207627 543201
rect 249797 543235 249855 543241
rect 249797 543201 249809 543235
rect 249843 543232 249855 543235
rect 259365 543235 259423 543241
rect 259365 543232 259377 543235
rect 249843 543204 259377 543232
rect 249843 543201 249855 543204
rect 249797 543195 249855 543201
rect 259365 543201 259377 543204
rect 259411 543201 259423 543235
rect 259365 543195 259423 543201
rect 280157 543235 280215 543241
rect 280157 543201 280169 543235
rect 280203 543232 280215 543235
rect 284849 543235 284907 543241
rect 284849 543232 284861 543235
rect 280203 543204 284861 543232
rect 280203 543201 280215 543204
rect 280157 543195 280215 543201
rect 284849 543201 284861 543204
rect 284895 543201 284907 543235
rect 284849 543195 284907 543201
rect 318797 543235 318855 543241
rect 318797 543201 318809 543235
rect 318843 543232 318855 543235
rect 323489 543235 323547 543241
rect 323489 543232 323501 543235
rect 318843 543204 323501 543232
rect 318843 543201 318855 543204
rect 318797 543195 318855 543201
rect 323489 543201 323501 543204
rect 323535 543201 323547 543235
rect 424965 543235 425023 543241
rect 424965 543232 424977 543235
rect 323489 543195 323547 543201
rect 417988 543204 424977 543232
rect 144917 543167 144975 543173
rect 144917 543133 144929 543167
rect 144963 543164 144975 543167
rect 154485 543167 154543 543173
rect 154485 543164 154497 543167
rect 144963 543136 154497 543164
rect 144963 543133 144975 543136
rect 144917 543127 144975 543133
rect 154485 543133 154497 543136
rect 154531 543133 154543 543167
rect 154485 543127 154543 543133
rect 176473 543167 176531 543173
rect 176473 543133 176485 543167
rect 176519 543164 176531 543167
rect 183465 543167 183523 543173
rect 183465 543164 183477 543167
rect 176519 543136 183477 543164
rect 176519 543133 176531 543136
rect 176473 543127 176531 543133
rect 183465 543133 183477 543136
rect 183511 543133 183523 543167
rect 183465 543127 183523 543133
rect 193309 543167 193367 543173
rect 193309 543133 193321 543167
rect 193355 543164 193367 543167
rect 202785 543167 202843 543173
rect 202785 543164 202797 543167
rect 193355 543136 202797 543164
rect 193355 543133 193367 543136
rect 193309 543127 193367 543133
rect 202785 543133 202797 543136
rect 202831 543133 202843 543167
rect 202785 543127 202843 543133
rect 211157 543167 211215 543173
rect 211157 543133 211169 543167
rect 211203 543164 211215 543167
rect 220725 543167 220783 543173
rect 220725 543164 220737 543167
rect 211203 543136 220737 543164
rect 211203 543133 211215 543136
rect 211157 543127 211215 543133
rect 220725 543133 220737 543136
rect 220771 543133 220783 543167
rect 220725 543127 220783 543133
rect 273073 543167 273131 543173
rect 273073 543133 273085 543167
rect 273119 543164 273131 543167
rect 280065 543167 280123 543173
rect 280065 543164 280077 543167
rect 273119 543136 280077 543164
rect 273119 543133 273131 543136
rect 273073 543127 273131 543133
rect 280065 543133 280077 543136
rect 280111 543133 280123 543167
rect 280065 543127 280123 543133
rect 292393 543167 292451 543173
rect 292393 543133 292405 543167
rect 292439 543164 292451 543167
rect 299385 543167 299443 543173
rect 299385 543164 299397 543167
rect 292439 543136 299397 543164
rect 292439 543133 292451 543136
rect 292393 543127 292451 543133
rect 299385 543133 299397 543136
rect 299431 543133 299443 543167
rect 299385 543127 299443 543133
rect 299477 543167 299535 543173
rect 299477 543133 299489 543167
rect 299523 543164 299535 543167
rect 308861 543167 308919 543173
rect 308861 543164 308873 543167
rect 299523 543136 308873 543164
rect 299523 543133 299535 543136
rect 299477 543127 299535 543133
rect 308861 543133 308873 543136
rect 308907 543133 308919 543167
rect 308861 543127 308919 543133
rect 311713 543167 311771 543173
rect 311713 543133 311725 543167
rect 311759 543164 311771 543167
rect 318705 543167 318763 543173
rect 318705 543164 318717 543167
rect 311759 543136 318717 543164
rect 311759 543133 311771 543136
rect 311713 543127 311771 543133
rect 318705 543133 318717 543136
rect 318751 543133 318763 543167
rect 318705 543127 318763 543133
rect 346581 543167 346639 543173
rect 346581 543133 346593 543167
rect 346627 543164 346639 543167
rect 355965 543167 356023 543173
rect 355965 543164 355977 543167
rect 346627 543136 355977 543164
rect 346627 543133 346639 543136
rect 346581 543127 346639 543133
rect 355965 543133 355977 543136
rect 356011 543133 356023 543167
rect 355965 543127 356023 543133
rect 19337 543099 19395 543105
rect 19337 543065 19349 543099
rect 19383 543096 19395 543099
rect 28905 543099 28963 543105
rect 28905 543096 28917 543099
rect 19383 543068 28917 543096
rect 19383 543065 19395 543068
rect 19337 543059 19395 543065
rect 28905 543065 28917 543068
rect 28951 543065 28963 543099
rect 28905 543059 28963 543065
rect 38657 543099 38715 543105
rect 38657 543065 38669 543099
rect 38703 543096 38715 543099
rect 48225 543099 48283 543105
rect 48225 543096 48237 543099
rect 38703 543068 48237 543096
rect 38703 543065 38715 543068
rect 38657 543059 38715 543065
rect 48225 543065 48237 543068
rect 48271 543065 48283 543099
rect 48225 543059 48283 543065
rect 57977 543099 58035 543105
rect 57977 543065 57989 543099
rect 58023 543096 58035 543099
rect 67545 543099 67603 543105
rect 67545 543096 67557 543099
rect 58023 543068 67557 543096
rect 58023 543065 58035 543068
rect 57977 543059 58035 543065
rect 67545 543065 67557 543068
rect 67591 543065 67603 543099
rect 67545 543059 67603 543065
rect 77297 543099 77355 543105
rect 77297 543065 77309 543099
rect 77343 543096 77355 543099
rect 86865 543099 86923 543105
rect 86865 543096 86877 543099
rect 77343 543068 86877 543096
rect 77343 543065 77355 543068
rect 77297 543059 77355 543065
rect 86865 543065 86877 543068
rect 86911 543065 86923 543099
rect 86865 543059 86923 543065
rect 96617 543099 96675 543105
rect 96617 543065 96629 543099
rect 96663 543096 96675 543099
rect 106185 543099 106243 543105
rect 106185 543096 106197 543099
rect 96663 543068 106197 543096
rect 96663 543065 96675 543068
rect 96617 543059 96675 543065
rect 106185 543065 106197 543068
rect 106231 543065 106243 543099
rect 106185 543059 106243 543065
rect 115937 543099 115995 543105
rect 115937 543065 115949 543099
rect 115983 543096 115995 543099
rect 125505 543099 125563 543105
rect 125505 543096 125517 543099
rect 115983 543068 125517 543096
rect 115983 543065 115995 543068
rect 115937 543059 115995 543065
rect 125505 543065 125517 543068
rect 125551 543065 125563 543099
rect 125505 543059 125563 543065
rect 173897 543099 173955 543105
rect 173897 543065 173909 543099
rect 173943 543096 173955 543099
rect 178681 543099 178739 543105
rect 178681 543096 178693 543099
rect 173943 543068 178693 543096
rect 173943 543065 173955 543068
rect 173897 543059 173955 543065
rect 178681 543065 178693 543068
rect 178727 543065 178739 543099
rect 178681 543059 178739 543065
rect 193217 543099 193275 543105
rect 193217 543065 193229 543099
rect 193263 543096 193275 543099
rect 198001 543099 198059 543105
rect 198001 543096 198013 543099
rect 193263 543068 198013 543096
rect 193263 543065 193275 543068
rect 193217 543059 193275 543065
rect 198001 543065 198013 543068
rect 198047 543065 198059 543099
rect 249797 543099 249855 543105
rect 249797 543096 249809 543099
rect 198001 543059 198059 543065
rect 234448 543068 249809 543096
rect 144917 543031 144975 543037
rect 144917 543028 144929 543031
rect 138216 543000 144929 543028
rect 12437 542963 12495 542969
rect 12437 542929 12449 542963
rect 12483 542960 12495 542963
rect 19337 542963 19395 542969
rect 19337 542960 19349 542963
rect 12483 542932 19349 542960
rect 12483 542929 12495 542932
rect 12437 542923 12495 542929
rect 19337 542929 19349 542932
rect 19383 542929 19395 542963
rect 19337 542923 19395 542929
rect 31757 542963 31815 542969
rect 31757 542929 31769 542963
rect 31803 542960 31815 542963
rect 38657 542963 38715 542969
rect 38657 542960 38669 542963
rect 31803 542932 38669 542960
rect 31803 542929 31815 542932
rect 31757 542923 31815 542929
rect 38657 542929 38669 542932
rect 38703 542929 38715 542963
rect 38657 542923 38715 542929
rect 51077 542963 51135 542969
rect 51077 542929 51089 542963
rect 51123 542960 51135 542963
rect 57977 542963 58035 542969
rect 57977 542960 57989 542963
rect 51123 542932 57989 542960
rect 51123 542929 51135 542932
rect 51077 542923 51135 542929
rect 57977 542929 57989 542932
rect 58023 542929 58035 542963
rect 57977 542923 58035 542929
rect 70397 542963 70455 542969
rect 70397 542929 70409 542963
rect 70443 542960 70455 542963
rect 77297 542963 77355 542969
rect 77297 542960 77309 542963
rect 70443 542932 77309 542960
rect 70443 542929 70455 542932
rect 70397 542923 70455 542929
rect 77297 542929 77309 542932
rect 77343 542929 77355 542963
rect 77297 542923 77355 542929
rect 89717 542963 89775 542969
rect 89717 542929 89729 542963
rect 89763 542960 89775 542963
rect 96617 542963 96675 542969
rect 96617 542960 96629 542963
rect 89763 542932 96629 542960
rect 89763 542929 89775 542932
rect 89717 542923 89775 542929
rect 96617 542929 96629 542932
rect 96663 542929 96675 542963
rect 96617 542923 96675 542929
rect 109037 542963 109095 542969
rect 109037 542929 109049 542963
rect 109083 542960 109095 542963
rect 115937 542963 115995 542969
rect 115937 542960 115949 542963
rect 109083 542932 115949 542960
rect 109083 542929 109095 542932
rect 109037 542923 109095 542929
rect 115937 542929 115949 542932
rect 115983 542929 115995 542963
rect 115937 542923 115995 542929
rect 128357 542963 128415 542969
rect 128357 542929 128369 542963
rect 128403 542960 128415 542963
rect 137925 542963 137983 542969
rect 137925 542960 137937 542963
rect 128403 542932 137937 542960
rect 128403 542929 128415 542932
rect 128357 542923 128415 542929
rect 137925 542929 137937 542932
rect 137971 542929 137983 542963
rect 137925 542923 137983 542929
rect 138017 542963 138075 542969
rect 138017 542929 138029 542963
rect 138063 542960 138075 542963
rect 138216 542960 138244 543000
rect 144917 542997 144929 543000
rect 144963 542997 144975 543031
rect 144917 542991 144975 542997
rect 168837 543031 168895 543037
rect 168837 542997 168849 543031
rect 168883 543028 168895 543031
rect 173805 543031 173863 543037
rect 173805 543028 173817 543031
rect 168883 543000 173817 543028
rect 168883 542997 168895 543000
rect 168837 542991 168895 542997
rect 173805 542997 173817 543000
rect 173851 542997 173863 543031
rect 173805 542991 173863 542997
rect 188157 543031 188215 543037
rect 188157 542997 188169 543031
rect 188203 543028 188215 543031
rect 193125 543031 193183 543037
rect 193125 543028 193137 543031
rect 188203 543000 193137 543028
rect 188203 542997 188215 543000
rect 188157 542991 188215 542997
rect 193125 542997 193137 543000
rect 193171 542997 193183 543031
rect 193125 542991 193183 542997
rect 207477 543031 207535 543037
rect 207477 542997 207489 543031
rect 207523 543028 207535 543031
rect 215757 543031 215815 543037
rect 215757 543028 215769 543031
rect 207523 543000 215769 543028
rect 207523 542997 207535 543000
rect 207477 542991 207535 542997
rect 215757 542997 215769 543000
rect 215803 542997 215815 543031
rect 215757 542991 215815 542997
rect 138063 542932 138244 542960
rect 154669 542963 154727 542969
rect 138063 542929 138075 542932
rect 138017 542923 138075 542929
rect 154669 542929 154681 542963
rect 154715 542960 154727 542963
rect 164237 542963 164295 542969
rect 164237 542960 164249 542963
rect 154715 542932 164249 542960
rect 154715 542929 154727 542932
rect 154669 542923 154727 542929
rect 164237 542929 164249 542932
rect 164283 542929 164295 542963
rect 164237 542923 164295 542929
rect 183465 542963 183523 542969
rect 183465 542929 183477 542963
rect 183511 542960 183523 542963
rect 183557 542963 183615 542969
rect 183557 542960 183569 542963
rect 183511 542932 183569 542960
rect 183511 542929 183523 542932
rect 183465 542923 183523 542929
rect 183557 542929 183569 542932
rect 183603 542929 183615 542963
rect 183557 542923 183615 542929
rect 202785 542963 202843 542969
rect 202785 542929 202797 542963
rect 202831 542960 202843 542963
rect 202877 542963 202935 542969
rect 202877 542960 202889 542963
rect 202831 542932 202889 542960
rect 202831 542929 202843 542932
rect 202785 542923 202843 542929
rect 202877 542929 202889 542932
rect 202923 542929 202935 542963
rect 202877 542923 202935 542929
rect 220725 542963 220783 542969
rect 220725 542929 220737 542963
rect 220771 542960 220783 542963
rect 234448 542960 234476 543068
rect 249797 543065 249809 543068
rect 249843 543065 249855 543099
rect 249797 543059 249855 543065
rect 270497 543099 270555 543105
rect 270497 543065 270509 543099
rect 270543 543096 270555 543099
rect 275281 543099 275339 543105
rect 275281 543096 275293 543099
rect 270543 543068 275293 543096
rect 270543 543065 270555 543068
rect 270497 543059 270555 543065
rect 275281 543065 275293 543068
rect 275327 543065 275339 543099
rect 275281 543059 275339 543065
rect 289817 543099 289875 543105
rect 289817 543065 289829 543099
rect 289863 543096 289875 543099
rect 294601 543099 294659 543105
rect 294601 543096 294613 543099
rect 289863 543068 294613 543096
rect 289863 543065 289875 543068
rect 289817 543059 289875 543065
rect 294601 543065 294613 543068
rect 294647 543065 294659 543099
rect 294601 543059 294659 543065
rect 309137 543099 309195 543105
rect 309137 543065 309149 543099
rect 309183 543096 309195 543099
rect 313921 543099 313979 543105
rect 313921 543096 313933 543099
rect 309183 543068 313933 543096
rect 309183 543065 309195 543068
rect 309137 543059 309195 543065
rect 313921 543065 313933 543068
rect 313967 543065 313979 543099
rect 313921 543059 313979 543065
rect 327077 543099 327135 543105
rect 327077 543065 327089 543099
rect 327123 543096 327135 543099
rect 417988 543096 418016 543204
rect 424965 543201 424977 543204
rect 425011 543201 425023 543235
rect 424965 543195 425023 543201
rect 437400 543164 437428 543680
rect 438213 543677 438225 543680
rect 438259 543677 438271 543711
rect 438213 543671 438271 543677
rect 427832 543136 437428 543164
rect 327123 543068 336688 543096
rect 327123 543065 327135 543068
rect 327077 543059 327135 543065
rect 259365 543031 259423 543037
rect 259365 542997 259377 543031
rect 259411 543028 259423 543031
rect 265161 543031 265219 543037
rect 265161 543028 265173 543031
rect 259411 543000 265173 543028
rect 259411 542997 259423 543000
rect 259365 542991 259423 542997
rect 265161 542997 265173 543000
rect 265207 542997 265219 543031
rect 265161 542991 265219 542997
rect 284757 543031 284815 543037
rect 284757 542997 284769 543031
rect 284803 543028 284815 543031
rect 289725 543031 289783 543037
rect 289725 543028 289737 543031
rect 284803 543000 289737 543028
rect 284803 542997 284815 543000
rect 284757 542991 284815 542997
rect 289725 542997 289737 543000
rect 289771 542997 289783 543031
rect 323397 543031 323455 543037
rect 289725 542991 289783 542997
rect 299492 543000 304212 543028
rect 220771 542932 234476 542960
rect 263689 542963 263747 542969
rect 220771 542929 220783 542932
rect 220725 542923 220783 542929
rect 263689 542929 263701 542963
rect 263735 542960 263747 542963
rect 280065 542963 280123 542969
rect 263735 542932 270448 542960
rect 263735 542929 263747 542932
rect 263689 542923 263747 542929
rect 28905 542895 28963 542901
rect 28905 542861 28917 542895
rect 28951 542892 28963 542895
rect 48225 542895 48283 542901
rect 28951 542864 31708 542892
rect 28951 542861 28963 542864
rect 28905 542855 28963 542861
rect 3510 542784 3516 542836
rect 3568 542824 3574 542836
rect 12437 542827 12495 542833
rect 12437 542824 12449 542827
rect 3568 542796 12449 542824
rect 3568 542784 3574 542796
rect 12437 542793 12449 542796
rect 12483 542793 12495 542827
rect 31680 542824 31708 542864
rect 48225 542861 48237 542895
rect 48271 542892 48283 542895
rect 67545 542895 67603 542901
rect 48271 542864 51028 542892
rect 48271 542861 48283 542864
rect 48225 542855 48283 542861
rect 31757 542827 31815 542833
rect 31757 542824 31769 542827
rect 31680 542796 31769 542824
rect 12437 542787 12495 542793
rect 31757 542793 31769 542796
rect 31803 542793 31815 542827
rect 51000 542824 51028 542864
rect 67545 542861 67557 542895
rect 67591 542892 67603 542895
rect 86865 542895 86923 542901
rect 67591 542864 70348 542892
rect 67591 542861 67603 542864
rect 67545 542855 67603 542861
rect 51077 542827 51135 542833
rect 51077 542824 51089 542827
rect 51000 542796 51089 542824
rect 31757 542787 31815 542793
rect 51077 542793 51089 542796
rect 51123 542793 51135 542827
rect 70320 542824 70348 542864
rect 86865 542861 86877 542895
rect 86911 542892 86923 542895
rect 106185 542895 106243 542901
rect 86911 542864 89668 542892
rect 86911 542861 86923 542864
rect 86865 542855 86923 542861
rect 70397 542827 70455 542833
rect 70397 542824 70409 542827
rect 70320 542796 70409 542824
rect 51077 542787 51135 542793
rect 70397 542793 70409 542796
rect 70443 542793 70455 542827
rect 89640 542824 89668 542864
rect 106185 542861 106197 542895
rect 106231 542892 106243 542895
rect 125505 542895 125563 542901
rect 106231 542864 108988 542892
rect 106231 542861 106243 542864
rect 106185 542855 106243 542861
rect 89717 542827 89775 542833
rect 89717 542824 89729 542827
rect 89640 542796 89729 542824
rect 70397 542787 70455 542793
rect 89717 542793 89729 542796
rect 89763 542793 89775 542827
rect 108960 542824 108988 542864
rect 125505 542861 125517 542895
rect 125551 542892 125563 542895
rect 154485 542895 154543 542901
rect 125551 542864 128308 542892
rect 125551 542861 125563 542864
rect 125505 542855 125563 542861
rect 109037 542827 109095 542833
rect 109037 542824 109049 542827
rect 108960 542796 109049 542824
rect 89717 542787 89775 542793
rect 109037 542793 109049 542796
rect 109083 542793 109095 542827
rect 128280 542824 128308 542864
rect 154485 542861 154497 542895
rect 154531 542892 154543 542895
rect 154577 542895 154635 542901
rect 154577 542892 154589 542895
rect 154531 542864 154589 542892
rect 154531 542861 154543 542864
rect 154485 542855 154543 542861
rect 154577 542861 154589 542864
rect 154623 542861 154635 542895
rect 154577 542855 154635 542861
rect 161845 542895 161903 542901
rect 161845 542861 161857 542895
rect 161891 542892 161903 542895
rect 168837 542895 168895 542901
rect 168837 542892 168849 542895
rect 161891 542864 168849 542892
rect 161891 542861 161903 542864
rect 161845 542855 161903 542861
rect 168837 542861 168849 542864
rect 168883 542861 168895 542895
rect 168837 542855 168895 542861
rect 168929 542895 168987 542901
rect 168929 542861 168941 542895
rect 168975 542861 168987 542895
rect 168929 542855 168987 542861
rect 173805 542895 173863 542901
rect 173805 542861 173817 542895
rect 173851 542892 173863 542895
rect 173897 542895 173955 542901
rect 173897 542892 173909 542895
rect 173851 542864 173909 542892
rect 173851 542861 173863 542864
rect 173805 542855 173863 542861
rect 173897 542861 173909 542864
rect 173943 542861 173955 542895
rect 173897 542855 173955 542861
rect 176473 542895 176531 542901
rect 176473 542861 176485 542895
rect 176519 542861 176531 542895
rect 176473 542855 176531 542861
rect 178681 542895 178739 542901
rect 178681 542861 178693 542895
rect 178727 542892 178739 542895
rect 188157 542895 188215 542901
rect 188157 542892 188169 542895
rect 178727 542864 188169 542892
rect 178727 542861 178739 542864
rect 178681 542855 178739 542861
rect 188157 542861 188169 542864
rect 188203 542861 188215 542895
rect 188157 542855 188215 542861
rect 188249 542895 188307 542901
rect 188249 542861 188261 542895
rect 188295 542861 188307 542895
rect 188249 542855 188307 542861
rect 193125 542895 193183 542901
rect 193125 542861 193137 542895
rect 193171 542892 193183 542895
rect 193217 542895 193275 542901
rect 193217 542892 193229 542895
rect 193171 542864 193229 542892
rect 193171 542861 193183 542864
rect 193125 542855 193183 542861
rect 193217 542861 193229 542864
rect 193263 542861 193275 542895
rect 193217 542855 193275 542861
rect 193309 542895 193367 542901
rect 193309 542861 193321 542895
rect 193355 542861 193367 542895
rect 193309 542855 193367 542861
rect 198001 542895 198059 542901
rect 198001 542861 198013 542895
rect 198047 542892 198059 542895
rect 207477 542895 207535 542901
rect 207477 542892 207489 542895
rect 198047 542864 207489 542892
rect 198047 542861 198059 542864
rect 198001 542855 198059 542861
rect 207477 542861 207489 542864
rect 207523 542861 207535 542895
rect 207477 542855 207535 542861
rect 207569 542895 207627 542901
rect 207569 542861 207581 542895
rect 207615 542861 207627 542895
rect 207569 542855 207627 542861
rect 211157 542895 211215 542901
rect 211157 542861 211169 542895
rect 211203 542861 211215 542895
rect 211157 542855 211215 542861
rect 215757 542895 215815 542901
rect 215757 542861 215769 542895
rect 215803 542892 215815 542895
rect 241517 542895 241575 542901
rect 241517 542892 241529 542895
rect 215803 542864 241529 542892
rect 215803 542861 215815 542864
rect 215757 542855 215815 542861
rect 241517 542861 241529 542864
rect 241563 542861 241575 542895
rect 241517 542855 241575 542861
rect 241701 542895 241759 542901
rect 241701 542861 241713 542895
rect 241747 542892 241759 542895
rect 263505 542895 263563 542901
rect 263505 542892 263517 542895
rect 241747 542864 263517 542892
rect 241747 542861 241759 542864
rect 241701 542855 241759 542861
rect 263505 542861 263517 542864
rect 263551 542861 263563 542895
rect 263505 542855 263563 542861
rect 265161 542895 265219 542901
rect 265161 542861 265173 542895
rect 265207 542861 265219 542895
rect 270420 542892 270448 542932
rect 280065 542929 280077 542963
rect 280111 542960 280123 542963
rect 280157 542963 280215 542969
rect 280157 542960 280169 542963
rect 280111 542932 280169 542960
rect 280111 542929 280123 542932
rect 280065 542923 280123 542929
rect 280157 542929 280169 542932
rect 280203 542929 280215 542963
rect 280157 542923 280215 542929
rect 299385 542963 299443 542969
rect 299385 542929 299397 542963
rect 299431 542960 299443 542963
rect 299492 542960 299520 543000
rect 299431 542932 299520 542960
rect 299431 542929 299443 542932
rect 299385 542923 299443 542929
rect 270497 542895 270555 542901
rect 270497 542892 270509 542895
rect 270420 542864 270509 542892
rect 265161 542855 265219 542861
rect 270497 542861 270509 542864
rect 270543 542861 270555 542895
rect 270497 542855 270555 542861
rect 273073 542895 273131 542901
rect 273073 542861 273085 542895
rect 273119 542861 273131 542895
rect 273073 542855 273131 542861
rect 275281 542895 275339 542901
rect 275281 542861 275293 542895
rect 275327 542892 275339 542895
rect 284757 542895 284815 542901
rect 284757 542892 284769 542895
rect 275327 542864 284769 542892
rect 275327 542861 275339 542864
rect 275281 542855 275339 542861
rect 284757 542861 284769 542864
rect 284803 542861 284815 542895
rect 284757 542855 284815 542861
rect 284849 542895 284907 542901
rect 284849 542861 284861 542895
rect 284895 542861 284907 542895
rect 284849 542855 284907 542861
rect 289725 542895 289783 542901
rect 289725 542861 289737 542895
rect 289771 542892 289783 542895
rect 289817 542895 289875 542901
rect 289817 542892 289829 542895
rect 289771 542864 289829 542892
rect 289771 542861 289783 542864
rect 289725 542855 289783 542861
rect 289817 542861 289829 542864
rect 289863 542861 289875 542895
rect 289817 542855 289875 542861
rect 292393 542895 292451 542901
rect 292393 542861 292405 542895
rect 292439 542861 292451 542895
rect 292393 542855 292451 542861
rect 294601 542895 294659 542901
rect 294601 542861 294613 542895
rect 294647 542892 294659 542895
rect 299477 542895 299535 542901
rect 299477 542892 299489 542895
rect 294647 542864 299489 542892
rect 294647 542861 294659 542864
rect 294601 542855 294659 542861
rect 299477 542861 299489 542864
rect 299523 542861 299535 542895
rect 299477 542855 299535 542861
rect 128357 542827 128415 542833
rect 128357 542824 128369 542827
rect 128280 542796 128369 542824
rect 109037 542787 109095 542793
rect 128357 542793 128369 542796
rect 128403 542793 128415 542827
rect 168944 542824 168972 542855
rect 176488 542824 176516 542855
rect 168944 542796 176516 542824
rect 188264 542824 188292 542855
rect 193324 542824 193352 542855
rect 188264 542796 193352 542824
rect 207584 542824 207612 542855
rect 211172 542824 211200 542855
rect 207584 542796 211200 542824
rect 265176 542824 265204 542855
rect 273088 542824 273116 542855
rect 265176 542796 273116 542824
rect 284864 542824 284892 542855
rect 292408 542824 292436 542855
rect 284864 542796 292436 542824
rect 304184 542824 304212 543000
rect 323397 542997 323409 543031
rect 323443 543028 323455 543031
rect 328457 543031 328515 543037
rect 328457 543028 328469 543031
rect 323443 543000 328469 543028
rect 323443 542997 323455 543000
rect 323397 542991 323455 542997
rect 328457 542997 328469 543000
rect 328503 542997 328515 543031
rect 328457 542991 328515 542997
rect 318705 542963 318763 542969
rect 318705 542929 318717 542963
rect 318751 542960 318763 542963
rect 318797 542963 318855 542969
rect 318797 542960 318809 542963
rect 318751 542932 318809 542960
rect 318751 542929 318763 542932
rect 318705 542923 318763 542929
rect 318797 542929 318809 542932
rect 318843 542929 318855 542963
rect 318797 542923 318855 542929
rect 328549 542963 328607 542969
rect 328549 542929 328561 542963
rect 328595 542960 328607 542963
rect 336660 542960 336688 543068
rect 346504 543068 355916 543096
rect 346504 542960 346532 543068
rect 328595 542932 331720 542960
rect 336660 542932 346532 542960
rect 346581 542963 346639 542969
rect 328595 542929 328607 542932
rect 328549 542923 328607 542929
rect 309045 542895 309103 542901
rect 309045 542861 309057 542895
rect 309091 542892 309103 542895
rect 309137 542895 309195 542901
rect 309137 542892 309149 542895
rect 309091 542864 309149 542892
rect 309091 542861 309103 542864
rect 309045 542855 309103 542861
rect 309137 542861 309149 542864
rect 309183 542861 309195 542895
rect 309137 542855 309195 542861
rect 311713 542895 311771 542901
rect 311713 542861 311725 542895
rect 311759 542861 311771 542895
rect 311713 542855 311771 542861
rect 313921 542895 313979 542901
rect 313921 542861 313933 542895
rect 313967 542892 313979 542895
rect 323397 542895 323455 542901
rect 323397 542892 323409 542895
rect 313967 542864 323409 542892
rect 313967 542861 313979 542864
rect 313921 542855 313979 542861
rect 323397 542861 323409 542864
rect 323443 542861 323455 542895
rect 323397 542855 323455 542861
rect 323489 542895 323547 542901
rect 323489 542861 323501 542895
rect 323535 542861 323547 542895
rect 323489 542855 323547 542861
rect 327077 542895 327135 542901
rect 327077 542861 327089 542895
rect 327123 542861 327135 542895
rect 331692 542892 331720 542932
rect 346581 542929 346593 542963
rect 346627 542929 346639 542963
rect 346581 542923 346639 542929
rect 346596 542892 346624 542923
rect 331692 542864 346624 542892
rect 327077 542855 327135 542861
rect 311728 542824 311756 542855
rect 304184 542796 311756 542824
rect 323504 542824 323532 542855
rect 327092 542824 327120 542855
rect 323504 542796 327120 542824
rect 355888 542824 355916 543068
rect 408696 543068 418016 543096
rect 424965 543099 425023 543105
rect 355965 543031 356023 543037
rect 355965 542997 355977 543031
rect 356011 542997 356023 543031
rect 355965 542991 356023 542997
rect 365809 543031 365867 543037
rect 365809 542997 365821 543031
rect 365855 543028 365867 543031
rect 370041 543031 370099 543037
rect 365855 543000 369992 543028
rect 365855 542997 365867 543000
rect 365809 542991 365867 542997
rect 355980 542892 356008 542991
rect 365809 542895 365867 542901
rect 365809 542892 365821 542895
rect 355980 542864 365821 542892
rect 365809 542861 365821 542864
rect 365855 542861 365867 542895
rect 369765 542895 369823 542901
rect 369765 542892 369777 542895
rect 365809 542855 365867 542861
rect 369688 542864 369777 542892
rect 369688 542824 369716 542864
rect 369765 542861 369777 542864
rect 369811 542861 369823 542895
rect 369964 542892 369992 543000
rect 370041 542997 370053 543031
rect 370087 543028 370099 543031
rect 389085 543031 389143 543037
rect 389085 543028 389097 543031
rect 370087 543000 389097 543028
rect 370087 542997 370099 543000
rect 370041 542991 370099 542997
rect 389085 542997 389097 543000
rect 389131 542997 389143 543031
rect 389085 542991 389143 542997
rect 389177 543031 389235 543037
rect 389177 542997 389189 543031
rect 389223 543028 389235 543031
rect 398745 543031 398803 543037
rect 398745 543028 398757 543031
rect 389223 543000 398757 543028
rect 389223 542997 389235 543000
rect 389177 542991 389235 542997
rect 398745 542997 398757 543000
rect 398791 542997 398803 543031
rect 398745 542991 398803 542997
rect 398929 543031 398987 543037
rect 398929 542997 398941 543031
rect 398975 543028 398987 543031
rect 408696 543028 408724 543068
rect 424965 543065 424977 543099
rect 425011 543096 425023 543099
rect 427832 543096 427860 543136
rect 425011 543068 427860 543096
rect 425011 543065 425023 543068
rect 424965 543059 425023 543065
rect 398975 543000 400904 543028
rect 398975 542997 398987 543000
rect 398929 542991 398987 542997
rect 400876 542960 400904 543000
rect 408512 543000 408724 543028
rect 408512 542960 408540 543000
rect 400876 542932 408540 542960
rect 580258 542892 580264 542904
rect 369964 542864 580264 542892
rect 369765 542855 369823 542861
rect 580258 542852 580264 542864
rect 580316 542852 580322 542904
rect 355888 542796 369716 542824
rect 128357 542787 128415 542793
rect 449066 534012 449072 534064
rect 449124 534052 449130 534064
rect 579890 534052 579896 534064
rect 449124 534024 579896 534052
rect 449124 534012 449130 534024
rect 579890 534012 579896 534024
rect 579948 534012 579954 534064
rect 449802 510552 449808 510604
rect 449860 510592 449866 510604
rect 579890 510592 579896 510604
rect 449860 510564 579896 510592
rect 449860 510552 449866 510564
rect 579890 510552 579896 510564
rect 579948 510552 579954 510604
rect 2958 509940 2964 509992
rect 3016 509980 3022 509992
rect 6454 509980 6460 509992
rect 3016 509952 6460 509980
rect 3016 509940 3022 509952
rect 6454 509940 6460 509952
rect 6512 509940 6518 509992
rect 2774 495524 2780 495576
rect 2832 495564 2838 495576
rect 4706 495564 4712 495576
rect 2832 495536 4712 495564
rect 2832 495524 2838 495536
rect 4706 495524 4712 495536
rect 4764 495524 4770 495576
rect 449710 487092 449716 487144
rect 449768 487132 449774 487144
rect 580074 487132 580080 487144
rect 449768 487104 580080 487132
rect 449768 487092 449774 487104
rect 580074 487092 580080 487104
rect 580132 487092 580138 487144
rect 2774 481108 2780 481160
rect 2832 481148 2838 481160
rect 5442 481148 5448 481160
rect 2832 481120 5448 481148
rect 2832 481108 2838 481120
rect 5442 481108 5448 481120
rect 5500 481108 5506 481160
rect 449618 463632 449624 463684
rect 449676 463672 449682 463684
rect 580074 463672 580080 463684
rect 449676 463644 580080 463672
rect 449676 463632 449682 463644
rect 580074 463632 580080 463644
rect 580132 463632 580138 463684
rect 449526 452548 449532 452600
rect 449584 452588 449590 452600
rect 580074 452588 580080 452600
rect 449584 452560 580080 452588
rect 449584 452548 449590 452560
rect 580074 452548 580080 452560
rect 580132 452548 580138 452600
rect 2774 438540 2780 438592
rect 2832 438580 2838 438592
rect 5350 438580 5356 438592
rect 2832 438552 5356 438580
rect 2832 438540 2838 438552
rect 5350 438540 5356 438552
rect 5408 438540 5414 438592
rect 2774 424804 2780 424856
rect 2832 424844 2838 424856
rect 5258 424844 5264 424856
rect 2832 424816 5264 424844
rect 2832 424804 2838 424816
rect 5258 424804 5264 424816
rect 5316 424804 5322 424856
rect 449434 416712 449440 416764
rect 449492 416752 449498 416764
rect 580074 416752 580080 416764
rect 449492 416724 580080 416752
rect 449492 416712 449498 416724
rect 580074 416712 580080 416724
rect 580132 416712 580138 416764
rect 449342 405628 449348 405680
rect 449400 405668 449406 405680
rect 580074 405668 580080 405680
rect 449400 405640 580080 405668
rect 449400 405628 449406 405640
rect 580074 405628 580080 405640
rect 580132 405628 580138 405680
rect 2958 380604 2964 380656
rect 3016 380644 3022 380656
rect 6362 380644 6368 380656
rect 3016 380616 6368 380644
rect 3016 380604 3022 380616
rect 6362 380604 6368 380616
rect 6420 380604 6426 380656
rect 2774 366936 2780 366988
rect 2832 366976 2838 366988
rect 5166 366976 5172 366988
rect 2832 366948 5172 366976
rect 2832 366936 2838 366948
rect 5166 366936 5172 366948
rect 5224 366936 5230 366988
rect 3142 324096 3148 324148
rect 3200 324136 3206 324148
rect 6270 324136 6276 324148
rect 3200 324108 6276 324136
rect 3200 324096 3206 324108
rect 6270 324096 6276 324108
rect 6328 324096 6334 324148
rect 3142 280100 3148 280152
rect 3200 280140 3206 280152
rect 6178 280140 6184 280152
rect 3200 280112 6184 280140
rect 3200 280100 3206 280112
rect 6178 280100 6184 280112
rect 6236 280100 6242 280152
rect 2774 266160 2780 266212
rect 2832 266200 2838 266212
rect 5074 266200 5080 266212
rect 2832 266172 5080 266200
rect 2832 266160 2838 266172
rect 5074 266160 5080 266172
rect 5132 266160 5138 266212
rect 346946 243176 346952 243228
rect 347004 243216 347010 243228
rect 355413 243219 355471 243225
rect 355413 243216 355425 243219
rect 347004 243188 355425 243216
rect 347004 243176 347010 243188
rect 355413 243185 355425 243188
rect 355459 243185 355471 243219
rect 355413 243179 355471 243185
rect 183557 243083 183615 243089
rect 183557 243049 183569 243083
rect 183603 243080 183615 243083
rect 190641 243083 190699 243089
rect 190641 243080 190653 243083
rect 183603 243052 190653 243080
rect 183603 243049 183615 243052
rect 183557 243043 183615 243049
rect 190641 243049 190653 243052
rect 190687 243049 190699 243083
rect 190641 243043 190699 243049
rect 368934 243040 368940 243092
rect 368992 243080 368998 243092
rect 369762 243080 369768 243092
rect 368992 243052 369768 243080
rect 368992 243040 368998 243052
rect 369762 243040 369768 243052
rect 369820 243040 369826 243092
rect 184201 243015 184259 243021
rect 184201 242981 184213 243015
rect 184247 243012 184259 243015
rect 186866 243012 186872 243024
rect 184247 242984 186872 243012
rect 184247 242981 184259 242984
rect 184201 242975 184259 242981
rect 186866 242972 186872 242984
rect 186924 242972 186930 243024
rect 48317 242947 48375 242953
rect 48317 242913 48329 242947
rect 48363 242944 48375 242947
rect 57885 242947 57943 242953
rect 57885 242944 57897 242947
rect 48363 242916 57897 242944
rect 48363 242913 48375 242916
rect 48317 242907 48375 242913
rect 57885 242913 57897 242916
rect 57931 242913 57943 242947
rect 57885 242907 57943 242913
rect 67637 242947 67695 242953
rect 67637 242913 67649 242947
rect 67683 242944 67695 242947
rect 77205 242947 77263 242953
rect 77205 242944 77217 242947
rect 67683 242916 77217 242944
rect 67683 242913 67695 242916
rect 67637 242907 67695 242913
rect 77205 242913 77217 242916
rect 77251 242913 77263 242947
rect 77205 242907 77263 242913
rect 82081 242947 82139 242953
rect 82081 242913 82093 242947
rect 82127 242944 82139 242947
rect 86865 242947 86923 242953
rect 86865 242944 86877 242947
rect 82127 242916 86877 242944
rect 82127 242913 82139 242916
rect 82081 242907 82139 242913
rect 86865 242913 86877 242916
rect 86911 242913 86923 242947
rect 86865 242907 86923 242913
rect 132497 242947 132555 242953
rect 132497 242913 132509 242947
rect 132543 242944 132555 242947
rect 142249 242947 142307 242953
rect 142249 242944 142261 242947
rect 132543 242916 142261 242944
rect 132543 242913 132555 242916
rect 132497 242907 132555 242913
rect 142249 242913 142261 242916
rect 142295 242913 142307 242947
rect 142249 242907 142307 242913
rect 273165 242947 273223 242953
rect 273165 242913 273177 242947
rect 273211 242944 273223 242947
rect 342901 242947 342959 242953
rect 273211 242916 273392 242944
rect 273211 242913 273223 242916
rect 273165 242907 273223 242913
rect 71038 242836 71044 242888
rect 71096 242876 71102 242888
rect 169754 242876 169760 242888
rect 71096 242848 169760 242876
rect 71096 242836 71102 242848
rect 169754 242836 169760 242848
rect 169812 242836 169818 242888
rect 171781 242879 171839 242885
rect 171781 242845 171793 242879
rect 171827 242876 171839 242879
rect 178773 242879 178831 242885
rect 171827 242848 178724 242876
rect 171827 242845 171839 242848
rect 171781 242839 171839 242845
rect 42058 242768 42064 242820
rect 42116 242808 42122 242820
rect 48317 242811 48375 242817
rect 48317 242808 48329 242811
rect 42116 242780 48329 242808
rect 42116 242768 42122 242780
rect 48317 242777 48329 242780
rect 48363 242777 48375 242811
rect 67637 242811 67695 242817
rect 67637 242808 67649 242811
rect 48317 242771 48375 242777
rect 61948 242780 67649 242808
rect 57885 242743 57943 242749
rect 57885 242709 57897 242743
rect 57931 242740 57943 242743
rect 60645 242743 60703 242749
rect 60645 242740 60657 242743
rect 57931 242712 60657 242740
rect 57931 242709 57943 242712
rect 57885 242703 57943 242709
rect 60645 242709 60657 242712
rect 60691 242709 60703 242743
rect 60645 242703 60703 242709
rect 60737 242743 60795 242749
rect 60737 242709 60749 242743
rect 60783 242740 60795 242743
rect 61948 242740 61976 242780
rect 67637 242777 67649 242780
rect 67683 242777 67695 242811
rect 67637 242771 67695 242777
rect 89625 242811 89683 242817
rect 89625 242777 89637 242811
rect 89671 242808 89683 242811
rect 94501 242811 94559 242817
rect 94501 242808 94513 242811
rect 89671 242780 94513 242808
rect 89671 242777 89683 242780
rect 89625 242771 89683 242777
rect 94501 242777 94513 242780
rect 94547 242777 94559 242811
rect 94501 242771 94559 242777
rect 103422 242768 103428 242820
rect 103480 242808 103486 242820
rect 113177 242811 113235 242817
rect 113177 242808 113189 242811
rect 103480 242780 113189 242808
rect 103480 242768 103486 242780
rect 113177 242777 113189 242780
rect 113223 242777 113235 242811
rect 113177 242771 113235 242777
rect 122745 242811 122803 242817
rect 122745 242777 122757 242811
rect 122791 242808 122803 242811
rect 132497 242811 132555 242817
rect 132497 242808 132509 242811
rect 122791 242780 132509 242808
rect 122791 242777 122803 242780
rect 122745 242771 122803 242777
rect 132497 242777 132509 242780
rect 132543 242777 132555 242811
rect 132497 242771 132555 242777
rect 152461 242811 152519 242817
rect 152461 242777 152473 242811
rect 152507 242808 152519 242811
rect 162121 242811 162179 242817
rect 162121 242808 162133 242811
rect 152507 242780 162133 242808
rect 152507 242777 152519 242780
rect 152461 242771 152519 242777
rect 162121 242777 162133 242780
rect 162167 242777 162179 242811
rect 178696 242808 178724 242848
rect 178773 242845 178785 242879
rect 178819 242876 178831 242879
rect 190546 242876 190552 242888
rect 178819 242848 190552 242876
rect 178819 242845 178831 242848
rect 178773 242839 178831 242845
rect 190546 242836 190552 242848
rect 190604 242836 190610 242888
rect 190641 242879 190699 242885
rect 190641 242845 190653 242879
rect 190687 242876 190699 242879
rect 199654 242876 199660 242888
rect 190687 242848 199660 242876
rect 190687 242845 190699 242848
rect 190641 242839 190699 242845
rect 199654 242836 199660 242848
rect 199712 242836 199718 242888
rect 200761 242879 200819 242885
rect 200761 242845 200773 242879
rect 200807 242876 200819 242879
rect 210694 242876 210700 242888
rect 200807 242848 210700 242876
rect 200807 242845 200819 242848
rect 200761 242839 200819 242845
rect 210694 242836 210700 242848
rect 210752 242836 210758 242888
rect 211890 242836 211896 242888
rect 211948 242876 211954 242888
rect 254118 242876 254124 242888
rect 211948 242848 254124 242876
rect 211948 242836 211954 242848
rect 254118 242836 254124 242848
rect 254176 242836 254182 242888
rect 257982 242836 257988 242888
rect 258040 242876 258046 242888
rect 273364 242876 273392 242916
rect 342901 242913 342913 242947
rect 342947 242944 342959 242947
rect 347685 242947 347743 242953
rect 347685 242944 347697 242947
rect 342947 242916 347697 242944
rect 342947 242913 342959 242916
rect 342901 242907 342959 242913
rect 347685 242913 347697 242916
rect 347731 242913 347743 242947
rect 350813 242947 350871 242953
rect 350813 242944 350825 242947
rect 347685 242907 347743 242913
rect 350276 242916 350825 242944
rect 286502 242876 286508 242888
rect 258040 242848 273300 242876
rect 273364 242848 286508 242876
rect 258040 242836 258046 242848
rect 183370 242808 183376 242820
rect 178696 242780 183376 242808
rect 162121 242771 162179 242777
rect 183370 242768 183376 242780
rect 183428 242768 183434 242820
rect 183465 242811 183523 242817
rect 183465 242777 183477 242811
rect 183511 242777 183523 242811
rect 183465 242771 183523 242777
rect 220081 242811 220139 242817
rect 220081 242777 220093 242811
rect 220127 242808 220139 242811
rect 260190 242808 260196 242820
rect 220127 242780 260196 242808
rect 220127 242777 220139 242780
rect 220081 242771 220139 242777
rect 60783 242712 61976 242740
rect 77205 242743 77263 242749
rect 60783 242709 60795 242712
rect 60737 242703 60795 242709
rect 77205 242709 77217 242743
rect 77251 242740 77263 242743
rect 82081 242743 82139 242749
rect 82081 242740 82093 242743
rect 77251 242712 82093 242740
rect 77251 242709 77263 242712
rect 77205 242703 77263 242709
rect 82081 242709 82093 242712
rect 82127 242709 82139 242743
rect 82081 242703 82139 242709
rect 86218 242700 86224 242752
rect 86276 242740 86282 242752
rect 183281 242743 183339 242749
rect 183281 242740 183293 242743
rect 86276 242712 183293 242740
rect 86276 242700 86282 242712
rect 183281 242709 183293 242712
rect 183327 242709 183339 242743
rect 183480 242740 183508 242771
rect 260190 242768 260196 242780
rect 260248 242768 260254 242820
rect 261481 242811 261539 242817
rect 261481 242777 261493 242811
rect 261527 242808 261539 242811
rect 267550 242808 267556 242820
rect 261527 242780 267556 242808
rect 261527 242777 261539 242780
rect 261481 242771 261539 242777
rect 267550 242768 267556 242780
rect 267608 242768 267614 242820
rect 267645 242811 267703 242817
rect 267645 242777 267657 242811
rect 267691 242808 267703 242811
rect 273165 242811 273223 242817
rect 273165 242808 273177 242811
rect 267691 242780 273177 242808
rect 267691 242777 267703 242780
rect 267645 242771 267703 242777
rect 273165 242777 273177 242780
rect 273211 242777 273223 242811
rect 273272 242808 273300 242848
rect 286502 242836 286508 242848
rect 286560 242836 286566 242888
rect 312722 242836 312728 242888
rect 312780 242876 312786 242888
rect 316034 242876 316040 242888
rect 312780 242848 316040 242876
rect 312780 242836 312786 242848
rect 316034 242836 316040 242848
rect 316092 242836 316098 242888
rect 341426 242836 341432 242888
rect 341484 242876 341490 242888
rect 345937 242879 345995 242885
rect 345937 242876 345949 242879
rect 341484 242848 345949 242876
rect 341484 242836 341490 242848
rect 345937 242845 345949 242848
rect 345983 242845 345995 242879
rect 345937 242839 345995 242845
rect 346302 242836 346308 242888
rect 346360 242876 346366 242888
rect 350169 242879 350227 242885
rect 350169 242876 350181 242879
rect 346360 242848 350181 242876
rect 346360 242836 346366 242848
rect 350169 242845 350181 242848
rect 350215 242845 350227 242879
rect 350169 242839 350227 242845
rect 282178 242808 282184 242820
rect 273272 242780 282184 242808
rect 273165 242771 273223 242777
rect 282178 242768 282184 242780
rect 282236 242768 282242 242820
rect 284938 242768 284944 242820
rect 284996 242808 285002 242820
rect 288894 242808 288900 242820
rect 284996 242780 288900 242808
rect 284996 242768 285002 242780
rect 288894 242768 288900 242780
rect 288952 242768 288958 242820
rect 331674 242768 331680 242820
rect 331732 242808 331738 242820
rect 341518 242808 341524 242820
rect 331732 242780 341524 242808
rect 331732 242768 331738 242780
rect 341518 242768 341524 242780
rect 341576 242768 341582 242820
rect 345106 242768 345112 242820
rect 345164 242808 345170 242820
rect 350276 242808 350304 242916
rect 350813 242913 350825 242916
rect 350859 242913 350871 242947
rect 350813 242907 350871 242913
rect 367738 242904 367744 242956
rect 367796 242944 367802 242956
rect 369949 242947 370007 242953
rect 369949 242944 369961 242947
rect 367796 242916 369961 242944
rect 367796 242904 367802 242916
rect 369949 242913 369961 242916
rect 369995 242913 370007 242947
rect 369949 242907 370007 242913
rect 414474 242904 414480 242956
rect 414532 242944 414538 242956
rect 418157 242947 418215 242953
rect 418157 242944 418169 242947
rect 414532 242916 418169 242944
rect 414532 242904 414538 242916
rect 418157 242913 418169 242916
rect 418203 242913 418215 242947
rect 418157 242907 418215 242913
rect 350353 242879 350411 242885
rect 350353 242845 350365 242879
rect 350399 242876 350411 242879
rect 377398 242876 377404 242888
rect 350399 242848 377404 242876
rect 350399 242845 350411 242848
rect 350353 242839 350411 242845
rect 377398 242836 377404 242848
rect 377456 242836 377462 242888
rect 379517 242879 379575 242885
rect 379517 242845 379529 242879
rect 379563 242876 379575 242879
rect 398098 242876 398104 242888
rect 379563 242848 398104 242876
rect 379563 242845 379575 242848
rect 379517 242839 379575 242845
rect 398098 242836 398104 242848
rect 398156 242836 398162 242888
rect 399478 242836 399484 242888
rect 399536 242876 399542 242888
rect 485774 242876 485780 242888
rect 399536 242848 485780 242876
rect 399536 242836 399542 242848
rect 485774 242836 485780 242848
rect 485832 242836 485838 242888
rect 345164 242780 350304 242808
rect 350445 242811 350503 242817
rect 345164 242768 345170 242780
rect 350445 242777 350457 242811
rect 350491 242808 350503 242811
rect 364613 242811 364671 242817
rect 364613 242808 364625 242811
rect 350491 242780 364625 242808
rect 350491 242777 350503 242780
rect 350445 242771 350503 242777
rect 364613 242777 364625 242780
rect 364659 242777 364671 242811
rect 364613 242771 364671 242777
rect 364702 242768 364708 242820
rect 364760 242808 364766 242820
rect 370041 242811 370099 242817
rect 370041 242808 370053 242811
rect 364760 242780 370053 242808
rect 364760 242768 364766 242780
rect 370041 242777 370053 242780
rect 370087 242777 370099 242811
rect 370041 242771 370099 242777
rect 370130 242768 370136 242820
rect 370188 242808 370194 242820
rect 371142 242808 371148 242820
rect 370188 242780 371148 242808
rect 370188 242768 370194 242780
rect 371142 242768 371148 242780
rect 371200 242768 371206 242820
rect 375650 242768 375656 242820
rect 375708 242808 375714 242820
rect 439038 242808 439044 242820
rect 375708 242780 439044 242808
rect 375708 242768 375714 242780
rect 439038 242768 439044 242780
rect 439096 242768 439102 242820
rect 443454 242768 443460 242820
rect 443512 242808 443518 242820
rect 449989 242811 450047 242817
rect 449989 242808 450001 242811
rect 443512 242780 450001 242808
rect 443512 242768 443518 242780
rect 449989 242777 450001 242780
rect 450035 242777 450047 242811
rect 449989 242771 450047 242777
rect 184201 242743 184259 242749
rect 184201 242740 184213 242743
rect 183480 242712 184213 242740
rect 183281 242703 183339 242709
rect 184201 242709 184213 242712
rect 184247 242709 184259 242743
rect 184201 242703 184259 242709
rect 199378 242700 199384 242752
rect 199436 242740 199442 242752
rect 245562 242740 245568 242752
rect 199436 242712 245568 242740
rect 199436 242700 199442 242712
rect 245562 242700 245568 242712
rect 245620 242700 245626 242752
rect 245654 242700 245660 242752
rect 245712 242740 245718 242752
rect 271325 242743 271383 242749
rect 271325 242740 271337 242743
rect 245712 242712 271337 242740
rect 245712 242700 245718 242712
rect 271325 242709 271337 242712
rect 271371 242709 271383 242743
rect 271325 242703 271383 242709
rect 276753 242743 276811 242749
rect 276753 242709 276765 242743
rect 276799 242740 276811 242743
rect 280338 242740 280344 242752
rect 276799 242712 280344 242740
rect 276799 242709 276811 242712
rect 276753 242703 276811 242709
rect 280338 242700 280344 242712
rect 280396 242700 280402 242752
rect 294782 242700 294788 242752
rect 294840 242740 294846 242752
rect 296806 242740 296812 242752
rect 294840 242712 296812 242740
rect 294840 242700 294846 242712
rect 296806 242700 296812 242712
rect 296864 242700 296870 242752
rect 314562 242700 314568 242752
rect 314620 242740 314626 242752
rect 316770 242740 316776 242752
rect 314620 242712 316776 242740
rect 314620 242700 314626 242712
rect 316770 242700 316776 242712
rect 316828 242700 316834 242752
rect 329834 242700 329840 242752
rect 329892 242740 329898 242752
rect 340138 242740 340144 242752
rect 329892 242712 340144 242740
rect 329892 242700 329898 242712
rect 340138 242700 340144 242712
rect 340196 242700 340202 242752
rect 343266 242700 343272 242752
rect 343324 242740 343330 242752
rect 350353 242743 350411 242749
rect 350353 242740 350365 242743
rect 343324 242712 350365 242740
rect 343324 242700 343330 242712
rect 350353 242709 350365 242712
rect 350399 242709 350411 242743
rect 367189 242743 367247 242749
rect 367189 242740 367201 242743
rect 350353 242703 350411 242709
rect 350460 242712 367201 242740
rect 88978 242632 88984 242684
rect 89036 242672 89042 242684
rect 178773 242675 178831 242681
rect 178773 242672 178785 242675
rect 89036 242644 178785 242672
rect 89036 242632 89042 242644
rect 178773 242641 178785 242644
rect 178819 242641 178831 242675
rect 178773 242635 178831 242641
rect 183462 242632 183468 242684
rect 183520 242672 183526 242684
rect 183557 242675 183615 242681
rect 183557 242672 183569 242675
rect 183520 242644 183569 242672
rect 183520 242632 183526 242644
rect 183557 242641 183569 242644
rect 183603 242641 183615 242675
rect 183557 242635 183615 242641
rect 188338 242632 188344 242684
rect 188396 242672 188402 242684
rect 200761 242675 200819 242681
rect 200761 242672 200773 242675
rect 188396 242644 200773 242672
rect 188396 242632 188402 242644
rect 200761 242641 200773 242644
rect 200807 242641 200819 242675
rect 200761 242635 200819 242641
rect 211798 242632 211804 242684
rect 211856 242672 211862 242684
rect 258350 242672 258356 242684
rect 211856 242644 258356 242672
rect 211856 242632 211862 242644
rect 258350 242632 258356 242644
rect 258408 242632 258414 242684
rect 259362 242632 259368 242684
rect 259420 242672 259426 242684
rect 282822 242672 282828 242684
rect 259420 242644 282828 242672
rect 259420 242632 259426 242644
rect 282822 242632 282828 242644
rect 282880 242632 282886 242684
rect 286318 242632 286324 242684
rect 286376 242672 286382 242684
rect 292574 242672 292580 242684
rect 286376 242644 292580 242672
rect 286376 242632 286382 242644
rect 292574 242632 292580 242644
rect 292632 242632 292638 242684
rect 313918 242632 313924 242684
rect 313976 242672 313982 242684
rect 319070 242672 319076 242684
rect 313976 242644 319076 242672
rect 313976 242632 313982 242644
rect 319070 242632 319076 242644
rect 319128 242632 319134 242684
rect 328638 242632 328644 242684
rect 328696 242672 328702 242684
rect 341981 242675 342039 242681
rect 341981 242672 341993 242675
rect 328696 242644 341993 242672
rect 328696 242632 328702 242644
rect 341981 242641 341993 242644
rect 342027 242641 342039 242675
rect 341981 242635 342039 242641
rect 342070 242632 342076 242684
rect 342128 242672 342134 242684
rect 350460 242672 350488 242712
rect 367189 242709 367201 242712
rect 367235 242709 367247 242743
rect 367189 242703 367247 242709
rect 378134 242700 378140 242752
rect 378192 242740 378198 242752
rect 379422 242740 379428 242752
rect 378192 242712 379428 242740
rect 378192 242700 378198 242712
rect 379422 242700 379428 242712
rect 379480 242700 379486 242752
rect 379517 242743 379575 242749
rect 379517 242709 379529 242743
rect 379563 242709 379575 242743
rect 379517 242703 379575 242709
rect 342128 242644 350488 242672
rect 350537 242675 350595 242681
rect 342128 242632 342134 242644
rect 350537 242641 350549 242675
rect 350583 242641 350595 242675
rect 350537 242635 350595 242641
rect 93118 242564 93124 242616
rect 93176 242604 93182 242616
rect 196066 242604 196072 242616
rect 93176 242576 196072 242604
rect 93176 242564 93182 242576
rect 196066 242564 196072 242576
rect 196124 242564 196130 242616
rect 208302 242564 208308 242616
rect 208360 242604 208366 242616
rect 256510 242604 256516 242616
rect 208360 242576 256516 242604
rect 208360 242564 208366 242576
rect 256510 242564 256516 242576
rect 256568 242564 256574 242616
rect 262030 242604 262036 242616
rect 256620 242576 262036 242604
rect 86865 242539 86923 242545
rect 86865 242505 86877 242539
rect 86911 242536 86923 242539
rect 89625 242539 89683 242545
rect 89625 242536 89637 242539
rect 86911 242508 89637 242536
rect 86911 242505 86923 242508
rect 86865 242499 86923 242505
rect 89625 242505 89637 242508
rect 89671 242505 89683 242539
rect 89625 242499 89683 242505
rect 94501 242539 94559 242545
rect 94501 242505 94513 242539
rect 94547 242536 94559 242539
rect 103517 242539 103575 242545
rect 103517 242536 103529 242539
rect 94547 242508 103529 242536
rect 94547 242505 94559 242508
rect 94501 242499 94559 242505
rect 103517 242505 103529 242508
rect 103563 242505 103575 242539
rect 103517 242499 103575 242505
rect 113085 242539 113143 242545
rect 113085 242505 113097 242539
rect 113131 242536 113143 242539
rect 113174 242536 113180 242548
rect 113131 242508 113180 242536
rect 113131 242505 113143 242508
rect 113085 242499 113143 242505
rect 113174 242496 113180 242508
rect 113232 242496 113238 242548
rect 122742 242496 122748 242548
rect 122800 242536 122806 242548
rect 142157 242539 142215 242545
rect 142157 242536 142169 242539
rect 122800 242508 142169 242536
rect 122800 242496 122806 242508
rect 142157 242505 142169 242508
rect 142203 242505 142215 242539
rect 142157 242499 142215 242505
rect 142249 242539 142307 242545
rect 142249 242505 142261 242539
rect 142295 242536 142307 242539
rect 152461 242539 152519 242545
rect 152461 242536 152473 242539
rect 142295 242508 152473 242536
rect 142295 242505 142307 242508
rect 142249 242499 142307 242505
rect 152461 242505 152473 242508
rect 152507 242505 152519 242539
rect 152461 242499 152519 242505
rect 152553 242539 152611 242545
rect 152553 242505 152565 242539
rect 152599 242536 152611 242539
rect 170398 242536 170404 242548
rect 152599 242508 170404 242536
rect 152599 242505 152611 242508
rect 152553 242499 152611 242505
rect 170398 242496 170404 242508
rect 170456 242496 170462 242548
rect 180058 242496 180064 242548
rect 180116 242536 180122 242548
rect 188706 242536 188712 242548
rect 180116 242508 188712 242536
rect 180116 242496 180122 242508
rect 188706 242496 188712 242508
rect 188764 242496 188770 242548
rect 203610 242496 203616 242548
rect 203668 242536 203674 242548
rect 252278 242536 252284 242548
rect 203668 242508 252284 242536
rect 203668 242496 203674 242508
rect 252278 242496 252284 242508
rect 252336 242496 252342 242548
rect 254578 242496 254584 242548
rect 254636 242536 254642 242548
rect 256620 242536 256648 242576
rect 262030 242564 262036 242576
rect 262088 242564 262094 242616
rect 266262 242564 266268 242616
rect 266320 242604 266326 242616
rect 267645 242607 267703 242613
rect 267645 242604 267657 242607
rect 266320 242576 267657 242604
rect 266320 242564 266326 242576
rect 267645 242573 267657 242576
rect 267691 242573 267703 242607
rect 267645 242567 267703 242573
rect 268289 242607 268347 242613
rect 268289 242573 268301 242607
rect 268335 242604 268347 242607
rect 284662 242604 284668 242616
rect 268335 242576 284668 242604
rect 268335 242573 268347 242576
rect 268289 242567 268347 242573
rect 284662 242564 284668 242576
rect 284720 242564 284726 242616
rect 313366 242564 313372 242616
rect 313424 242604 313430 242616
rect 316678 242604 316684 242616
rect 313424 242576 316684 242604
rect 313424 242564 313430 242576
rect 316678 242564 316684 242576
rect 316736 242564 316742 242616
rect 325602 242564 325608 242616
rect 325660 242604 325666 242616
rect 338758 242604 338764 242616
rect 325660 242576 338764 242604
rect 325660 242564 325666 242576
rect 338758 242564 338764 242576
rect 338816 242564 338822 242616
rect 347685 242607 347743 242613
rect 347685 242573 347697 242607
rect 347731 242604 347743 242607
rect 350552 242604 350580 242635
rect 351822 242632 351828 242684
rect 351880 242672 351886 242684
rect 367094 242672 367100 242684
rect 351880 242644 367100 242672
rect 351880 242632 351886 242644
rect 367094 242632 367100 242644
rect 367152 242632 367158 242684
rect 367281 242675 367339 242681
rect 367281 242641 367293 242675
rect 367327 242672 367339 242675
rect 367646 242672 367652 242684
rect 367327 242644 367652 242672
rect 367327 242641 367339 242644
rect 367281 242635 367339 242641
rect 367646 242632 367652 242644
rect 367704 242632 367710 242684
rect 376938 242632 376944 242684
rect 376996 242672 377002 242684
rect 379532 242672 379560 242703
rect 404998 242700 405004 242752
rect 405056 242740 405062 242752
rect 435358 242740 435364 242752
rect 405056 242712 435364 242740
rect 405056 242700 405062 242712
rect 435358 242700 435364 242712
rect 435416 242700 435422 242752
rect 436186 242700 436192 242752
rect 436244 242740 436250 242752
rect 525058 242740 525064 242752
rect 436244 242712 525064 242740
rect 436244 242700 436250 242712
rect 525058 242700 525064 242712
rect 525116 242700 525122 242752
rect 376996 242644 379560 242672
rect 379609 242675 379667 242681
rect 376996 242632 377002 242644
rect 379609 242641 379621 242675
rect 379655 242672 379667 242675
rect 385678 242672 385684 242684
rect 379655 242644 385684 242672
rect 379655 242641 379667 242644
rect 379609 242635 379667 242641
rect 385678 242632 385684 242644
rect 385736 242632 385742 242684
rect 403158 242632 403164 242684
rect 403216 242672 403222 242684
rect 492674 242672 492680 242684
rect 403216 242644 492680 242672
rect 403216 242632 403222 242644
rect 492674 242632 492680 242644
rect 492732 242632 492738 242684
rect 347731 242576 350580 242604
rect 350813 242607 350871 242613
rect 347731 242573 347743 242576
rect 347685 242567 347743 242573
rect 350813 242573 350825 242607
rect 350859 242604 350871 242607
rect 367189 242607 367247 242613
rect 367189 242604 367201 242607
rect 350859 242576 367201 242604
rect 350859 242573 350871 242576
rect 350813 242567 350871 242573
rect 367189 242573 367201 242576
rect 367235 242573 367247 242607
rect 367189 242567 367247 242573
rect 367373 242607 367431 242613
rect 367373 242573 367385 242607
rect 367419 242604 367431 242607
rect 379698 242604 379704 242616
rect 367419 242576 379704 242604
rect 367419 242573 367431 242576
rect 367373 242567 367431 242573
rect 379698 242564 379704 242576
rect 379756 242564 379762 242616
rect 401318 242564 401324 242616
rect 401376 242604 401382 242616
rect 422941 242607 422999 242613
rect 422941 242604 422953 242607
rect 401376 242576 422953 242604
rect 401376 242564 401382 242576
rect 422941 242573 422953 242576
rect 422987 242573 422999 242607
rect 422941 242567 422999 242573
rect 425146 242564 425152 242616
rect 425204 242604 425210 242616
rect 431865 242607 431923 242613
rect 431865 242604 431877 242607
rect 425204 242576 431877 242604
rect 425204 242564 425210 242576
rect 431865 242573 431877 242576
rect 431911 242573 431923 242607
rect 431865 242567 431923 242573
rect 432506 242564 432512 242616
rect 432564 242604 432570 242616
rect 523678 242604 523684 242616
rect 432564 242576 523684 242604
rect 432564 242564 432570 242576
rect 523678 242564 523684 242576
rect 523736 242564 523742 242616
rect 254636 242508 256648 242536
rect 254636 242496 254642 242508
rect 256694 242496 256700 242548
rect 256752 242536 256758 242548
rect 281534 242536 281540 242548
rect 256752 242508 281540 242536
rect 256752 242496 256758 242508
rect 281534 242496 281540 242508
rect 281592 242496 281598 242548
rect 288250 242496 288256 242548
rect 288308 242536 288314 242548
rect 297450 242536 297456 242548
rect 288308 242508 297456 242536
rect 288308 242496 288314 242508
rect 297450 242496 297456 242508
rect 297508 242496 297514 242548
rect 333514 242496 333520 242548
rect 333572 242536 333578 242548
rect 342901 242539 342959 242545
rect 342901 242536 342913 242539
rect 333572 242508 342913 242536
rect 333572 242496 333578 242508
rect 342901 242505 342913 242508
rect 342947 242505 342959 242539
rect 342901 242499 342959 242505
rect 345661 242539 345719 242545
rect 345661 242505 345673 242539
rect 345707 242536 345719 242539
rect 350537 242539 350595 242545
rect 350537 242536 350549 242539
rect 345707 242508 350549 242536
rect 345707 242505 345719 242508
rect 345661 242499 345719 242505
rect 350537 242505 350549 242508
rect 350583 242505 350595 242539
rect 350537 242499 350595 242505
rect 350629 242539 350687 242545
rect 350629 242505 350641 242539
rect 350675 242536 350687 242539
rect 350675 242508 355364 242536
rect 350675 242505 350687 242508
rect 350629 242499 350687 242505
rect 35158 242428 35164 242480
rect 35216 242468 35222 242480
rect 166718 242468 166724 242480
rect 35216 242440 166724 242468
rect 35216 242428 35222 242440
rect 166718 242428 166724 242440
rect 166776 242428 166782 242480
rect 176102 242428 176108 242480
rect 176160 242468 176166 242480
rect 181346 242468 181352 242480
rect 176160 242440 181352 242468
rect 176160 242428 176166 242440
rect 181346 242428 181352 242440
rect 181404 242428 181410 242480
rect 184198 242428 184204 242480
rect 184256 242468 184262 242480
rect 194226 242468 194232 242480
rect 184256 242440 194232 242468
rect 184256 242428 184262 242440
rect 194226 242428 194232 242440
rect 194284 242428 194290 242480
rect 198274 242428 198280 242480
rect 198332 242468 198338 242480
rect 247402 242468 247408 242480
rect 198332 242440 247408 242468
rect 198332 242428 198338 242440
rect 247402 242428 247408 242440
rect 247460 242428 247466 242480
rect 248322 242428 248328 242480
rect 248380 242468 248386 242480
rect 277302 242468 277308 242480
rect 248380 242440 277308 242468
rect 248380 242428 248386 242440
rect 277302 242428 277308 242440
rect 277360 242428 277366 242480
rect 277394 242428 277400 242480
rect 277452 242468 277458 242480
rect 291930 242468 291936 242480
rect 277452 242440 291936 242468
rect 277452 242428 277458 242440
rect 291930 242428 291936 242440
rect 291988 242428 291994 242480
rect 292482 242428 292488 242480
rect 292540 242468 292546 242480
rect 299934 242468 299940 242480
rect 292540 242440 299940 242468
rect 292540 242428 292546 242440
rect 299934 242428 299940 242440
rect 299992 242428 299998 242480
rect 341981 242471 342039 242477
rect 341981 242437 341993 242471
rect 342027 242468 342039 242471
rect 347958 242468 347964 242480
rect 342027 242440 347964 242468
rect 342027 242437 342039 242440
rect 341981 242431 342039 242437
rect 347958 242428 347964 242440
rect 348016 242428 348022 242480
rect 349982 242428 349988 242480
rect 350040 242468 350046 242480
rect 355229 242471 355287 242477
rect 355229 242468 355241 242471
rect 350040 242440 355241 242468
rect 350040 242428 350046 242440
rect 355229 242437 355241 242440
rect 355275 242437 355287 242471
rect 355336 242468 355364 242508
rect 357342 242496 357348 242548
rect 357400 242536 357406 242548
rect 367094 242536 367100 242548
rect 357400 242508 367100 242536
rect 357400 242496 357406 242508
rect 367094 242496 367100 242508
rect 367152 242496 367158 242548
rect 367462 242496 367468 242548
rect 367520 242536 367526 242548
rect 391198 242536 391204 242548
rect 367520 242508 391204 242536
rect 367520 242496 367526 242508
rect 391198 242496 391204 242508
rect 391256 242496 391262 242548
rect 397638 242496 397644 242548
rect 397696 242536 397702 242548
rect 403618 242536 403624 242548
rect 397696 242508 403624 242536
rect 397696 242496 397702 242508
rect 403618 242496 403624 242508
rect 403676 242496 403682 242548
rect 414017 242539 414075 242545
rect 414017 242505 414029 242539
rect 414063 242536 414075 242539
rect 502978 242536 502984 242548
rect 414063 242508 502984 242536
rect 414063 242505 414075 242508
rect 414017 242499 414075 242505
rect 502978 242496 502984 242508
rect 503036 242496 503042 242548
rect 359458 242468 359464 242480
rect 355336 242440 359464 242468
rect 355229 242431 355287 242437
rect 359458 242428 359464 242440
rect 359516 242428 359522 242480
rect 361850 242468 361856 242480
rect 359660 242440 361856 242468
rect 31018 242360 31024 242412
rect 31076 242400 31082 242412
rect 163038 242400 163044 242412
rect 31076 242372 163044 242400
rect 31076 242360 31082 242372
rect 163038 242360 163044 242372
rect 163096 242360 163102 242412
rect 187142 242360 187148 242412
rect 187200 242400 187206 242412
rect 201494 242400 201500 242412
rect 187200 242372 201500 242400
rect 187200 242360 187206 242372
rect 201494 242360 201500 242372
rect 201552 242360 201558 242412
rect 204162 242360 204168 242412
rect 204220 242400 204226 242412
rect 254670 242400 254676 242412
rect 204220 242372 254676 242400
rect 204220 242360 204226 242372
rect 254670 242360 254676 242372
rect 254728 242360 254734 242412
rect 255222 242360 255228 242412
rect 255280 242400 255286 242412
rect 280982 242400 280988 242412
rect 255280 242372 280988 242400
rect 255280 242360 255286 242372
rect 280982 242360 280988 242372
rect 281040 242360 281046 242412
rect 288342 242360 288348 242412
rect 288400 242400 288406 242412
rect 298094 242400 298100 242412
rect 288400 242372 298100 242400
rect 288400 242360 288406 242372
rect 298094 242360 298100 242372
rect 298152 242360 298158 242412
rect 326798 242360 326804 242412
rect 326856 242400 326862 242412
rect 342898 242400 342904 242412
rect 326856 242372 342904 242400
rect 326856 242360 326862 242372
rect 342898 242360 342904 242372
rect 342956 242360 342962 242412
rect 24118 242292 24124 242344
rect 24176 242332 24182 242344
rect 158162 242332 158168 242344
rect 24176 242304 158168 242332
rect 24176 242292 24182 242304
rect 158162 242292 158168 242304
rect 158220 242292 158226 242344
rect 162121 242335 162179 242341
rect 162121 242301 162133 242335
rect 162167 242332 162179 242335
rect 171781 242335 171839 242341
rect 171781 242332 171793 242335
rect 162167 242304 171793 242332
rect 162167 242301 162179 242304
rect 162121 242295 162179 242301
rect 171781 242301 171793 242304
rect 171827 242301 171839 242335
rect 171781 242295 171839 242301
rect 185578 242292 185584 242344
rect 185636 242332 185642 242344
rect 197906 242332 197912 242344
rect 185636 242304 197912 242332
rect 185636 242292 185642 242304
rect 197906 242292 197912 242304
rect 197964 242292 197970 242344
rect 198182 242292 198188 242344
rect 198240 242332 198246 242344
rect 238481 242335 238539 242341
rect 238481 242332 238493 242335
rect 198240 242304 238493 242332
rect 198240 242292 198246 242304
rect 238481 242301 238493 242304
rect 238527 242301 238539 242335
rect 238481 242295 238539 242301
rect 249702 242292 249708 242344
rect 249760 242332 249766 242344
rect 277946 242332 277952 242344
rect 249760 242304 277952 242332
rect 249760 242292 249766 242304
rect 277946 242292 277952 242304
rect 278004 242292 278010 242344
rect 284202 242292 284208 242344
rect 284260 242332 284266 242344
rect 295610 242332 295616 242344
rect 284260 242304 295616 242332
rect 284260 242292 284266 242304
rect 295610 242292 295616 242304
rect 295668 242292 295674 242344
rect 315206 242292 315212 242344
rect 315264 242332 315270 242344
rect 321646 242332 321652 242344
rect 315264 242304 321652 242332
rect 315264 242292 315270 242304
rect 321646 242292 321652 242304
rect 321704 242292 321710 242344
rect 324958 242292 324964 242344
rect 325016 242332 325022 242344
rect 330478 242332 330484 242344
rect 325016 242304 330484 242332
rect 325016 242292 325022 242304
rect 330478 242292 330484 242304
rect 330536 242292 330542 242344
rect 335998 242292 336004 242344
rect 336056 242332 336062 242344
rect 355226 242332 355232 242344
rect 336056 242304 355232 242332
rect 336056 242292 336062 242304
rect 355226 242292 355232 242304
rect 355284 242292 355290 242344
rect 355502 242292 355508 242344
rect 355560 242332 355566 242344
rect 359660 242332 359688 242440
rect 361850 242428 361856 242440
rect 361908 242428 361914 242480
rect 364613 242471 364671 242477
rect 364613 242437 364625 242471
rect 364659 242468 364671 242471
rect 367189 242471 367247 242477
rect 367189 242468 367201 242471
rect 364659 242440 367201 242468
rect 364659 242437 364671 242440
rect 364613 242431 364671 242437
rect 367189 242437 367201 242440
rect 367235 242437 367247 242471
rect 367189 242431 367247 242437
rect 369213 242471 369271 242477
rect 369213 242437 369225 242471
rect 369259 242468 369271 242471
rect 395338 242468 395344 242480
rect 369259 242440 395344 242468
rect 369259 242437 369271 242440
rect 369213 242431 369271 242437
rect 395338 242428 395344 242440
rect 395396 242428 395402 242480
rect 397086 242428 397092 242480
rect 397144 242468 397150 242480
rect 412729 242471 412787 242477
rect 412729 242468 412741 242471
rect 397144 242440 412741 242468
rect 397144 242428 397150 242440
rect 412729 242437 412741 242440
rect 412775 242437 412787 242471
rect 412729 242431 412787 242437
rect 412913 242471 412971 242477
rect 412913 242437 412925 242471
rect 412959 242468 412971 242471
rect 421558 242468 421564 242480
rect 412959 242440 421564 242468
rect 412959 242437 412971 242440
rect 412913 242431 412971 242437
rect 421558 242428 421564 242440
rect 421616 242428 421622 242480
rect 422941 242471 422999 242477
rect 422941 242437 422953 242471
rect 422987 242468 422999 242471
rect 431218 242468 431224 242480
rect 422987 242440 431224 242468
rect 422987 242437 422999 242440
rect 422941 242431 422999 242437
rect 431218 242428 431224 242440
rect 431276 242428 431282 242480
rect 431957 242471 432015 242477
rect 431957 242437 431969 242471
rect 432003 242468 432015 242471
rect 518158 242468 518164 242480
rect 432003 242440 518164 242468
rect 432003 242437 432015 242440
rect 431957 242431 432015 242437
rect 518158 242428 518164 242440
rect 518216 242428 518222 242480
rect 369578 242360 369584 242412
rect 369636 242400 369642 242412
rect 382458 242400 382464 242412
rect 369636 242372 382464 242400
rect 369636 242360 369642 242372
rect 382458 242360 382464 242372
rect 382516 242360 382522 242412
rect 389726 242360 389732 242412
rect 389784 242400 389790 242412
rect 394237 242403 394295 242409
rect 394237 242400 394249 242403
rect 389784 242372 394249 242400
rect 389784 242360 389790 242372
rect 394237 242369 394249 242372
rect 394283 242369 394295 242403
rect 394237 242363 394295 242369
rect 395246 242360 395252 242412
rect 395304 242400 395310 242412
rect 420178 242400 420184 242412
rect 395304 242372 420184 242400
rect 395304 242360 395310 242372
rect 420178 242360 420184 242372
rect 420236 242360 420242 242412
rect 421466 242360 421472 242412
rect 421524 242400 421530 242412
rect 514018 242400 514024 242412
rect 421524 242372 514024 242400
rect 421524 242360 421530 242372
rect 514018 242360 514024 242372
rect 514076 242360 514082 242412
rect 355560 242304 359688 242332
rect 355560 242292 355566 242304
rect 361022 242292 361028 242344
rect 361080 242332 361086 242344
rect 369213 242335 369271 242341
rect 369213 242332 369225 242335
rect 361080 242304 369225 242332
rect 361080 242292 361086 242304
rect 369213 242301 369225 242304
rect 369259 242301 369271 242335
rect 369213 242295 369271 242301
rect 370041 242335 370099 242341
rect 370041 242301 370053 242335
rect 370087 242332 370099 242335
rect 409138 242332 409144 242344
rect 370087 242304 409144 242332
rect 370087 242301 370099 242304
rect 370041 242295 370099 242301
rect 409138 242292 409144 242304
rect 409196 242292 409202 242344
rect 410518 242292 410524 242344
rect 410576 242332 410582 242344
rect 414017 242335 414075 242341
rect 414017 242332 414029 242335
rect 410576 242304 414029 242332
rect 410576 242292 410582 242304
rect 414017 242301 414029 242304
rect 414063 242301 414075 242335
rect 414017 242295 414075 242301
rect 416038 242292 416044 242344
rect 416096 242332 416102 242344
rect 416682 242332 416688 242344
rect 416096 242304 416688 242332
rect 416096 242292 416102 242304
rect 416682 242292 416688 242304
rect 416740 242292 416746 242344
rect 418157 242335 418215 242341
rect 418157 242301 418169 242335
rect 418203 242332 418215 242335
rect 507118 242332 507124 242344
rect 418203 242304 507124 242332
rect 418203 242301 418215 242304
rect 418157 242295 418215 242301
rect 507118 242292 507124 242304
rect 507176 242292 507182 242344
rect 28258 242224 28264 242276
rect 28316 242264 28322 242276
rect 162394 242264 162400 242276
rect 28316 242236 162400 242264
rect 28316 242224 28322 242236
rect 162394 242224 162400 242236
rect 162452 242224 162458 242276
rect 163498 242224 163504 242276
rect 163556 242264 163562 242276
rect 200942 242264 200948 242276
rect 163556 242236 200948 242264
rect 163556 242224 163562 242236
rect 200942 242224 200948 242236
rect 201000 242224 201006 242276
rect 201402 242224 201408 242276
rect 201460 242264 201466 242276
rect 252830 242264 252836 242276
rect 201460 242236 252836 242264
rect 201460 242224 201466 242236
rect 252830 242224 252836 242236
rect 252888 242224 252894 242276
rect 254670 242224 254676 242276
rect 254728 242264 254734 242276
rect 276753 242267 276811 242273
rect 276753 242264 276765 242267
rect 254728 242236 276765 242264
rect 254728 242224 254734 242236
rect 276753 242233 276765 242236
rect 276799 242233 276811 242267
rect 276753 242227 276811 242233
rect 281442 242224 281448 242276
rect 281500 242264 281506 242276
rect 294414 242264 294420 242276
rect 281500 242236 294420 242264
rect 281500 242224 281506 242236
rect 294414 242224 294420 242236
rect 294472 242224 294478 242276
rect 317598 242224 317604 242276
rect 317656 242264 317662 242276
rect 325786 242264 325792 242276
rect 317656 242236 325792 242264
rect 317656 242224 317662 242236
rect 325786 242224 325792 242236
rect 325844 242224 325850 242276
rect 337746 242224 337752 242276
rect 337804 242264 337810 242276
rect 355321 242267 355379 242273
rect 355321 242264 355333 242267
rect 337804 242236 355333 242264
rect 337804 242224 337810 242236
rect 355321 242233 355333 242236
rect 355367 242233 355379 242267
rect 355321 242227 355379 242233
rect 355413 242267 355471 242273
rect 355413 242233 355425 242267
rect 355459 242264 355471 242267
rect 357434 242264 357440 242276
rect 355459 242236 357440 242264
rect 355459 242233 355471 242236
rect 355413 242227 355471 242233
rect 357434 242224 357440 242236
rect 357492 242224 357498 242276
rect 368382 242224 368388 242276
rect 368440 242264 368446 242276
rect 411254 242264 411260 242276
rect 368440 242236 411260 242264
rect 368440 242224 368446 242236
rect 411254 242224 411260 242236
rect 411312 242224 411318 242276
rect 411714 242224 411720 242276
rect 411772 242264 411778 242276
rect 412542 242264 412548 242276
rect 411772 242236 412548 242264
rect 411772 242224 411778 242236
rect 412542 242224 412548 242236
rect 412600 242224 412606 242276
rect 412821 242267 412879 242273
rect 412821 242233 412833 242267
rect 412867 242264 412879 242267
rect 418249 242267 418307 242273
rect 418249 242264 418261 242267
rect 412867 242236 418261 242264
rect 412867 242233 412879 242236
rect 412821 242227 412879 242233
rect 418249 242233 418261 242236
rect 418295 242233 418307 242267
rect 418249 242227 418307 242233
rect 418341 242267 418399 242273
rect 418341 242233 418353 242267
rect 418387 242264 418399 242267
rect 422938 242264 422944 242276
rect 418387 242236 422944 242264
rect 418387 242233 418399 242236
rect 418341 242227 418399 242233
rect 422938 242224 422944 242236
rect 422996 242224 423002 242276
rect 428826 242224 428832 242276
rect 428884 242264 428890 242276
rect 520918 242264 520924 242276
rect 428884 242236 520924 242264
rect 428884 242224 428890 242236
rect 520918 242224 520924 242236
rect 520976 242224 520982 242276
rect 17218 242156 17224 242208
rect 17276 242196 17282 242208
rect 157518 242196 157524 242208
rect 17276 242168 157524 242196
rect 17276 242156 17282 242168
rect 157518 242156 157524 242168
rect 157576 242156 157582 242208
rect 181622 242156 181628 242208
rect 181680 242196 181686 242208
rect 192386 242196 192392 242208
rect 181680 242168 192392 242196
rect 181680 242156 181686 242168
rect 192386 242156 192392 242168
rect 192444 242156 192450 242208
rect 197262 242156 197268 242208
rect 197320 242196 197326 242208
rect 238389 242199 238447 242205
rect 238389 242196 238401 242199
rect 197320 242168 238401 242196
rect 197320 242156 197326 242168
rect 238389 242165 238401 242168
rect 238435 242165 238447 242199
rect 238389 242159 238447 242165
rect 238481 242199 238539 242205
rect 238481 242165 238493 242199
rect 238527 242196 238539 242199
rect 249150 242196 249156 242208
rect 238527 242168 249156 242196
rect 238527 242165 238539 242168
rect 238481 242159 238539 242165
rect 249150 242156 249156 242168
rect 249208 242156 249214 242208
rect 252462 242156 252468 242208
rect 252520 242196 252526 242208
rect 279142 242196 279148 242208
rect 252520 242168 279148 242196
rect 252520 242156 252526 242168
rect 279142 242156 279148 242168
rect 279200 242156 279206 242208
rect 280062 242156 280068 242208
rect 280120 242196 280126 242208
rect 293770 242196 293776 242208
rect 280120 242168 293776 242196
rect 280120 242156 280126 242168
rect 293770 242156 293776 242168
rect 293828 242156 293834 242208
rect 318242 242156 318248 242208
rect 318300 242196 318306 242208
rect 327258 242196 327264 242208
rect 318300 242168 327264 242196
rect 318300 242156 318306 242168
rect 327258 242156 327264 242168
rect 327316 242156 327322 242208
rect 332318 242156 332324 242208
rect 332376 242196 332382 242208
rect 345661 242199 345719 242205
rect 345661 242196 345673 242199
rect 332376 242168 345673 242196
rect 332376 242156 332382 242168
rect 345661 242165 345673 242168
rect 345707 242165 345719 242199
rect 345661 242159 345719 242165
rect 348786 242156 348792 242208
rect 348844 242196 348850 242208
rect 379517 242199 379575 242205
rect 379517 242196 379529 242199
rect 348844 242168 379529 242196
rect 348844 242156 348850 242168
rect 379517 242165 379529 242168
rect 379563 242165 379575 242199
rect 379517 242159 379575 242165
rect 379609 242199 379667 242205
rect 379609 242165 379621 242199
rect 379655 242196 379667 242199
rect 388622 242196 388628 242208
rect 379655 242168 388628 242196
rect 379655 242165 379667 242168
rect 379609 242159 379667 242165
rect 388622 242156 388628 242168
rect 388680 242156 388686 242208
rect 392210 242156 392216 242208
rect 392268 242196 392274 242208
rect 395525 242199 395583 242205
rect 395525 242196 395537 242199
rect 392268 242168 395537 242196
rect 392268 242156 392274 242168
rect 395525 242165 395537 242168
rect 395571 242165 395583 242199
rect 395525 242159 395583 242165
rect 406838 242156 406844 242208
rect 406896 242196 406902 242208
rect 499574 242196 499580 242208
rect 406896 242168 499580 242196
rect 406896 242156 406902 242168
rect 499574 242156 499580 242168
rect 499632 242156 499638 242208
rect 98638 242088 98644 242140
rect 98696 242128 98702 242140
rect 103422 242128 103428 242140
rect 98696 242100 103428 242128
rect 98696 242088 98702 242100
rect 103422 242088 103428 242100
rect 103480 242088 103486 242140
rect 104802 242088 104808 242140
rect 104860 242128 104866 242140
rect 203334 242128 203340 242140
rect 104860 242100 203340 242128
rect 104860 242088 104866 242100
rect 203334 242088 203340 242100
rect 203392 242088 203398 242140
rect 215202 242088 215208 242140
rect 215260 242128 215266 242140
rect 220081 242131 220139 242137
rect 220081 242128 220093 242131
rect 215260 242100 220093 242128
rect 215260 242088 215266 242100
rect 220081 242097 220093 242100
rect 220127 242097 220139 242131
rect 220081 242091 220139 242097
rect 226242 242088 226248 242140
rect 226300 242128 226306 242140
rect 265710 242128 265716 242140
rect 226300 242100 265716 242128
rect 226300 242088 226306 242100
rect 265710 242088 265716 242100
rect 265768 242088 265774 242140
rect 267642 242088 267648 242140
rect 267700 242128 267706 242140
rect 287054 242128 287060 242140
rect 267700 242100 287060 242128
rect 267700 242088 267706 242100
rect 287054 242088 287060 242100
rect 287112 242088 287118 242140
rect 343910 242088 343916 242140
rect 343968 242128 343974 242140
rect 343968 242100 374224 242128
rect 343968 242088 343974 242100
rect 77938 242020 77944 242072
rect 77996 242060 78002 242072
rect 175826 242060 175832 242072
rect 77996 242032 175832 242060
rect 77996 242020 78002 242032
rect 175826 242020 175832 242032
rect 175884 242020 175890 242072
rect 202138 242020 202144 242072
rect 202196 242060 202202 242072
rect 243722 242060 243728 242072
rect 202196 242032 243728 242060
rect 202196 242020 202202 242032
rect 243722 242020 243728 242032
rect 243780 242020 243786 242072
rect 244182 242020 244188 242072
rect 244240 242060 244246 242072
rect 268381 242063 268439 242069
rect 268381 242060 268393 242063
rect 244240 242032 268393 242060
rect 244240 242020 244246 242032
rect 268381 242029 268393 242032
rect 268427 242029 268439 242063
rect 268381 242023 268439 242029
rect 268470 242020 268476 242072
rect 268528 242060 268534 242072
rect 275462 242060 275468 242072
rect 268528 242032 275468 242060
rect 268528 242020 268534 242032
rect 275462 242020 275468 242032
rect 275520 242020 275526 242072
rect 275922 242020 275928 242072
rect 275980 242060 275986 242072
rect 291378 242060 291384 242072
rect 275980 242032 291384 242060
rect 275980 242020 275986 242032
rect 291378 242020 291384 242032
rect 291436 242020 291442 242072
rect 342714 242020 342720 242072
rect 342772 242060 342778 242072
rect 374086 242060 374092 242072
rect 342772 242032 374092 242060
rect 342772 242020 342778 242032
rect 374086 242020 374092 242032
rect 374144 242020 374150 242072
rect 374196 242060 374224 242100
rect 374270 242088 374276 242140
rect 374328 242128 374334 242140
rect 384298 242128 384304 242140
rect 374328 242100 384304 242128
rect 374328 242088 374334 242100
rect 384298 242088 384304 242100
rect 384356 242088 384362 242140
rect 384850 242088 384856 242140
rect 384908 242128 384914 242140
rect 393961 242131 394019 242137
rect 393961 242128 393973 242131
rect 384908 242100 393973 242128
rect 384908 242088 384914 242100
rect 393961 242097 393973 242100
rect 394007 242097 394019 242131
rect 393961 242091 394019 242097
rect 408678 242088 408684 242140
rect 408736 242128 408742 242140
rect 412821 242131 412879 242137
rect 412821 242128 412833 242131
rect 408736 242100 412833 242128
rect 408736 242088 408742 242100
rect 412821 242097 412833 242100
rect 412867 242097 412879 242131
rect 412821 242091 412879 242097
rect 412910 242088 412916 242140
rect 412968 242128 412974 242140
rect 413922 242128 413928 242140
rect 412968 242100 413928 242128
rect 412968 242088 412974 242100
rect 413922 242088 413928 242100
rect 413980 242088 413986 242140
rect 415394 242088 415400 242140
rect 415452 242128 415458 242140
rect 416498 242128 416504 242140
rect 415452 242100 416504 242128
rect 415452 242088 415458 242100
rect 416498 242088 416504 242100
rect 416556 242088 416562 242140
rect 417234 242088 417240 242140
rect 417292 242128 417298 242140
rect 418062 242128 418068 242140
rect 417292 242100 418068 242128
rect 417292 242088 417298 242100
rect 418062 242088 418068 242100
rect 418120 242088 418126 242140
rect 418249 242131 418307 242137
rect 418249 242097 418261 242131
rect 418295 242128 418307 242131
rect 419537 242131 419595 242137
rect 419537 242128 419549 242131
rect 418295 242100 419549 242128
rect 418295 242097 418307 242100
rect 418249 242091 418307 242097
rect 419537 242097 419549 242100
rect 419583 242097 419595 242131
rect 419537 242091 419595 242097
rect 419626 242088 419632 242140
rect 419684 242128 419690 242140
rect 421650 242128 421656 242140
rect 419684 242100 421656 242128
rect 419684 242088 419690 242100
rect 421650 242088 421656 242100
rect 421708 242088 421714 242140
rect 440418 242088 440424 242140
rect 440476 242128 440482 242140
rect 441522 242128 441528 242140
rect 440476 242100 441528 242128
rect 440476 242088 440482 242100
rect 441522 242088 441528 242100
rect 441580 242088 441586 242140
rect 441706 242088 441712 242140
rect 441764 242128 441770 242140
rect 442994 242128 443000 242140
rect 441764 242100 443000 242128
rect 441764 242088 441770 242100
rect 442994 242088 443000 242100
rect 443052 242088 443058 242140
rect 443089 242131 443147 242137
rect 443089 242097 443101 242131
rect 443135 242128 443147 242131
rect 445754 242128 445760 242140
rect 443135 242100 445760 242128
rect 443135 242097 443147 242100
rect 443089 242091 443147 242097
rect 445754 242088 445760 242100
rect 445812 242088 445818 242140
rect 447134 242088 447140 242140
rect 447192 242128 447198 242140
rect 449989 242131 450047 242137
rect 447192 242100 449940 242128
rect 447192 242088 447198 242100
rect 376018 242060 376024 242072
rect 374196 242032 376024 242060
rect 376018 242020 376024 242032
rect 376076 242020 376082 242072
rect 379330 242020 379336 242072
rect 379388 242060 379394 242072
rect 442629 242063 442687 242069
rect 442629 242060 442641 242063
rect 379388 242032 442641 242060
rect 379388 242020 379394 242032
rect 442629 242029 442641 242032
rect 442675 242029 442687 242063
rect 442629 242023 442687 242029
rect 442718 242020 442724 242072
rect 442776 242060 442782 242072
rect 442902 242060 442908 242072
rect 442776 242032 442908 242060
rect 442776 242020 442782 242032
rect 442902 242020 442908 242032
rect 442960 242020 442966 242072
rect 444742 242020 444748 242072
rect 444800 242060 444806 242072
rect 445570 242060 445576 242072
rect 444800 242032 445576 242060
rect 444800 242020 444806 242032
rect 445570 242020 445576 242032
rect 445628 242020 445634 242072
rect 445938 242020 445944 242072
rect 445996 242060 446002 242072
rect 447042 242060 447048 242072
rect 445996 242032 447048 242060
rect 445996 242020 446002 242032
rect 447042 242020 447048 242032
rect 447100 242020 447106 242072
rect 447778 242020 447784 242072
rect 447836 242060 447842 242072
rect 448422 242060 448428 242072
rect 447836 242032 448428 242060
rect 447836 242020 447842 242032
rect 448422 242020 448428 242032
rect 448480 242020 448486 242072
rect 448974 242020 448980 242072
rect 449032 242060 449038 242072
rect 449802 242060 449808 242072
rect 449032 242032 449808 242060
rect 449032 242020 449038 242032
rect 449802 242020 449808 242032
rect 449860 242020 449866 242072
rect 449912 242060 449940 242100
rect 449989 242097 450001 242131
rect 450035 242128 450047 242131
rect 529198 242128 529204 242140
rect 450035 242100 529204 242128
rect 450035 242097 450047 242100
rect 449989 242091 450047 242097
rect 529198 242088 529204 242100
rect 529256 242088 529262 242140
rect 530578 242060 530584 242072
rect 449912 242032 530584 242060
rect 530578 242020 530584 242032
rect 530636 242020 530642 242072
rect 75178 241952 75184 242004
rect 75236 241992 75242 242004
rect 173434 241992 173440 242004
rect 75236 241964 173440 241992
rect 75236 241952 75242 241964
rect 173434 241952 173440 241964
rect 173492 241952 173498 242004
rect 177298 241952 177304 242004
rect 177356 241992 177362 242004
rect 185026 241992 185032 242004
rect 177356 241964 185032 241992
rect 177356 241952 177362 241964
rect 185026 241952 185032 241964
rect 185084 241952 185090 242004
rect 200758 241952 200764 242004
rect 200816 241992 200822 242004
rect 228450 241992 228456 242004
rect 200816 241964 228456 241992
rect 200816 241952 200822 241964
rect 228450 241952 228456 241964
rect 228508 241952 228514 242004
rect 231762 241952 231768 242004
rect 231820 241992 231826 242004
rect 268746 241992 268752 242004
rect 231820 241964 268752 241992
rect 231820 241952 231826 241964
rect 268746 241952 268752 241964
rect 268804 241952 268810 242004
rect 269022 241952 269028 242004
rect 269080 241992 269086 242004
rect 287698 241992 287704 242004
rect 269080 241964 287704 241992
rect 269080 241952 269086 241964
rect 287698 241952 287704 241964
rect 287756 241952 287762 242004
rect 345937 241995 345995 242001
rect 345937 241961 345949 241995
rect 345983 241992 345995 241995
rect 372798 241992 372804 242004
rect 345983 241964 372804 241992
rect 345983 241961 345995 241964
rect 345937 241955 345995 241961
rect 372798 241952 372804 241964
rect 372856 241952 372862 242004
rect 375098 241952 375104 242004
rect 375156 241992 375162 242004
rect 394050 241992 394056 242004
rect 375156 241964 394056 241992
rect 375156 241952 375162 241964
rect 394050 241952 394056 241964
rect 394108 241952 394114 242004
rect 395798 241952 395804 242004
rect 395856 241992 395862 242004
rect 477586 241992 477592 242004
rect 395856 241964 477592 241992
rect 395856 241952 395862 241964
rect 477586 241952 477592 241964
rect 477644 241952 477650 242004
rect 111702 241884 111708 241936
rect 111760 241924 111766 241936
rect 207014 241924 207020 241936
rect 111760 241896 207020 241924
rect 111760 241884 111766 241896
rect 207014 241884 207020 241896
rect 207072 241884 207078 241936
rect 232498 241884 232504 241936
rect 232556 241924 232562 241936
rect 261481 241927 261539 241933
rect 261481 241924 261493 241927
rect 232556 241896 261493 241924
rect 232556 241884 232562 241896
rect 261481 241893 261493 241896
rect 261527 241893 261539 241927
rect 261481 241887 261539 241893
rect 261570 241884 261576 241936
rect 261628 241924 261634 241936
rect 263870 241924 263876 241936
rect 261628 241896 263876 241924
rect 261628 241884 261634 241896
rect 263870 241884 263876 241896
rect 263928 241884 263934 241936
rect 271782 241884 271788 241936
rect 271840 241924 271846 241936
rect 289538 241924 289544 241936
rect 271840 241896 289544 241924
rect 271840 241884 271846 241896
rect 289538 241884 289544 241896
rect 289596 241884 289602 241936
rect 335354 241884 335360 241936
rect 335412 241924 335418 241936
rect 344005 241927 344063 241933
rect 344005 241924 344017 241927
rect 335412 241896 344017 241924
rect 335412 241884 335418 241896
rect 344005 241893 344017 241896
rect 344051 241893 344063 241927
rect 344005 241887 344063 241893
rect 344097 241927 344155 241933
rect 344097 241893 344109 241927
rect 344143 241924 344155 241927
rect 350810 241924 350816 241936
rect 344143 241896 350816 241924
rect 344143 241893 344155 241896
rect 344097 241887 344155 241893
rect 350810 241884 350816 241896
rect 350868 241884 350874 241936
rect 350905 241927 350963 241933
rect 350905 241893 350917 241927
rect 350951 241924 350963 241927
rect 355137 241927 355195 241933
rect 355137 241924 355149 241927
rect 350951 241896 355149 241924
rect 350951 241893 350963 241896
rect 350905 241887 350963 241893
rect 355137 241893 355149 241896
rect 355183 241893 355195 241927
rect 355137 241887 355195 241893
rect 355229 241927 355287 241933
rect 355229 241893 355241 241927
rect 355275 241924 355287 241927
rect 380158 241924 380164 241936
rect 355275 241896 380164 241924
rect 355275 241893 355287 241896
rect 355229 241887 355287 241893
rect 380158 241884 380164 241896
rect 380216 241884 380222 241936
rect 391382 241924 391388 241936
rect 384316 241896 391388 241924
rect 84838 241816 84844 241868
rect 84896 241856 84902 241868
rect 179506 241856 179512 241868
rect 84896 241828 179512 241856
rect 84896 241816 84902 241828
rect 179506 241816 179512 241828
rect 179564 241816 179570 241868
rect 188430 241816 188436 241868
rect 188488 241856 188494 241868
rect 204806 241856 204812 241868
rect 188488 241828 204812 241856
rect 188488 241816 188494 241828
rect 204806 241816 204812 241828
rect 204864 241816 204870 241868
rect 204898 241816 204904 241868
rect 204956 241856 204962 241868
rect 241238 241856 241244 241868
rect 204956 241828 241244 241856
rect 204956 241816 204962 241828
rect 241238 241816 241244 241828
rect 241296 241816 241302 241868
rect 241422 241816 241428 241868
rect 241480 241856 241486 241868
rect 273622 241856 273628 241868
rect 241480 241828 273628 241856
rect 241480 241816 241486 241828
rect 273622 241816 273628 241828
rect 273680 241816 273686 241868
rect 274361 241859 274419 241865
rect 274361 241825 274373 241859
rect 274407 241856 274419 241859
rect 278498 241856 278504 241868
rect 274407 241828 278504 241856
rect 274407 241825 274419 241828
rect 274361 241819 274419 241825
rect 278498 241816 278504 241828
rect 278556 241816 278562 241868
rect 339586 241816 339592 241868
rect 339644 241856 339650 241868
rect 368474 241856 368480 241868
rect 339644 241828 368480 241856
rect 339644 241816 339650 241828
rect 368474 241816 368480 241828
rect 368532 241816 368538 241868
rect 371418 241816 371424 241868
rect 371476 241856 371482 241868
rect 384316 241856 384344 241896
rect 391382 241884 391388 241896
rect 391440 241884 391446 241936
rect 393406 241884 393412 241936
rect 393464 241924 393470 241936
rect 473354 241924 473360 241936
rect 393464 241896 473360 241924
rect 393464 241884 393470 241896
rect 473354 241884 473360 241896
rect 473412 241884 473418 241936
rect 371476 241828 384344 241856
rect 371476 241816 371482 241828
rect 388530 241816 388536 241868
rect 388588 241856 388594 241868
rect 395525 241859 395583 241865
rect 388588 241828 393912 241856
rect 388588 241816 388594 241828
rect 103517 241791 103575 241797
rect 103517 241757 103529 241791
rect 103563 241788 103575 241791
rect 113085 241791 113143 241797
rect 113085 241788 113097 241791
rect 103563 241760 113097 241788
rect 103563 241757 103575 241760
rect 103517 241751 103575 241757
rect 113085 241757 113097 241760
rect 113131 241757 113143 241791
rect 113085 241751 113143 241757
rect 115842 241748 115848 241800
rect 115900 241788 115906 241800
rect 208854 241788 208860 241800
rect 115900 241760 208860 241788
rect 115900 241748 115906 241760
rect 208854 241748 208860 241760
rect 208912 241748 208918 241800
rect 238665 241791 238723 241797
rect 238665 241757 238677 241791
rect 238711 241788 238723 241791
rect 272426 241788 272432 241800
rect 238711 241760 272432 241788
rect 238711 241757 238723 241760
rect 238665 241751 238723 241757
rect 272426 241748 272432 241760
rect 272484 241748 272490 241800
rect 273162 241748 273168 241800
rect 273220 241788 273226 241800
rect 290090 241788 290096 241800
rect 273220 241760 290096 241788
rect 273220 241748 273226 241760
rect 290090 241748 290096 241760
rect 290148 241748 290154 241800
rect 291102 241748 291108 241800
rect 291160 241788 291166 241800
rect 299290 241788 299296 241800
rect 291160 241760 299296 241788
rect 291160 241748 291166 241760
rect 299290 241748 299296 241760
rect 299348 241748 299354 241800
rect 334158 241748 334164 241800
rect 334216 241788 334222 241800
rect 355321 241791 355379 241797
rect 334216 241760 353984 241788
rect 334216 241748 334222 241760
rect 113177 241723 113235 241729
rect 113177 241689 113189 241723
rect 113223 241720 113235 241723
rect 122653 241723 122711 241729
rect 122653 241720 122665 241723
rect 113223 241692 122665 241720
rect 113223 241689 113235 241692
rect 113177 241683 113235 241689
rect 122653 241689 122665 241692
rect 122699 241689 122711 241723
rect 122653 241683 122711 241689
rect 122742 241680 122748 241732
rect 122800 241720 122806 241732
rect 212534 241720 212540 241732
rect 122800 241692 212540 241720
rect 122800 241680 122806 241692
rect 212534 241680 212540 241692
rect 212592 241680 212598 241732
rect 226978 241680 226984 241732
rect 227036 241720 227042 241732
rect 255866 241720 255872 241732
rect 227036 241692 255872 241720
rect 227036 241680 227042 241692
rect 255866 241680 255872 241692
rect 255924 241680 255930 241732
rect 257338 241680 257344 241732
rect 257396 241720 257402 241732
rect 261386 241720 261392 241732
rect 257396 241692 261392 241720
rect 257396 241680 257402 241692
rect 261386 241680 261392 241692
rect 261444 241680 261450 241732
rect 262858 241680 262864 241732
rect 262916 241720 262922 241732
rect 265066 241720 265072 241732
rect 262916 241692 265072 241720
rect 262916 241680 262922 241692
rect 265066 241680 265072 241692
rect 265124 241680 265130 241732
rect 270402 241680 270408 241732
rect 270460 241720 270466 241732
rect 287974 241720 287980 241732
rect 270460 241692 287980 241720
rect 270460 241680 270466 241692
rect 287974 241680 287980 241692
rect 288032 241680 288038 241732
rect 318886 241680 318892 241732
rect 318944 241720 318950 241732
rect 323578 241720 323584 241732
rect 318944 241692 323584 241720
rect 318944 241680 318950 241692
rect 323578 241680 323584 241692
rect 323636 241680 323642 241732
rect 330754 241680 330760 241732
rect 330812 241720 330818 241732
rect 344097 241723 344155 241729
rect 344097 241720 344109 241723
rect 330812 241692 344109 241720
rect 330812 241680 330818 241692
rect 344097 241689 344109 241692
rect 344143 241689 344155 241723
rect 344097 241683 344155 241689
rect 344189 241723 344247 241729
rect 344189 241689 344201 241723
rect 344235 241720 344247 241723
rect 345658 241720 345664 241732
rect 344235 241692 345664 241720
rect 344235 241689 344247 241692
rect 344189 241683 344247 241689
rect 345658 241680 345664 241692
rect 345716 241680 345722 241732
rect 349430 241680 349436 241732
rect 349488 241720 349494 241732
rect 350442 241720 350448 241732
rect 349488 241692 350448 241720
rect 349488 241680 349494 241692
rect 350442 241680 350448 241692
rect 350500 241680 350506 241732
rect 350537 241723 350595 241729
rect 350537 241689 350549 241723
rect 350583 241720 350595 241723
rect 353297 241723 353355 241729
rect 353297 241720 353309 241723
rect 350583 241692 353309 241720
rect 350583 241689 350595 241692
rect 350537 241683 350595 241689
rect 353297 241689 353309 241692
rect 353343 241689 353355 241723
rect 353956 241720 353984 241760
rect 355321 241757 355333 241791
rect 355367 241788 355379 241791
rect 365806 241788 365812 241800
rect 355367 241760 365812 241788
rect 355367 241757 355379 241760
rect 355321 241751 355379 241757
rect 365806 241748 365812 241760
rect 365864 241748 365870 241800
rect 367370 241748 367376 241800
rect 367428 241788 367434 241800
rect 368382 241788 368388 241800
rect 367428 241760 368388 241788
rect 367428 241748 367434 241760
rect 368382 241748 368388 241760
rect 368440 241748 368446 241800
rect 369118 241748 369124 241800
rect 369176 241788 369182 241800
rect 379517 241791 379575 241797
rect 379517 241788 379529 241791
rect 369176 241760 379529 241788
rect 369176 241748 369182 241760
rect 379517 241757 379529 241760
rect 379563 241757 379575 241791
rect 384482 241788 384488 241800
rect 379517 241751 379575 241757
rect 379624 241760 384488 241788
rect 357434 241720 357440 241732
rect 353956 241692 357440 241720
rect 353297 241683 353355 241689
rect 357434 241680 357440 241692
rect 357492 241680 357498 241732
rect 379624 241720 379652 241760
rect 384482 241748 384488 241760
rect 384540 241748 384546 241800
rect 391290 241720 391296 241732
rect 360304 241692 379652 241720
rect 381004 241692 391296 241720
rect 95878 241612 95884 241664
rect 95936 241652 95942 241664
rect 174078 241652 174084 241664
rect 95936 241624 174084 241652
rect 95936 241612 95942 241624
rect 174078 241612 174084 241624
rect 174136 241612 174142 241664
rect 174538 241612 174544 241664
rect 174596 241652 174602 241664
rect 177666 241652 177672 241664
rect 174596 241624 177672 241652
rect 174596 241612 174602 241624
rect 177666 241612 177672 241624
rect 177724 241612 177730 241664
rect 191098 241612 191104 241664
rect 191156 241652 191162 241664
rect 214374 241652 214380 241664
rect 191156 241624 214380 241652
rect 191156 241612 191162 241624
rect 214374 241612 214380 241624
rect 214432 241612 214438 241664
rect 243538 241612 243544 241664
rect 243596 241652 243602 241664
rect 271230 241652 271236 241664
rect 243596 241624 271236 241652
rect 243596 241612 243602 241624
rect 271230 241612 271236 241624
rect 271288 241612 271294 241664
rect 271325 241655 271383 241661
rect 271325 241621 271337 241655
rect 271371 241652 271383 241655
rect 271371 241624 274496 241652
rect 271371 241621 271383 241624
rect 271325 241615 271383 241621
rect 106918 241544 106924 241596
rect 106976 241584 106982 241596
rect 183186 241584 183192 241596
rect 106976 241556 183192 241584
rect 106976 241544 106982 241556
rect 183186 241544 183192 241556
rect 183244 241544 183250 241596
rect 238389 241587 238447 241593
rect 238389 241553 238401 241587
rect 238435 241584 238447 241587
rect 250990 241584 250996 241596
rect 238435 241556 250996 241584
rect 238435 241553 238447 241556
rect 238389 241547 238447 241553
rect 250990 241544 250996 241556
rect 251048 241544 251054 241596
rect 251082 241544 251088 241596
rect 251140 241584 251146 241596
rect 274361 241587 274419 241593
rect 274361 241584 274373 241587
rect 251140 241556 274373 241584
rect 251140 241544 251146 241556
rect 274361 241553 274373 241556
rect 274407 241553 274419 241587
rect 274468 241584 274496 241624
rect 274542 241612 274548 241664
rect 274600 241652 274606 241664
rect 290734 241652 290740 241664
rect 274600 241624 290740 241652
rect 274600 241612 274606 241624
rect 290734 241612 290740 241624
rect 290792 241612 290798 241664
rect 298738 241612 298744 241664
rect 298796 241652 298802 241664
rect 301774 241652 301780 241664
rect 298796 241624 301780 241652
rect 298796 241612 298802 241624
rect 301774 241612 301780 241624
rect 301832 241612 301838 241664
rect 302878 241612 302884 241664
rect 302936 241652 302942 241664
rect 304810 241652 304816 241664
rect 302936 241624 304816 241652
rect 302936 241612 302942 241624
rect 304810 241612 304816 241624
rect 304868 241612 304874 241664
rect 317046 241612 317052 241664
rect 317104 241652 317110 241664
rect 322198 241652 322204 241664
rect 317104 241624 322204 241652
rect 317104 241612 317110 241624
rect 322198 241612 322204 241624
rect 322256 241612 322262 241664
rect 337194 241612 337200 241664
rect 337252 241652 337258 241664
rect 337252 241624 338988 241652
rect 337252 241612 337258 241624
rect 276106 241584 276112 241596
rect 274468 241556 276112 241584
rect 274361 241547 274419 241553
rect 276106 241544 276112 241556
rect 276164 241544 276170 241596
rect 290458 241544 290464 241596
rect 290516 241584 290522 241596
rect 296254 241584 296260 241596
rect 290516 241556 296260 241584
rect 290516 241544 290522 241556
rect 296254 241544 296260 241556
rect 296312 241544 296318 241596
rect 297450 241544 297456 241596
rect 297508 241584 297514 241596
rect 301130 241584 301136 241596
rect 297508 241556 301136 241584
rect 297508 241544 297514 241556
rect 301130 241544 301136 241556
rect 301188 241544 301194 241596
rect 301498 241544 301504 241596
rect 301556 241584 301562 241596
rect 303614 241584 303620 241596
rect 301556 241556 303620 241584
rect 301556 241544 301562 241556
rect 303614 241544 303620 241556
rect 303672 241544 303678 241596
rect 304258 241544 304264 241596
rect 304316 241584 304322 241596
rect 305362 241584 305368 241596
rect 304316 241556 305368 241584
rect 304316 241544 304322 241556
rect 305362 241544 305368 241556
rect 305420 241544 305426 241596
rect 310330 241544 310336 241596
rect 310388 241584 310394 241596
rect 311894 241584 311900 241596
rect 310388 241556 311900 241584
rect 310388 241544 310394 241556
rect 311894 241544 311900 241556
rect 311952 241544 311958 241596
rect 312170 241544 312176 241596
rect 312228 241584 312234 241596
rect 314838 241584 314844 241596
rect 312228 241556 314844 241584
rect 312228 241544 312234 241556
rect 314838 241544 314844 241556
rect 314896 241544 314902 241596
rect 316402 241544 316408 241596
rect 316460 241584 316466 241596
rect 320818 241584 320824 241596
rect 316460 241556 320824 241584
rect 316460 241544 316466 241556
rect 320818 241544 320824 241556
rect 320876 241544 320882 241596
rect 329190 241544 329196 241596
rect 329248 241584 329254 241596
rect 333238 241584 333244 241596
rect 329248 241556 333244 241584
rect 329248 241544 329254 241556
rect 333238 241544 333244 241556
rect 333296 241544 333302 241596
rect 336550 241544 336556 241596
rect 336608 241584 336614 241596
rect 338850 241584 338856 241596
rect 336608 241556 338856 241584
rect 336608 241544 336614 241556
rect 338850 241544 338856 241556
rect 338908 241544 338914 241596
rect 338960 241584 338988 241624
rect 339034 241612 339040 241664
rect 339092 241652 339098 241664
rect 358078 241652 358084 241664
rect 339092 241624 358084 241652
rect 339092 241612 339098 241624
rect 358078 241612 358084 241624
rect 358136 241612 358142 241664
rect 356698 241584 356704 241596
rect 338960 241556 356704 241584
rect 356698 241544 356704 241556
rect 356756 241544 356762 241596
rect 357066 241544 357072 241596
rect 357124 241584 357130 241596
rect 360304 241584 360332 241692
rect 360378 241612 360384 241664
rect 360436 241652 360442 241664
rect 369118 241652 369124 241664
rect 360436 241624 369124 241652
rect 360436 241612 360442 241624
rect 369118 241612 369124 241624
rect 369176 241612 369182 241664
rect 377490 241612 377496 241664
rect 377548 241652 377554 241664
rect 380250 241652 380256 241664
rect 377548 241624 380256 241652
rect 377548 241612 377554 241624
rect 380250 241612 380256 241624
rect 380308 241612 380314 241664
rect 357124 241556 360332 241584
rect 367189 241587 367247 241593
rect 357124 241544 357130 241556
rect 367189 241553 367201 241587
rect 367235 241584 367247 241587
rect 375558 241584 375564 241596
rect 367235 241556 375564 241584
rect 367235 241553 367247 241556
rect 367189 241547 367247 241553
rect 375558 241544 375564 241556
rect 375616 241544 375622 241596
rect 381004 241584 381032 241692
rect 391290 241680 391296 241692
rect 391348 241680 391354 241732
rect 393884 241720 393912 241828
rect 395525 241825 395537 241859
rect 395571 241856 395583 241859
rect 470594 241856 470600 241868
rect 395571 241828 470600 241856
rect 395571 241825 395583 241828
rect 395525 241819 395583 241825
rect 470594 241816 470600 241828
rect 470652 241816 470658 241868
rect 394237 241791 394295 241797
rect 394237 241757 394249 241791
rect 394283 241788 394295 241791
rect 466454 241788 466460 241800
rect 394283 241760 466460 241788
rect 394283 241757 394295 241760
rect 394237 241751 394295 241757
rect 466454 241748 466460 241760
rect 466512 241748 466518 241800
rect 463694 241720 463700 241732
rect 393884 241692 463700 241720
rect 463694 241680 463700 241692
rect 463752 241680 463758 241732
rect 383010 241612 383016 241664
rect 383068 241652 383074 241664
rect 383068 241624 388668 241652
rect 383068 241612 383074 241624
rect 379900 241556 381032 241584
rect 113174 241476 113180 241528
rect 113232 241516 113238 241528
rect 122650 241516 122656 241528
rect 113232 241488 122656 241516
rect 113232 241476 113238 241488
rect 122650 241476 122656 241488
rect 122708 241476 122714 241528
rect 142157 241519 142215 241525
rect 142157 241485 142169 241519
rect 142203 241516 142215 241519
rect 152553 241519 152611 241525
rect 152553 241516 152565 241519
rect 142203 241488 152565 241516
rect 142203 241485 142215 241488
rect 142157 241479 142215 241485
rect 152553 241485 152565 241488
rect 152599 241485 152611 241519
rect 152553 241479 152611 241485
rect 160830 241476 160836 241528
rect 160888 241516 160894 241528
rect 208210 241516 208216 241528
rect 160888 241488 208216 241516
rect 160888 241476 160894 241488
rect 208210 241476 208216 241488
rect 208268 241476 208274 241528
rect 238662 241516 238668 241528
rect 238623 241488 238668 241516
rect 238662 241476 238668 241488
rect 238720 241476 238726 241528
rect 250438 241476 250444 241528
rect 250496 241516 250502 241528
rect 257706 241516 257712 241528
rect 250496 241488 257712 241516
rect 250496 241476 250502 241488
rect 257706 241476 257712 241488
rect 257764 241476 257770 241528
rect 261478 241476 261484 241528
rect 261536 241516 261542 241528
rect 263226 241516 263232 241528
rect 261536 241488 263232 241516
rect 261536 241476 261542 241488
rect 263226 241476 263232 241488
rect 263284 241476 263290 241528
rect 263502 241476 263508 241528
rect 263560 241516 263566 241528
rect 268289 241519 268347 241525
rect 268289 241516 268301 241519
rect 263560 241488 268301 241516
rect 263560 241476 263566 241488
rect 268289 241485 268301 241488
rect 268335 241485 268347 241519
rect 268289 241479 268347 241485
rect 268381 241519 268439 241525
rect 268381 241485 268393 241519
rect 268427 241516 268439 241519
rect 274818 241516 274824 241528
rect 268427 241488 274824 241516
rect 268427 241485 268439 241488
rect 268381 241479 268439 241485
rect 274818 241476 274824 241488
rect 274876 241476 274882 241528
rect 280798 241476 280804 241528
rect 280856 241516 280862 241528
rect 283374 241516 283380 241528
rect 280856 241488 283380 241516
rect 280856 241476 280862 241488
rect 283374 241476 283380 241488
rect 283432 241476 283438 241528
rect 291838 241476 291844 241528
rect 291896 241516 291902 241528
rect 293218 241516 293224 241528
rect 291896 241488 293224 241516
rect 291896 241476 291902 241488
rect 293218 241476 293224 241488
rect 293276 241476 293282 241528
rect 297358 241476 297364 241528
rect 297416 241516 297422 241528
rect 298646 241516 298652 241528
rect 297416 241488 298652 241516
rect 297416 241476 297422 241488
rect 298646 241476 298652 241488
rect 298704 241476 298710 241528
rect 298830 241476 298836 241528
rect 298888 241516 298894 241528
rect 300486 241516 300492 241528
rect 298888 241488 300492 241516
rect 298888 241476 298894 241488
rect 300486 241476 300492 241488
rect 300544 241476 300550 241528
rect 301590 241476 301596 241528
rect 301648 241516 301654 241528
rect 302970 241516 302976 241528
rect 301648 241488 302976 241516
rect 301648 241476 301654 241488
rect 302970 241476 302976 241488
rect 303028 241476 303034 241528
rect 304902 241476 304908 241528
rect 304960 241516 304966 241528
rect 306006 241516 306012 241528
rect 304960 241488 306012 241516
rect 304960 241476 304966 241488
rect 306006 241476 306012 241488
rect 306064 241476 306070 241528
rect 307202 241516 307208 241528
rect 306300 241488 307208 241516
rect 306300 241460 306328 241488
rect 307202 241476 307208 241488
rect 307260 241476 307266 241528
rect 309686 241476 309692 241528
rect 309744 241516 309750 241528
rect 310422 241516 310428 241528
rect 309744 241488 310428 241516
rect 309744 241476 309750 241488
rect 310422 241476 310428 241488
rect 310480 241476 310486 241528
rect 310882 241476 310888 241528
rect 310940 241516 310946 241528
rect 312538 241516 312544 241528
rect 310940 241488 312544 241516
rect 310940 241476 310946 241488
rect 312538 241476 312544 241488
rect 312596 241476 312602 241528
rect 320634 241476 320640 241528
rect 320692 241516 320698 241528
rect 321462 241516 321468 241528
rect 320692 241488 321468 241516
rect 320692 241476 320698 241488
rect 321462 241476 321468 241488
rect 321520 241476 321526 241528
rect 321922 241476 321928 241528
rect 321980 241516 321986 241528
rect 322842 241516 322848 241528
rect 321980 241488 322848 241516
rect 321980 241476 321986 241488
rect 322842 241476 322848 241488
rect 322900 241476 322906 241528
rect 323118 241476 323124 241528
rect 323176 241516 323182 241528
rect 324130 241516 324136 241528
rect 323176 241488 324136 241516
rect 323176 241476 323182 241488
rect 324130 241476 324136 241488
rect 324188 241476 324194 241528
rect 324314 241476 324320 241528
rect 324372 241516 324378 241528
rect 325602 241516 325608 241528
rect 324372 241488 325608 241516
rect 324372 241476 324378 241488
rect 325602 241476 325608 241488
rect 325660 241476 325666 241528
rect 326154 241476 326160 241528
rect 326212 241516 326218 241528
rect 326982 241516 326988 241528
rect 326212 241488 326988 241516
rect 326212 241476 326218 241488
rect 326982 241476 326988 241488
rect 327040 241476 327046 241528
rect 327442 241476 327448 241528
rect 327500 241516 327506 241528
rect 328362 241516 328368 241528
rect 327500 241488 328368 241516
rect 327500 241476 327506 241488
rect 328362 241476 328368 241488
rect 328420 241476 328426 241528
rect 332870 241476 332876 241528
rect 332928 241516 332934 241528
rect 333882 241516 333888 241528
rect 332928 241488 333888 241516
rect 332928 241476 332934 241488
rect 333882 241476 333888 241488
rect 333940 241476 333946 241528
rect 338390 241476 338396 241528
rect 338448 241516 338454 241528
rect 339402 241516 339408 241528
rect 338448 241488 339408 241516
rect 338448 241476 338454 241488
rect 339402 241476 339408 241488
rect 339460 241476 339466 241528
rect 340874 241476 340880 241528
rect 340932 241516 340938 241528
rect 340932 241488 348096 241516
rect 340932 241476 340938 241488
rect 198274 241448 198280 241460
rect 198235 241420 198280 241448
rect 198274 241408 198280 241420
rect 198332 241408 198338 241460
rect 303798 241448 303804 241460
rect 303759 241420 303804 241448
rect 303798 241408 303804 241420
rect 303856 241408 303862 241460
rect 306282 241408 306288 241460
rect 306340 241408 306346 241460
rect 348068 241448 348096 241488
rect 348142 241476 348148 241528
rect 348200 241516 348206 241528
rect 349062 241516 349068 241528
rect 348200 241488 349068 241516
rect 348200 241476 348206 241488
rect 349062 241476 349068 241488
rect 349120 241476 349126 241528
rect 350537 241519 350595 241525
rect 350537 241516 350549 241519
rect 349172 241488 350549 241516
rect 349172 241448 349200 241488
rect 350537 241485 350549 241488
rect 350583 241485 350595 241519
rect 350537 241479 350595 241485
rect 352466 241476 352472 241528
rect 352524 241516 352530 241528
rect 353202 241516 353208 241528
rect 352524 241488 353208 241516
rect 352524 241476 352530 241488
rect 353202 241476 353208 241488
rect 353260 241476 353266 241528
rect 353297 241519 353355 241525
rect 353297 241485 353309 241519
rect 353343 241516 353355 241519
rect 354766 241516 354772 241528
rect 353343 241488 354772 241516
rect 353343 241485 353355 241488
rect 353297 241479 353355 241485
rect 354766 241476 354772 241488
rect 354824 241476 354830 241528
rect 354858 241476 354864 241528
rect 354916 241516 354922 241528
rect 355870 241516 355876 241528
rect 354916 241488 355876 241516
rect 354916 241476 354922 241488
rect 355870 241476 355876 241488
rect 355928 241476 355934 241528
rect 356146 241476 356152 241528
rect 356204 241516 356210 241528
rect 357342 241516 357348 241528
rect 356204 241488 357348 241516
rect 356204 241476 356210 241488
rect 357342 241476 357348 241488
rect 357400 241476 357406 241528
rect 357986 241476 357992 241528
rect 358044 241516 358050 241528
rect 358722 241516 358728 241528
rect 358044 241488 358728 241516
rect 358044 241476 358050 241488
rect 358722 241476 358728 241488
rect 358780 241476 358786 241528
rect 359182 241476 359188 241528
rect 359240 241516 359246 241528
rect 360102 241516 360108 241528
rect 359240 241488 360108 241516
rect 359240 241476 359246 241488
rect 360102 241476 360108 241488
rect 360160 241476 360166 241528
rect 361574 241476 361580 241528
rect 361632 241516 361638 241528
rect 362770 241516 362776 241528
rect 361632 241488 362776 241516
rect 361632 241476 361638 241488
rect 362770 241476 362776 241488
rect 362828 241476 362834 241528
rect 363414 241476 363420 241528
rect 363472 241516 363478 241528
rect 364242 241516 364248 241528
rect 363472 241488 364248 241516
rect 363472 241476 363478 241488
rect 364242 241476 364248 241488
rect 364300 241476 364306 241528
rect 365898 241476 365904 241528
rect 365956 241516 365962 241528
rect 367002 241516 367008 241528
rect 365956 241488 367008 241516
rect 365956 241476 365962 241488
rect 367002 241476 367008 241488
rect 367060 241476 367066 241528
rect 369949 241519 370007 241525
rect 369949 241485 369961 241519
rect 369995 241516 370007 241519
rect 369995 241488 370084 241516
rect 369995 241485 370007 241488
rect 369949 241479 370007 241485
rect 348068 241420 349200 241448
rect 355137 241451 355195 241457
rect 355137 241417 355149 241451
rect 355183 241448 355195 241451
rect 356330 241448 356336 241460
rect 355183 241420 356336 241448
rect 355183 241417 355195 241420
rect 355137 241411 355195 241417
rect 356330 241408 356336 241420
rect 356388 241408 356394 241460
rect 370056 241448 370084 241488
rect 371252 241488 372568 241516
rect 371252 241448 371280 241488
rect 370056 241420 371280 241448
rect 372540 241448 372568 241488
rect 372614 241476 372620 241528
rect 372672 241516 372678 241528
rect 373810 241516 373816 241528
rect 372672 241488 373816 241516
rect 372672 241476 372678 241488
rect 373810 241476 373816 241488
rect 373868 241476 373874 241528
rect 374454 241476 374460 241528
rect 374512 241516 374518 241528
rect 375282 241516 375288 241528
rect 374512 241488 375288 241516
rect 374512 241476 374518 241488
rect 375282 241476 375288 241488
rect 375340 241476 375346 241528
rect 379900 241516 379928 241556
rect 381170 241544 381176 241596
rect 381228 241584 381234 241596
rect 384390 241584 384396 241596
rect 381228 241556 384396 241584
rect 381228 241544 381234 241556
rect 384390 241544 384396 241556
rect 384448 241544 384454 241596
rect 386690 241544 386696 241596
rect 386748 241584 386754 241596
rect 388530 241584 388536 241596
rect 386748 241556 388536 241584
rect 386748 241544 386754 241556
rect 388530 241544 388536 241556
rect 388588 241544 388594 241596
rect 388640 241584 388668 241624
rect 390370 241612 390376 241664
rect 390428 241652 390434 241664
rect 392578 241652 392584 241664
rect 390428 241624 392584 241652
rect 390428 241612 390434 241624
rect 392578 241612 392584 241624
rect 392636 241612 392642 241664
rect 393961 241655 394019 241661
rect 393961 241621 393973 241655
rect 394007 241652 394019 241655
rect 456794 241652 456800 241664
rect 394007 241624 456800 241652
rect 394007 241621 394019 241624
rect 393961 241615 394019 241621
rect 456794 241612 456800 241624
rect 456852 241612 456858 241664
rect 452654 241584 452660 241596
rect 388640 241556 452660 241584
rect 452654 241544 452660 241556
rect 452712 241544 452718 241596
rect 375392 241488 379928 241516
rect 375392 241448 375420 241488
rect 379974 241476 379980 241528
rect 380032 241516 380038 241528
rect 380802 241516 380808 241528
rect 380032 241488 380808 241516
rect 380032 241476 380038 241488
rect 380802 241476 380808 241488
rect 380860 241476 380866 241528
rect 382366 241476 382372 241528
rect 382424 241516 382430 241528
rect 383562 241516 383568 241528
rect 382424 241488 383568 241516
rect 382424 241476 382430 241488
rect 383562 241476 383568 241488
rect 383620 241476 383626 241528
rect 383654 241476 383660 241528
rect 383712 241516 383718 241528
rect 384942 241516 384948 241528
rect 383712 241488 384948 241516
rect 383712 241476 383718 241488
rect 384942 241476 384948 241488
rect 385000 241476 385006 241528
rect 385402 241476 385408 241528
rect 385460 241516 385466 241528
rect 386322 241516 386328 241528
rect 385460 241488 386328 241516
rect 385460 241476 385466 241488
rect 386322 241476 386328 241488
rect 386380 241476 386386 241528
rect 387886 241476 387892 241528
rect 387944 241516 387950 241528
rect 388990 241516 388996 241528
rect 387944 241488 388996 241516
rect 387944 241476 387950 241488
rect 388990 241476 388996 241488
rect 389048 241476 389054 241528
rect 390922 241476 390928 241528
rect 390980 241516 390986 241528
rect 391842 241516 391848 241528
rect 390980 241488 391848 241516
rect 390980 241476 390986 241488
rect 391842 241476 391848 241488
rect 391900 241476 391906 241528
rect 393958 241476 393964 241528
rect 394016 241516 394022 241528
rect 395430 241516 395436 241528
rect 394016 241488 395436 241516
rect 394016 241476 394022 241488
rect 395430 241476 395436 241488
rect 395488 241476 395494 241528
rect 396442 241476 396448 241528
rect 396500 241516 396506 241528
rect 397362 241516 397368 241528
rect 396500 241488 397368 241516
rect 396500 241476 396506 241488
rect 397362 241476 397368 241488
rect 397420 241476 397426 241528
rect 398926 241476 398932 241528
rect 398984 241516 398990 241528
rect 400122 241516 400128 241528
rect 398984 241488 400128 241516
rect 398984 241476 398990 241488
rect 400122 241476 400128 241488
rect 400180 241476 400186 241528
rect 400766 241476 400772 241528
rect 400824 241516 400830 241528
rect 401502 241516 401508 241528
rect 400824 241488 401508 241516
rect 400824 241476 400830 241488
rect 401502 241476 401508 241488
rect 401560 241476 401566 241528
rect 401962 241476 401968 241528
rect 402020 241516 402026 241528
rect 402790 241516 402796 241528
rect 402020 241488 402796 241516
rect 402020 241476 402026 241488
rect 402790 241476 402796 241488
rect 402848 241476 402854 241528
rect 404354 241476 404360 241528
rect 404412 241516 404418 241528
rect 405642 241516 405648 241528
rect 404412 241488 405648 241516
rect 404412 241476 404418 241488
rect 405642 241476 405648 241488
rect 405700 241476 405706 241528
rect 406194 241476 406200 241528
rect 406252 241516 406258 241528
rect 407022 241516 407028 241528
rect 406252 241488 407028 241516
rect 406252 241476 406258 241488
rect 407022 241476 407028 241488
rect 407080 241476 407086 241528
rect 407482 241476 407488 241528
rect 407540 241516 407546 241528
rect 408310 241516 408316 241528
rect 407540 241488 408316 241516
rect 407540 241476 407546 241488
rect 408310 241476 408316 241488
rect 408368 241476 408374 241528
rect 409874 241476 409880 241528
rect 409932 241516 409938 241528
rect 411162 241516 411168 241528
rect 409932 241488 411168 241516
rect 409932 241476 409938 241488
rect 411162 241476 411168 241488
rect 411220 241476 411226 241528
rect 411254 241476 411260 241528
rect 411312 241516 411318 241528
rect 411898 241516 411904 241528
rect 411312 241488 411904 241516
rect 411312 241476 411318 241488
rect 411898 241476 411904 241488
rect 411956 241476 411962 241528
rect 412358 241476 412364 241528
rect 412416 241516 412422 241528
rect 418341 241519 418399 241525
rect 418341 241516 418353 241519
rect 412416 241488 418353 241516
rect 412416 241476 412422 241488
rect 418341 241485 418353 241488
rect 418387 241485 418399 241519
rect 418341 241479 418399 241485
rect 418430 241476 418436 241528
rect 418488 241516 418494 241528
rect 419442 241516 419448 241528
rect 418488 241488 419448 241516
rect 418488 241476 418494 241488
rect 419442 241476 419448 241488
rect 419500 241476 419506 241528
rect 419537 241519 419595 241525
rect 419537 241485 419549 241519
rect 419583 241516 419595 241519
rect 419583 241488 420868 241516
rect 419583 241485 419595 241488
rect 419537 241479 419595 241485
rect 372540 241420 375420 241448
rect 420840 241448 420868 241488
rect 420914 241476 420920 241528
rect 420972 241516 420978 241528
rect 422110 241516 422116 241528
rect 420972 241488 422116 241516
rect 420972 241476 420978 241488
rect 422110 241476 422116 241488
rect 422168 241476 422174 241528
rect 423858 241516 423864 241528
rect 422220 241488 423864 241516
rect 422220 241448 422248 241488
rect 423858 241476 423864 241488
rect 423916 241476 423922 241528
rect 423950 241476 423956 241528
rect 424008 241516 424014 241528
rect 424778 241516 424784 241528
rect 424008 241488 424784 241516
rect 424008 241476 424014 241488
rect 424778 241476 424784 241488
rect 424836 241476 424842 241528
rect 425790 241476 425796 241528
rect 425848 241516 425854 241528
rect 426342 241516 426348 241528
rect 425848 241488 426348 241516
rect 425848 241476 425854 241488
rect 426342 241476 426348 241488
rect 426400 241476 426406 241528
rect 426986 241476 426992 241528
rect 427044 241516 427050 241528
rect 427722 241516 427728 241528
rect 427044 241488 427728 241516
rect 427044 241476 427050 241488
rect 427722 241476 427728 241488
rect 427780 241476 427786 241528
rect 428182 241476 428188 241528
rect 428240 241516 428246 241528
rect 429102 241516 429108 241528
rect 428240 241488 429108 241516
rect 428240 241476 428246 241488
rect 429102 241476 429108 241488
rect 429160 241476 429166 241528
rect 429470 241476 429476 241528
rect 429528 241516 429534 241528
rect 430482 241516 430488 241528
rect 429528 241488 430488 241516
rect 429528 241476 429534 241488
rect 430482 241476 430488 241488
rect 430540 241476 430546 241528
rect 430666 241476 430672 241528
rect 430724 241516 430730 241528
rect 430724 241488 431632 241516
rect 430724 241476 430730 241488
rect 423214 241448 423220 241460
rect 420840 241420 422248 241448
rect 423175 241420 423220 241448
rect 423214 241408 423220 241420
rect 423272 241408 423278 241460
rect 431604 241380 431632 241488
rect 431678 241476 431684 241528
rect 431736 241516 431742 241528
rect 431862 241516 431868 241528
rect 431736 241488 431868 241516
rect 431736 241476 431742 241488
rect 431862 241476 431868 241488
rect 431920 241476 431926 241528
rect 433702 241476 433708 241528
rect 433760 241516 433766 241528
rect 434530 241516 434536 241528
rect 433760 241488 434536 241516
rect 433760 241476 433766 241488
rect 434530 241476 434536 241488
rect 434588 241476 434594 241528
rect 434898 241476 434904 241528
rect 434956 241516 434962 241528
rect 436002 241516 436008 241528
rect 434956 241488 436008 241516
rect 434956 241476 434962 241488
rect 436002 241476 436008 241488
rect 436060 241476 436066 241528
rect 436738 241476 436744 241528
rect 436796 241516 436802 241528
rect 437382 241516 437388 241528
rect 436796 241488 437388 241516
rect 436796 241476 436802 241488
rect 437382 241476 437388 241488
rect 437440 241476 437446 241528
rect 438026 241476 438032 241528
rect 438084 241516 438090 241528
rect 438762 241516 438768 241528
rect 438084 241488 438768 241516
rect 438084 241476 438090 241488
rect 438762 241476 438768 241488
rect 438820 241476 438826 241528
rect 439222 241476 439228 241528
rect 439280 241516 439286 241528
rect 440142 241516 440148 241528
rect 439280 241488 440148 241516
rect 439280 241476 439286 241488
rect 440142 241476 440148 241488
rect 440200 241476 440206 241528
rect 440234 241476 440240 241528
rect 440292 241516 440298 241528
rect 527818 241516 527824 241528
rect 440292 241488 527824 241516
rect 440292 241476 440298 241488
rect 527818 241476 527824 241488
rect 527876 241476 527882 241528
rect 431862 241380 431868 241392
rect 431604 241352 431868 241380
rect 431862 241340 431868 241352
rect 431920 241340 431926 241392
rect 237653 239411 237711 239417
rect 237653 239377 237665 239411
rect 237699 239408 237711 239411
rect 237742 239408 237748 239420
rect 237699 239380 237748 239408
rect 237699 239377 237711 239380
rect 237653 239371 237711 239377
rect 237742 239368 237748 239380
rect 237800 239368 237806 239420
rect 149054 239300 149060 239352
rect 149112 239340 149118 239352
rect 149974 239340 149980 239352
rect 149112 239312 149980 239340
rect 149112 239300 149118 239312
rect 149974 239300 149980 239312
rect 150032 239300 150038 239352
rect 150710 239300 150716 239352
rect 150768 239340 150774 239352
rect 151170 239340 151176 239352
rect 150768 239312 151176 239340
rect 150768 239300 150774 239312
rect 151170 239300 151176 239312
rect 151228 239300 151234 239352
rect 158714 239300 158720 239352
rect 158772 239340 158778 239352
rect 159726 239340 159732 239352
rect 158772 239312 159732 239340
rect 158772 239300 158778 239312
rect 159726 239300 159732 239312
rect 159784 239300 159790 239352
rect 164326 239300 164332 239352
rect 164384 239340 164390 239352
rect 165246 239340 165252 239352
rect 164384 239312 165252 239340
rect 164384 239300 164390 239312
rect 165246 239300 165252 239312
rect 165304 239300 165310 239352
rect 166994 239300 167000 239352
rect 167052 239340 167058 239352
rect 167638 239340 167644 239352
rect 167052 239312 167644 239340
rect 167052 239300 167058 239312
rect 167638 239300 167644 239312
rect 167696 239300 167702 239352
rect 171134 239300 171140 239352
rect 171192 239340 171198 239352
rect 171870 239340 171876 239352
rect 171192 239312 171876 239340
rect 171192 239300 171198 239312
rect 171870 239300 171876 239312
rect 171928 239300 171934 239352
rect 190546 239300 190552 239352
rect 190604 239340 190610 239352
rect 191374 239340 191380 239352
rect 190604 239312 191380 239340
rect 190604 239300 190610 239312
rect 191374 239300 191380 239312
rect 191432 239300 191438 239352
rect 196066 239300 196072 239352
rect 196124 239340 196130 239352
rect 196894 239340 196900 239352
rect 196124 239312 196900 239340
rect 196124 239300 196130 239312
rect 196894 239300 196900 239312
rect 196952 239300 196958 239352
rect 201586 239300 201592 239352
rect 201644 239340 201650 239352
rect 202414 239340 202420 239352
rect 201644 239312 202420 239340
rect 201644 239300 201650 239312
rect 202414 239300 202420 239312
rect 202472 239300 202478 239352
rect 212626 239300 212632 239352
rect 212684 239340 212690 239352
rect 213454 239340 213460 239352
rect 212684 239312 213460 239340
rect 212684 239300 212690 239312
rect 213454 239300 213460 239312
rect 213512 239300 213518 239352
rect 215294 239300 215300 239352
rect 215352 239340 215358 239352
rect 215846 239340 215852 239352
rect 215352 239312 215852 239340
rect 215352 239300 215358 239312
rect 215846 239300 215852 239312
rect 215904 239300 215910 239352
rect 220814 239300 220820 239352
rect 220872 239340 220878 239352
rect 221366 239340 221372 239352
rect 220872 239312 221372 239340
rect 220872 239300 220878 239312
rect 221366 239300 221372 239312
rect 221424 239300 221430 239352
rect 222194 239300 222200 239352
rect 222252 239340 222258 239352
rect 223206 239340 223212 239352
rect 222252 239312 223212 239340
rect 222252 239300 222258 239312
rect 223206 239300 223212 239312
rect 223264 239300 223270 239352
rect 227806 239300 227812 239352
rect 227864 239340 227870 239352
rect 228726 239340 228732 239352
rect 227864 239312 228732 239340
rect 227864 239300 227870 239312
rect 228726 239300 228732 239312
rect 228784 239300 228790 239352
rect 230474 239300 230480 239352
rect 230532 239340 230538 239352
rect 231118 239340 231124 239352
rect 230532 239312 231124 239340
rect 230532 239300 230538 239312
rect 231118 239300 231124 239312
rect 231176 239300 231182 239352
rect 231854 239300 231860 239352
rect 231912 239340 231918 239352
rect 232406 239340 232412 239352
rect 231912 239312 232412 239340
rect 231912 239300 231918 239312
rect 232406 239300 232412 239312
rect 232464 239300 232470 239352
rect 233326 239300 233332 239352
rect 233384 239340 233390 239352
rect 234246 239340 234252 239352
rect 233384 239312 234252 239340
rect 233384 239300 233390 239312
rect 234246 239300 234252 239312
rect 234304 239300 234310 239352
rect 241514 239300 241520 239352
rect 241572 239340 241578 239352
rect 242158 239340 242164 239352
rect 241572 239312 242164 239340
rect 241572 239300 241578 239312
rect 242158 239300 242164 239312
rect 242216 239300 242222 239352
rect 244366 239300 244372 239352
rect 244424 239340 244430 239352
rect 244550 239340 244556 239352
rect 244424 239312 244556 239340
rect 244424 239300 244430 239312
rect 244550 239300 244556 239312
rect 244608 239300 244614 239352
rect 247218 239300 247224 239352
rect 247276 239340 247282 239352
rect 247770 239340 247776 239352
rect 247276 239312 247776 239340
rect 247276 239300 247282 239312
rect 247770 239300 247776 239312
rect 247828 239300 247834 239352
rect 249886 239300 249892 239352
rect 249944 239340 249950 239352
rect 250070 239340 250076 239352
rect 249944 239312 250076 239340
rect 249944 239300 249950 239312
rect 250070 239300 250076 239312
rect 250128 239300 250134 239352
rect 270494 239300 270500 239352
rect 270552 239340 270558 239352
rect 271506 239340 271512 239352
rect 270552 239312 271512 239340
rect 270552 239300 270558 239312
rect 271506 239300 271512 239312
rect 271564 239300 271570 239352
rect 272058 239300 272064 239352
rect 272116 239340 272122 239352
rect 272794 239340 272800 239352
rect 272116 239312 272800 239340
rect 272116 239300 272122 239312
rect 272794 239300 272800 239312
rect 272852 239300 272858 239352
rect 276014 239300 276020 239352
rect 276072 239340 276078 239352
rect 276474 239340 276480 239352
rect 276072 239312 276480 239340
rect 276072 239300 276078 239312
rect 276474 239300 276480 239312
rect 276532 239300 276538 239352
rect 423217 239275 423275 239281
rect 423217 239241 423229 239275
rect 423263 239272 423275 239275
rect 423306 239272 423312 239284
rect 423263 239244 423312 239272
rect 423263 239241 423275 239244
rect 423217 239235 423275 239241
rect 423306 239232 423312 239244
rect 423364 239232 423370 239284
rect 269206 238688 269212 238740
rect 269264 238728 269270 238740
rect 269574 238728 269580 238740
rect 269264 238700 269580 238728
rect 269264 238688 269270 238700
rect 269574 238688 269580 238700
rect 269632 238688 269638 238740
rect 3050 237328 3056 237380
rect 3108 237368 3114 237380
rect 10318 237368 10324 237380
rect 3108 237340 10324 237368
rect 3108 237328 3114 237340
rect 10318 237328 10324 237340
rect 10376 237328 10382 237380
rect 222470 236648 222476 236700
rect 222528 236688 222534 236700
rect 222654 236688 222660 236700
rect 222528 236660 222660 236688
rect 222528 236648 222534 236660
rect 222654 236648 222660 236660
rect 222712 236648 222718 236700
rect 223758 236648 223764 236700
rect 223816 236688 223822 236700
rect 224402 236688 224408 236700
rect 223816 236660 224408 236688
rect 223816 236648 223822 236660
rect 224402 236648 224408 236660
rect 224460 236648 224466 236700
rect 233234 236648 233240 236700
rect 233292 236688 233298 236700
rect 233510 236688 233516 236700
rect 233292 236660 233516 236688
rect 233292 236648 233298 236660
rect 233510 236648 233516 236660
rect 233568 236648 233574 236700
rect 194962 235940 194968 235952
rect 194923 235912 194968 235940
rect 194962 235900 194968 235912
rect 195020 235900 195026 235952
rect 265158 234812 265164 234864
rect 265216 234852 265222 234864
rect 265986 234852 265992 234864
rect 265216 234824 265992 234852
rect 265216 234812 265222 234824
rect 265986 234812 265992 234824
rect 266044 234812 266050 234864
rect 164234 234744 164240 234796
rect 164292 234784 164298 234796
rect 164510 234784 164516 234796
rect 164292 234756 164516 234784
rect 164292 234744 164298 234756
rect 164510 234744 164516 234756
rect 164568 234744 164574 234796
rect 403618 234716 403624 234728
rect 403544 234688 403624 234716
rect 245930 234608 245936 234660
rect 245988 234648 245994 234660
rect 246482 234648 246488 234660
rect 245988 234620 246488 234648
rect 245988 234608 245994 234620
rect 246482 234608 246488 234620
rect 246540 234608 246546 234660
rect 350994 234608 351000 234660
rect 351052 234648 351058 234660
rect 351730 234648 351736 234660
rect 351052 234620 351736 234648
rect 351052 234608 351058 234620
rect 351730 234608 351736 234620
rect 351788 234608 351794 234660
rect 403544 234592 403572 234688
rect 403618 234676 403624 234688
rect 403676 234676 403682 234728
rect 270494 234540 270500 234592
rect 270552 234580 270558 234592
rect 270678 234580 270684 234592
rect 270552 234552 270684 234580
rect 270552 234540 270558 234552
rect 270678 234540 270684 234552
rect 270736 234540 270742 234592
rect 403526 234540 403532 234592
rect 403584 234540 403590 234592
rect 185026 231888 185032 231940
rect 185084 231928 185090 231940
rect 185854 231928 185860 231940
rect 185084 231900 185860 231928
rect 185084 231888 185090 231900
rect 185854 231888 185860 231900
rect 185912 231888 185918 231940
rect 163038 231820 163044 231872
rect 163096 231860 163102 231872
rect 163222 231860 163228 231872
rect 163096 231832 163228 231860
rect 163096 231820 163102 231832
rect 163222 231820 163228 231832
rect 163280 231820 163286 231872
rect 174078 231820 174084 231872
rect 174136 231860 174142 231872
rect 174354 231860 174360 231872
rect 174136 231832 174360 231860
rect 174136 231820 174142 231832
rect 174354 231820 174360 231832
rect 174412 231820 174418 231872
rect 179598 231820 179604 231872
rect 179656 231860 179662 231872
rect 179874 231860 179880 231872
rect 179656 231832 179880 231860
rect 179656 231820 179662 231832
rect 179874 231820 179880 231832
rect 179932 231820 179938 231872
rect 185118 231820 185124 231872
rect 185176 231860 185182 231872
rect 185394 231860 185400 231872
rect 185176 231832 185400 231860
rect 185176 231820 185182 231832
rect 185394 231820 185400 231832
rect 185452 231820 185458 231872
rect 190638 231820 190644 231872
rect 190696 231860 190702 231872
rect 190730 231860 190736 231872
rect 190696 231832 190736 231860
rect 190696 231820 190702 231832
rect 190730 231820 190736 231832
rect 190788 231820 190794 231872
rect 196158 231820 196164 231872
rect 196216 231860 196222 231872
rect 196250 231860 196256 231872
rect 196216 231832 196256 231860
rect 196216 231820 196222 231832
rect 196250 231820 196256 231832
rect 196308 231820 196314 231872
rect 198274 231860 198280 231872
rect 198235 231832 198280 231860
rect 198274 231820 198280 231832
rect 198332 231820 198338 231872
rect 208486 231820 208492 231872
rect 208544 231860 208550 231872
rect 209130 231860 209136 231872
rect 208544 231832 209136 231860
rect 208544 231820 208550 231832
rect 209130 231820 209136 231832
rect 209188 231820 209194 231872
rect 211246 231820 211252 231872
rect 211304 231860 211310 231872
rect 211522 231860 211528 231872
rect 211304 231832 211528 231860
rect 211304 231820 211310 231832
rect 211522 231820 211528 231832
rect 211580 231820 211586 231872
rect 225046 231820 225052 231872
rect 225104 231860 225110 231872
rect 225690 231860 225696 231872
rect 225104 231832 225696 231860
rect 225104 231820 225110 231832
rect 225690 231820 225696 231832
rect 225748 231820 225754 231872
rect 226610 231820 226616 231872
rect 226668 231860 226674 231872
rect 226794 231860 226800 231872
rect 226668 231832 226800 231860
rect 226668 231820 226674 231832
rect 226794 231820 226800 231832
rect 226852 231820 226858 231872
rect 229370 231820 229376 231872
rect 229428 231860 229434 231872
rect 229830 231860 229836 231872
rect 229428 231832 229836 231860
rect 229428 231820 229434 231832
rect 229830 231820 229836 231832
rect 229888 231820 229894 231872
rect 234890 231820 234896 231872
rect 234948 231860 234954 231872
rect 235442 231860 235448 231872
rect 234948 231832 235448 231860
rect 234948 231820 234954 231832
rect 235442 231820 235448 231832
rect 235500 231820 235506 231872
rect 236362 231820 236368 231872
rect 236420 231860 236426 231872
rect 236546 231860 236552 231872
rect 236420 231832 236552 231860
rect 236420 231820 236426 231832
rect 236546 231820 236552 231832
rect 236604 231820 236610 231872
rect 237650 231860 237656 231872
rect 237611 231832 237656 231860
rect 237650 231820 237656 231832
rect 237708 231820 237714 231872
rect 239122 231820 239128 231872
rect 239180 231860 239186 231872
rect 239674 231860 239680 231872
rect 239180 231832 239680 231860
rect 239180 231820 239186 231832
rect 239674 231820 239680 231832
rect 239732 231820 239738 231872
rect 303801 231863 303859 231869
rect 303801 231829 303813 231863
rect 303847 231860 303859 231863
rect 303890 231860 303896 231872
rect 303847 231832 303896 231860
rect 303847 231829 303859 231832
rect 303801 231823 303859 231829
rect 303890 231820 303896 231832
rect 303948 231820 303954 231872
rect 393774 231820 393780 231872
rect 393832 231860 393838 231872
rect 393958 231860 393964 231872
rect 393832 231832 393964 231860
rect 393832 231820 393838 231832
rect 393958 231820 393964 231832
rect 394016 231820 394022 231872
rect 403526 231792 403532 231804
rect 403487 231764 403532 231792
rect 403526 231752 403532 231764
rect 403584 231752 403590 231804
rect 207106 230460 207112 230512
rect 207164 230500 207170 230512
rect 207198 230500 207204 230512
rect 207164 230472 207204 230500
rect 207164 230460 207170 230472
rect 207198 230460 207204 230472
rect 207256 230460 207262 230512
rect 238478 230460 238484 230512
rect 238536 230500 238542 230512
rect 238662 230500 238668 230512
rect 238536 230472 238668 230500
rect 238536 230460 238542 230472
rect 238662 230460 238668 230472
rect 238720 230460 238726 230512
rect 248138 230460 248144 230512
rect 248196 230500 248202 230512
rect 248230 230500 248236 230512
rect 248196 230472 248236 230500
rect 248196 230460 248202 230472
rect 248230 230460 248236 230472
rect 248288 230460 248294 230512
rect 374270 230460 374276 230512
rect 374328 230500 374334 230512
rect 374454 230500 374460 230512
rect 374328 230472 374460 230500
rect 374328 230460 374334 230472
rect 374454 230460 374460 230472
rect 374512 230460 374518 230512
rect 449250 229032 449256 229084
rect 449308 229072 449314 229084
rect 580166 229072 580172 229084
rect 449308 229044 580172 229072
rect 449308 229032 449314 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 169938 227032 169944 227044
rect 169899 227004 169944 227032
rect 169938 226992 169944 227004
rect 169996 226992 170002 227044
rect 194962 226352 194968 226364
rect 194923 226324 194968 226352
rect 194962 226312 194968 226324
rect 195020 226312 195026 226364
rect 168650 225060 168656 225072
rect 168576 225032 168656 225060
rect 154850 224992 154856 225004
rect 154811 224964 154856 224992
rect 154850 224952 154856 224964
rect 154908 224952 154914 225004
rect 156138 224992 156144 225004
rect 156099 224964 156144 224992
rect 156138 224952 156144 224964
rect 156196 224952 156202 225004
rect 168576 224936 168604 225032
rect 168650 225020 168656 225032
rect 168708 225020 168714 225072
rect 245930 225060 245936 225072
rect 245856 225032 245936 225060
rect 191926 224992 191932 225004
rect 191887 224964 191932 224992
rect 191926 224952 191932 224964
rect 191984 224952 191990 225004
rect 198274 224952 198280 225004
rect 198332 224952 198338 225004
rect 218422 224992 218428 225004
rect 218256 224964 218428 224992
rect 168558 224884 168564 224936
rect 168616 224884 168622 224936
rect 198292 224856 198320 224952
rect 218256 224936 218284 224964
rect 218422 224952 218428 224964
rect 218480 224952 218486 225004
rect 245856 224936 245884 225032
rect 245930 225020 245936 225032
rect 245988 225020 245994 225072
rect 278869 225063 278927 225069
rect 278869 225029 278881 225063
rect 278915 225060 278927 225063
rect 278958 225060 278964 225072
rect 278915 225032 278964 225060
rect 278915 225029 278927 225032
rect 278869 225023 278927 225029
rect 278958 225020 278964 225032
rect 279016 225020 279022 225072
rect 247218 224952 247224 225004
rect 247276 224952 247282 225004
rect 252646 224952 252652 225004
rect 252704 224992 252710 225004
rect 252830 224992 252836 225004
rect 252704 224964 252836 224992
rect 252704 224952 252710 224964
rect 252830 224952 252836 224964
rect 252888 224952 252894 225004
rect 307846 224952 307852 225004
rect 307904 224992 307910 225004
rect 308030 224992 308036 225004
rect 307904 224964 308036 224992
rect 307904 224952 307910 224964
rect 308030 224952 308036 224964
rect 308088 224952 308094 225004
rect 346118 224952 346124 225004
rect 346176 224992 346182 225004
rect 346302 224992 346308 225004
rect 346176 224964 346308 224992
rect 346176 224952 346182 224964
rect 346302 224952 346308 224964
rect 346360 224952 346366 225004
rect 357158 224952 357164 225004
rect 357216 224992 357222 225004
rect 357342 224992 357348 225004
rect 357216 224964 357348 224992
rect 357216 224952 357222 224964
rect 357342 224952 357348 224964
rect 357400 224952 357406 225004
rect 423214 224992 423220 225004
rect 423175 224964 423220 224992
rect 423214 224952 423220 224964
rect 423272 224952 423278 225004
rect 218238 224884 218244 224936
rect 218296 224884 218302 224936
rect 245838 224884 245844 224936
rect 245896 224884 245902 224936
rect 198366 224856 198372 224868
rect 198292 224828 198372 224856
rect 198366 224816 198372 224828
rect 198424 224816 198430 224868
rect 247236 224856 247264 224952
rect 247310 224856 247316 224868
rect 247236 224828 247316 224856
rect 247310 224816 247316 224828
rect 247368 224816 247374 224868
rect 3326 223524 3332 223576
rect 3384 223564 3390 223576
rect 149698 223564 149704 223576
rect 3384 223536 149704 223564
rect 3384 223524 3390 223536
rect 149698 223524 149704 223536
rect 149756 223524 149762 223576
rect 424686 222232 424692 222284
rect 424744 222272 424750 222284
rect 424778 222272 424784 222284
rect 424744 222244 424784 222272
rect 424744 222232 424750 222244
rect 424778 222232 424784 222244
rect 424836 222232 424842 222284
rect 154850 222204 154856 222216
rect 154811 222176 154856 222204
rect 154850 222164 154856 222176
rect 154908 222164 154914 222216
rect 156138 222204 156144 222216
rect 156099 222176 156144 222204
rect 156138 222164 156144 222176
rect 156196 222164 156202 222216
rect 169941 222207 169999 222213
rect 169941 222173 169953 222207
rect 169987 222204 169999 222207
rect 170030 222204 170036 222216
rect 169987 222176 170036 222204
rect 169987 222173 169999 222176
rect 169941 222167 169999 222173
rect 170030 222164 170036 222176
rect 170088 222164 170094 222216
rect 179598 222164 179604 222216
rect 179656 222204 179662 222216
rect 179782 222204 179788 222216
rect 179656 222176 179788 222204
rect 179656 222164 179662 222176
rect 179782 222164 179788 222176
rect 179840 222164 179846 222216
rect 185118 222164 185124 222216
rect 185176 222204 185182 222216
rect 185302 222204 185308 222216
rect 185176 222176 185308 222204
rect 185176 222164 185182 222176
rect 185302 222164 185308 222176
rect 185360 222164 185366 222216
rect 191926 222204 191932 222216
rect 191887 222176 191932 222204
rect 191926 222164 191932 222176
rect 191984 222164 191990 222216
rect 196158 222164 196164 222216
rect 196216 222204 196222 222216
rect 196342 222204 196348 222216
rect 196216 222176 196348 222204
rect 196216 222164 196222 222176
rect 196342 222164 196348 222176
rect 196400 222164 196406 222216
rect 205818 222164 205824 222216
rect 205876 222204 205882 222216
rect 205910 222204 205916 222216
rect 205876 222176 205916 222204
rect 205876 222164 205882 222176
rect 205910 222164 205916 222176
rect 205968 222164 205974 222216
rect 223850 222204 223856 222216
rect 223811 222176 223856 222204
rect 223850 222164 223856 222176
rect 223908 222164 223914 222216
rect 225138 222204 225144 222216
rect 225099 222176 225144 222204
rect 225138 222164 225144 222176
rect 225196 222164 225202 222216
rect 265158 222164 265164 222216
rect 265216 222204 265222 222216
rect 265342 222204 265348 222216
rect 265216 222176 265348 222204
rect 265216 222164 265222 222176
rect 265342 222164 265348 222176
rect 265400 222164 265406 222216
rect 278866 222204 278872 222216
rect 278827 222176 278872 222204
rect 278866 222164 278872 222176
rect 278924 222164 278930 222216
rect 403529 222207 403587 222213
rect 403529 222173 403541 222207
rect 403575 222204 403587 222207
rect 403710 222204 403716 222216
rect 403575 222176 403716 222204
rect 403575 222173 403587 222176
rect 403529 222167 403587 222173
rect 403710 222164 403716 222176
rect 403768 222164 403774 222216
rect 423214 222204 423220 222216
rect 423175 222176 423220 222204
rect 423214 222164 423220 222176
rect 423272 222164 423278 222216
rect 168558 222096 168564 222148
rect 168616 222096 168622 222148
rect 245838 222096 245844 222148
rect 245896 222096 245902 222148
rect 424686 222136 424692 222148
rect 424647 222108 424692 222136
rect 424686 222096 424692 222108
rect 424744 222096 424750 222148
rect 168576 222000 168604 222096
rect 168650 222000 168656 222012
rect 168576 221972 168656 222000
rect 168650 221960 168656 221972
rect 168708 221960 168714 222012
rect 245856 222000 245884 222096
rect 245930 222000 245936 222012
rect 245856 221972 245936 222000
rect 245930 221960 245936 221972
rect 245988 221960 245994 222012
rect 216766 220872 216772 220924
rect 216824 220912 216830 220924
rect 216858 220912 216864 220924
rect 216824 220884 216864 220912
rect 216824 220872 216830 220884
rect 216858 220872 216864 220884
rect 216916 220872 216922 220924
rect 223850 220844 223856 220856
rect 223811 220816 223856 220844
rect 223850 220804 223856 220816
rect 223908 220804 223914 220856
rect 225138 220844 225144 220856
rect 225099 220816 225144 220844
rect 225138 220804 225144 220816
rect 225196 220804 225202 220856
rect 247954 220804 247960 220856
rect 248012 220844 248018 220856
rect 248322 220844 248328 220856
rect 248012 220816 248328 220844
rect 248012 220804 248018 220816
rect 248322 220804 248328 220816
rect 248380 220804 248386 220856
rect 379054 220804 379060 220856
rect 379112 220844 379118 220856
rect 379238 220844 379244 220856
rect 379112 220816 379244 220844
rect 379112 220804 379118 220816
rect 379238 220804 379244 220816
rect 379296 220804 379302 220856
rect 384574 220804 384580 220856
rect 384632 220844 384638 220856
rect 384850 220844 384856 220856
rect 384632 220816 384856 220844
rect 384632 220804 384638 220816
rect 384850 220804 384856 220816
rect 384908 220804 384914 220856
rect 216766 220736 216772 220788
rect 216824 220776 216830 220788
rect 216950 220776 216956 220788
rect 216824 220748 216956 220776
rect 216824 220736 216830 220748
rect 216950 220736 216956 220748
rect 217008 220736 217014 220788
rect 218238 220736 218244 220788
rect 218296 220776 218302 220788
rect 218330 220776 218336 220788
rect 218296 220748 218336 220776
rect 218296 220736 218302 220748
rect 218330 220736 218336 220748
rect 218388 220736 218394 220788
rect 379146 220736 379152 220788
rect 379204 220776 379210 220788
rect 379330 220776 379336 220788
rect 379204 220748 379336 220776
rect 379204 220736 379210 220748
rect 379330 220736 379336 220748
rect 379388 220736 379394 220788
rect 216950 219416 216956 219428
rect 216911 219388 216956 219416
rect 216950 219376 216956 219388
rect 217008 219376 217014 219428
rect 218241 219419 218299 219425
rect 218241 219385 218253 219419
rect 218287 219416 218299 219419
rect 218330 219416 218336 219428
rect 218287 219388 218336 219416
rect 218287 219385 218299 219388
rect 218241 219379 218299 219385
rect 218330 219376 218336 219388
rect 218388 219376 218394 219428
rect 194502 216588 194508 216640
rect 194560 216628 194566 216640
rect 194962 216628 194968 216640
rect 194560 216600 194968 216628
rect 194560 216588 194566 216600
rect 194962 216588 194968 216600
rect 195020 216588 195026 216640
rect 179509 215407 179567 215413
rect 179509 215373 179521 215407
rect 179555 215404 179567 215407
rect 179598 215404 179604 215416
rect 179555 215376 179604 215404
rect 179555 215373 179567 215376
rect 179509 215367 179567 215373
rect 179598 215364 179604 215376
rect 179656 215364 179662 215416
rect 222562 215404 222568 215416
rect 222488 215376 222568 215404
rect 222488 215280 222516 215376
rect 222562 215364 222568 215376
rect 222620 215364 222626 215416
rect 265069 215407 265127 215413
rect 265069 215373 265081 215407
rect 265115 215404 265127 215407
rect 265158 215404 265164 215416
rect 265115 215376 265164 215404
rect 265115 215373 265127 215376
rect 265069 215367 265127 215373
rect 265158 215364 265164 215376
rect 265216 215364 265222 215416
rect 270589 215407 270647 215413
rect 270589 215373 270601 215407
rect 270635 215404 270647 215407
rect 270678 215404 270684 215416
rect 270635 215376 270684 215404
rect 270635 215373 270647 215376
rect 270589 215367 270647 215373
rect 270678 215364 270684 215376
rect 270736 215364 270742 215416
rect 423214 215364 423220 215416
rect 423272 215364 423278 215416
rect 278866 215296 278872 215348
rect 278924 215296 278930 215348
rect 178218 215268 178224 215280
rect 178179 215240 178224 215268
rect 178218 215228 178224 215240
rect 178276 215228 178282 215280
rect 222470 215228 222476 215280
rect 222528 215228 222534 215280
rect 258166 215228 258172 215280
rect 258224 215268 258230 215280
rect 258350 215268 258356 215280
rect 258224 215240 258356 215268
rect 258224 215228 258230 215240
rect 258350 215228 258356 215240
rect 258408 215228 258414 215280
rect 263778 215268 263784 215280
rect 263739 215240 263784 215268
rect 263778 215228 263784 215240
rect 263836 215228 263842 215280
rect 272058 215268 272064 215280
rect 272019 215240 272064 215268
rect 272058 215228 272064 215240
rect 272116 215228 272122 215280
rect 278884 215212 278912 215296
rect 423232 215280 423260 215364
rect 423214 215228 423220 215280
rect 423272 215228 423278 215280
rect 278866 215160 278872 215212
rect 278924 215160 278930 215212
rect 403526 215160 403532 215212
rect 403584 215200 403590 215212
rect 403710 215200 403716 215212
rect 403584 215172 403716 215200
rect 403584 215160 403590 215172
rect 403710 215160 403716 215172
rect 403768 215160 403774 215212
rect 154758 212508 154764 212560
rect 154816 212548 154822 212560
rect 154850 212548 154856 212560
rect 154816 212520 154856 212548
rect 154816 212508 154822 212520
rect 154850 212508 154856 212520
rect 154908 212508 154914 212560
rect 170030 212508 170036 212560
rect 170088 212548 170094 212560
rect 170122 212548 170128 212560
rect 170088 212520 170128 212548
rect 170088 212508 170094 212520
rect 170122 212508 170128 212520
rect 170180 212508 170186 212560
rect 178218 212548 178224 212560
rect 178179 212520 178224 212548
rect 178218 212508 178224 212520
rect 178276 212508 178282 212560
rect 179506 212548 179512 212560
rect 179467 212520 179512 212548
rect 179506 212508 179512 212520
rect 179564 212508 179570 212560
rect 185118 212508 185124 212560
rect 185176 212548 185182 212560
rect 185210 212548 185216 212560
rect 185176 212520 185216 212548
rect 185176 212508 185182 212520
rect 185210 212508 185216 212520
rect 185268 212508 185274 212560
rect 190730 212508 190736 212560
rect 190788 212548 190794 212560
rect 190914 212548 190920 212560
rect 190788 212520 190920 212548
rect 190788 212508 190794 212520
rect 190914 212508 190920 212520
rect 190972 212508 190978 212560
rect 191742 212508 191748 212560
rect 191800 212548 191806 212560
rect 192018 212548 192024 212560
rect 191800 212520 192024 212548
rect 191800 212508 191806 212520
rect 192018 212508 192024 212520
rect 192076 212508 192082 212560
rect 247310 212508 247316 212560
rect 247368 212548 247374 212560
rect 247402 212548 247408 212560
rect 247368 212520 247408 212548
rect 247368 212508 247374 212520
rect 247402 212508 247408 212520
rect 247460 212508 247466 212560
rect 263778 212548 263784 212560
rect 263739 212520 263784 212548
rect 263778 212508 263784 212520
rect 263836 212508 263842 212560
rect 265066 212548 265072 212560
rect 265027 212520 265072 212548
rect 265066 212508 265072 212520
rect 265124 212508 265130 212560
rect 270586 212548 270592 212560
rect 270547 212520 270592 212548
rect 270586 212508 270592 212520
rect 270644 212508 270650 212560
rect 272058 212548 272064 212560
rect 272019 212520 272064 212548
rect 272058 212508 272064 212520
rect 272116 212508 272122 212560
rect 424689 212551 424747 212557
rect 424689 212517 424701 212551
rect 424735 212548 424747 212551
rect 424778 212548 424784 212560
rect 424735 212520 424784 212548
rect 424735 212517 424747 212520
rect 424689 212511 424747 212517
rect 424778 212508 424784 212520
rect 424836 212508 424842 212560
rect 196250 211216 196256 211268
rect 196308 211256 196314 211268
rect 196342 211256 196348 211268
rect 196308 211228 196348 211256
rect 196308 211216 196314 211228
rect 196342 211216 196348 211228
rect 196400 211216 196406 211268
rect 248138 211148 248144 211200
rect 248196 211188 248202 211200
rect 248230 211188 248236 211200
rect 248196 211160 248236 211188
rect 248196 211148 248202 211160
rect 248230 211148 248236 211160
rect 248288 211148 248294 211200
rect 198182 211080 198188 211132
rect 198240 211120 198246 211132
rect 198366 211120 198372 211132
rect 198240 211092 198372 211120
rect 198240 211080 198246 211092
rect 198366 211080 198372 211092
rect 198424 211080 198430 211132
rect 216950 211120 216956 211132
rect 216911 211092 216956 211120
rect 216950 211080 216956 211092
rect 217008 211080 217014 211132
rect 219526 211080 219532 211132
rect 219584 211080 219590 211132
rect 379146 211080 379152 211132
rect 379204 211120 379210 211132
rect 379238 211120 379244 211132
rect 379204 211092 379244 211120
rect 379204 211080 379210 211092
rect 379238 211080 379244 211092
rect 379296 211080 379302 211132
rect 384666 211120 384672 211132
rect 384627 211092 384672 211120
rect 384666 211080 384672 211092
rect 384724 211080 384730 211132
rect 219544 211052 219572 211080
rect 219618 211052 219624 211064
rect 219544 211024 219624 211052
rect 219618 211012 219624 211024
rect 219676 211012 219682 211064
rect 150802 209788 150808 209840
rect 150860 209828 150866 209840
rect 150894 209828 150900 209840
rect 150860 209800 150900 209828
rect 150860 209788 150866 209800
rect 150894 209788 150900 209800
rect 150952 209788 150958 209840
rect 214006 209828 214012 209840
rect 213967 209800 214012 209828
rect 214006 209788 214012 209800
rect 214064 209788 214070 209840
rect 205910 206252 205916 206304
rect 205968 206292 205974 206304
rect 206094 206292 206100 206304
rect 205968 206264 206100 206292
rect 205968 206252 205974 206264
rect 206094 206252 206100 206264
rect 206152 206252 206158 206304
rect 238478 206252 238484 206304
rect 238536 206292 238542 206304
rect 238662 206292 238668 206304
rect 238536 206264 238668 206292
rect 238536 206252 238542 206264
rect 238662 206252 238668 206264
rect 238720 206252 238726 206304
rect 192018 205708 192024 205760
rect 192076 205708 192082 205760
rect 150802 205640 150808 205692
rect 150860 205640 150866 205692
rect 162854 205640 162860 205692
rect 162912 205680 162918 205692
rect 163038 205680 163044 205692
rect 162912 205652 163044 205680
rect 162912 205640 162918 205652
rect 163038 205640 163044 205652
rect 163096 205640 163102 205692
rect 173894 205640 173900 205692
rect 173952 205680 173958 205692
rect 174078 205680 174084 205692
rect 173952 205652 174084 205680
rect 173952 205640 173958 205652
rect 174078 205640 174084 205652
rect 174136 205640 174142 205692
rect 150820 205556 150848 205640
rect 192036 205624 192064 205708
rect 252646 205640 252652 205692
rect 252704 205680 252710 205692
rect 252830 205680 252836 205692
rect 252704 205652 252836 205680
rect 252704 205640 252710 205652
rect 252830 205640 252836 205652
rect 252888 205640 252894 205692
rect 284294 205640 284300 205692
rect 284352 205680 284358 205692
rect 284478 205680 284484 205692
rect 284352 205652 284484 205680
rect 284352 205640 284358 205652
rect 284478 205640 284484 205652
rect 284536 205640 284542 205692
rect 307846 205640 307852 205692
rect 307904 205680 307910 205692
rect 308030 205680 308036 205692
rect 307904 205652 308036 205680
rect 307904 205640 307910 205652
rect 308030 205640 308036 205652
rect 308088 205640 308094 205692
rect 346118 205640 346124 205692
rect 346176 205680 346182 205692
rect 346302 205680 346308 205692
rect 346176 205652 346308 205680
rect 346176 205640 346182 205652
rect 346302 205640 346308 205652
rect 346360 205640 346366 205692
rect 357158 205640 357164 205692
rect 357216 205680 357222 205692
rect 357342 205680 357348 205692
rect 357216 205652 357348 205680
rect 357216 205640 357222 205652
rect 357342 205640 357348 205652
rect 357400 205640 357406 205692
rect 423214 205680 423220 205692
rect 423175 205652 423220 205680
rect 423214 205640 423220 205652
rect 423272 205640 423278 205692
rect 192018 205572 192024 205624
rect 192076 205572 192082 205624
rect 218238 205612 218244 205624
rect 218199 205584 218244 205612
rect 218238 205572 218244 205584
rect 218296 205572 218302 205624
rect 384666 205612 384672 205624
rect 384627 205584 384672 205612
rect 384666 205572 384672 205584
rect 384724 205572 384730 205624
rect 403526 205572 403532 205624
rect 403584 205612 403590 205624
rect 403710 205612 403716 205624
rect 403584 205584 403716 205612
rect 403584 205572 403590 205584
rect 403710 205572 403716 205584
rect 403768 205572 403774 205624
rect 578050 205572 578056 205624
rect 578108 205612 578114 205624
rect 580810 205612 580816 205624
rect 578108 205584 580816 205612
rect 578108 205572 578114 205584
rect 580810 205572 580816 205584
rect 580868 205572 580874 205624
rect 150802 205504 150808 205556
rect 150860 205504 150866 205556
rect 190454 202852 190460 202904
rect 190512 202892 190518 202904
rect 190638 202892 190644 202904
rect 190512 202864 190644 202892
rect 190512 202852 190518 202864
rect 190638 202852 190644 202864
rect 190696 202852 190702 202904
rect 208486 202852 208492 202904
rect 208544 202892 208550 202904
rect 208578 202892 208584 202904
rect 208544 202864 208584 202892
rect 208544 202852 208550 202864
rect 208578 202852 208584 202864
rect 208636 202852 208642 202904
rect 211246 202852 211252 202904
rect 211304 202892 211310 202904
rect 211338 202892 211344 202904
rect 211304 202864 211344 202892
rect 211304 202852 211310 202864
rect 211338 202852 211344 202864
rect 211396 202852 211402 202904
rect 214006 202892 214012 202904
rect 213967 202864 214012 202892
rect 214006 202852 214012 202864
rect 214064 202852 214070 202904
rect 222470 202852 222476 202904
rect 222528 202892 222534 202904
rect 222562 202892 222568 202904
rect 222528 202864 222568 202892
rect 222528 202852 222534 202864
rect 222562 202852 222568 202864
rect 222620 202852 222626 202904
rect 223850 202852 223856 202904
rect 223908 202892 223914 202904
rect 223942 202892 223948 202904
rect 223908 202864 223948 202892
rect 223908 202852 223914 202864
rect 223942 202852 223948 202864
rect 224000 202852 224006 202904
rect 226518 202852 226524 202904
rect 226576 202892 226582 202904
rect 226610 202892 226616 202904
rect 226576 202864 226616 202892
rect 226576 202852 226582 202864
rect 226610 202852 226616 202864
rect 226668 202852 226674 202904
rect 229278 202852 229284 202904
rect 229336 202892 229342 202904
rect 229370 202892 229376 202904
rect 229336 202864 229376 202892
rect 229336 202852 229342 202864
rect 229370 202852 229376 202864
rect 229428 202852 229434 202904
rect 248138 202852 248144 202904
rect 248196 202892 248202 202904
rect 248322 202892 248328 202904
rect 248196 202864 248328 202892
rect 248196 202852 248202 202864
rect 248322 202852 248328 202864
rect 248380 202852 248386 202904
rect 423214 202892 423220 202904
rect 423175 202864 423220 202892
rect 423214 202852 423220 202864
rect 423272 202852 423278 202904
rect 424594 202852 424600 202904
rect 424652 202892 424658 202904
rect 424686 202892 424692 202904
rect 424652 202864 424692 202892
rect 424652 202852 424658 202864
rect 424686 202852 424692 202864
rect 424744 202852 424750 202904
rect 423214 202756 423220 202768
rect 423175 202728 423220 202756
rect 423214 202716 423220 202728
rect 423272 202716 423278 202768
rect 195974 201560 195980 201612
rect 196032 201600 196038 201612
rect 196250 201600 196256 201612
rect 196032 201572 196256 201600
rect 196032 201560 196038 201572
rect 196250 201560 196256 201572
rect 196308 201560 196314 201612
rect 198366 201560 198372 201612
rect 198424 201560 198430 201612
rect 198384 201476 198412 201560
rect 150713 201467 150771 201473
rect 150713 201433 150725 201467
rect 150759 201464 150771 201467
rect 150802 201464 150808 201476
rect 150759 201436 150808 201464
rect 150759 201433 150771 201436
rect 150713 201427 150771 201433
rect 150802 201424 150808 201436
rect 150860 201424 150866 201476
rect 198366 201424 198372 201476
rect 198424 201424 198430 201476
rect 205910 201424 205916 201476
rect 205968 201424 205974 201476
rect 208394 201424 208400 201476
rect 208452 201464 208458 201476
rect 208578 201464 208584 201476
rect 208452 201436 208584 201464
rect 208452 201424 208458 201436
rect 208578 201424 208584 201436
rect 208636 201424 208642 201476
rect 218238 201464 218244 201476
rect 218199 201436 218244 201464
rect 218238 201424 218244 201436
rect 218296 201424 218302 201476
rect 222562 201424 222568 201476
rect 222620 201464 222626 201476
rect 222654 201464 222660 201476
rect 222620 201436 222660 201464
rect 222620 201424 222626 201436
rect 222654 201424 222660 201436
rect 222712 201424 222718 201476
rect 226610 201424 226616 201476
rect 226668 201464 226674 201476
rect 226794 201464 226800 201476
rect 226668 201436 226800 201464
rect 226668 201424 226674 201436
rect 226794 201424 226800 201436
rect 226852 201424 226858 201476
rect 229370 201424 229376 201476
rect 229428 201464 229434 201476
rect 229462 201464 229468 201476
rect 229428 201436 229468 201464
rect 229428 201424 229434 201436
rect 229462 201424 229468 201436
rect 229520 201424 229526 201476
rect 238478 201424 238484 201476
rect 238536 201464 238542 201476
rect 238662 201464 238668 201476
rect 238536 201436 238668 201464
rect 238536 201424 238542 201436
rect 238662 201424 238668 201436
rect 238720 201424 238726 201476
rect 248141 201467 248199 201473
rect 248141 201433 248153 201467
rect 248187 201464 248199 201467
rect 248322 201464 248328 201476
rect 248187 201436 248328 201464
rect 248187 201433 248199 201436
rect 248141 201427 248199 201433
rect 248322 201424 248328 201436
rect 248380 201424 248386 201476
rect 374270 201424 374276 201476
rect 374328 201464 374334 201476
rect 374454 201464 374460 201476
rect 374328 201436 374460 201464
rect 374328 201424 374334 201436
rect 374454 201424 374460 201436
rect 374512 201424 374518 201476
rect 205928 201396 205956 201424
rect 206002 201396 206008 201408
rect 205928 201368 206008 201396
rect 206002 201356 206008 201368
rect 206060 201356 206066 201408
rect 226702 200064 226708 200116
rect 226760 200104 226766 200116
rect 226794 200104 226800 200116
rect 226760 200076 226800 200104
rect 226760 200064 226766 200076
rect 226794 200064 226800 200076
rect 226852 200064 226858 200116
rect 223850 196092 223856 196104
rect 223776 196064 223856 196092
rect 223776 195968 223804 196064
rect 223850 196052 223856 196064
rect 223908 196052 223914 196104
rect 223758 195916 223764 195968
rect 223816 195916 223822 195968
rect 2774 193876 2780 193928
rect 2832 193916 2838 193928
rect 4982 193916 4988 193928
rect 2832 193888 4988 193916
rect 2832 193876 2838 193888
rect 4982 193876 4988 193888
rect 5040 193876 5046 193928
rect 234890 193304 234896 193316
rect 234816 193276 234896 193304
rect 234816 193248 234844 193276
rect 234890 193264 234896 193276
rect 234948 193264 234954 193316
rect 423217 193307 423275 193313
rect 423217 193273 423229 193307
rect 423263 193304 423275 193307
rect 423306 193304 423312 193316
rect 423263 193276 423312 193304
rect 423263 193273 423275 193276
rect 423217 193267 423275 193273
rect 423306 193264 423312 193276
rect 423364 193264 423370 193316
rect 168650 193196 168656 193248
rect 168708 193236 168714 193248
rect 168834 193236 168840 193248
rect 168708 193208 168840 193236
rect 168708 193196 168714 193208
rect 168834 193196 168840 193208
rect 168892 193196 168898 193248
rect 169754 193196 169760 193248
rect 169812 193236 169818 193248
rect 170030 193236 170036 193248
rect 169812 193208 170036 193236
rect 169812 193196 169818 193208
rect 170030 193196 170036 193208
rect 170088 193196 170094 193248
rect 178218 193196 178224 193248
rect 178276 193236 178282 193248
rect 178402 193236 178408 193248
rect 178276 193208 178408 193236
rect 178276 193196 178282 193208
rect 178402 193196 178408 193208
rect 178460 193196 178466 193248
rect 190454 193196 190460 193248
rect 190512 193236 190518 193248
rect 190730 193236 190736 193248
rect 190512 193208 190736 193236
rect 190512 193196 190518 193208
rect 190730 193196 190736 193208
rect 190788 193196 190794 193248
rect 191834 193196 191840 193248
rect 191892 193236 191898 193248
rect 192018 193236 192024 193248
rect 191892 193208 192024 193236
rect 191892 193196 191898 193208
rect 192018 193196 192024 193208
rect 192076 193196 192082 193248
rect 207014 193196 207020 193248
rect 207072 193236 207078 193248
rect 207198 193236 207204 193248
rect 207072 193208 207204 193236
rect 207072 193196 207078 193208
rect 207198 193196 207204 193208
rect 207256 193196 207262 193248
rect 214006 193196 214012 193248
rect 214064 193236 214070 193248
rect 214098 193236 214104 193248
rect 214064 193208 214104 193236
rect 214064 193196 214070 193208
rect 214098 193196 214104 193208
rect 214156 193196 214162 193248
rect 234798 193196 234804 193248
rect 234856 193196 234862 193248
rect 236270 193196 236276 193248
rect 236328 193236 236334 193248
rect 236454 193236 236460 193248
rect 236328 193208 236460 193236
rect 236328 193196 236334 193208
rect 236454 193196 236460 193208
rect 236512 193196 236518 193248
rect 237558 193196 237564 193248
rect 237616 193236 237622 193248
rect 237742 193236 237748 193248
rect 237616 193208 237748 193236
rect 237616 193196 237622 193208
rect 237742 193196 237748 193208
rect 237800 193196 237806 193248
rect 239030 193196 239036 193248
rect 239088 193236 239094 193248
rect 239214 193236 239220 193248
rect 239088 193208 239220 193236
rect 239088 193196 239094 193208
rect 239214 193196 239220 193208
rect 239272 193196 239278 193248
rect 245930 193196 245936 193248
rect 245988 193236 245994 193248
rect 246114 193236 246120 193248
rect 245988 193208 246120 193236
rect 245988 193196 245994 193208
rect 246114 193196 246120 193208
rect 246172 193196 246178 193248
rect 247034 193196 247040 193248
rect 247092 193236 247098 193248
rect 247310 193236 247316 193248
rect 247092 193208 247316 193236
rect 247092 193196 247098 193208
rect 247310 193196 247316 193208
rect 247368 193196 247374 193248
rect 258074 193196 258080 193248
rect 258132 193236 258138 193248
rect 258350 193236 258356 193248
rect 258132 193208 258356 193236
rect 258132 193196 258138 193208
rect 258350 193196 258356 193208
rect 258408 193196 258414 193248
rect 263594 193196 263600 193248
rect 263652 193236 263658 193248
rect 263778 193236 263784 193248
rect 263652 193208 263784 193236
rect 263652 193196 263658 193208
rect 263778 193196 263784 193208
rect 263836 193196 263842 193248
rect 271874 193196 271880 193248
rect 271932 193236 271938 193248
rect 272058 193236 272064 193248
rect 271932 193208 272064 193236
rect 271932 193196 271938 193208
rect 272058 193196 272064 193208
rect 272116 193196 272122 193248
rect 403802 193196 403808 193248
rect 403860 193236 403866 193248
rect 403986 193236 403992 193248
rect 403860 193208 403992 193236
rect 403860 193196 403866 193208
rect 403986 193196 403992 193208
rect 404044 193196 404050 193248
rect 424502 193196 424508 193248
rect 424560 193236 424566 193248
rect 424778 193236 424784 193248
rect 424560 193208 424784 193236
rect 424560 193196 424566 193208
rect 424778 193196 424784 193208
rect 424836 193196 424842 193248
rect 218241 193171 218299 193177
rect 218241 193137 218253 193171
rect 218287 193168 218299 193171
rect 218330 193168 218336 193180
rect 218287 193140 218336 193168
rect 218287 193137 218299 193140
rect 218241 193131 218299 193137
rect 218330 193128 218336 193140
rect 218388 193128 218394 193180
rect 248138 191876 248144 191888
rect 248099 191848 248144 191876
rect 248138 191836 248144 191848
rect 248196 191836 248202 191888
rect 223758 191768 223764 191820
rect 223816 191808 223822 191820
rect 224034 191808 224040 191820
rect 223816 191780 224040 191808
rect 223816 191768 223822 191780
rect 224034 191768 224040 191780
rect 224092 191768 224098 191820
rect 226426 190408 226432 190460
rect 226484 190448 226490 190460
rect 226794 190448 226800 190460
rect 226484 190420 226800 190448
rect 226484 190408 226490 190420
rect 226794 190408 226800 190420
rect 226852 190408 226858 190460
rect 198274 189048 198280 189100
rect 198332 189088 198338 189100
rect 198366 189088 198372 189100
rect 198332 189060 198372 189088
rect 198332 189048 198338 189060
rect 198366 189048 198372 189060
rect 198424 189048 198430 189100
rect 196253 189023 196311 189029
rect 196253 188989 196265 189023
rect 196299 189020 196311 189023
rect 196342 189020 196348 189032
rect 196299 188992 196348 189020
rect 196299 188989 196311 188992
rect 196253 188983 196311 188989
rect 196342 188980 196348 188992
rect 196400 188980 196406 189032
rect 162854 186328 162860 186380
rect 162912 186368 162918 186380
rect 163038 186368 163044 186380
rect 162912 186340 163044 186368
rect 162912 186328 162918 186340
rect 163038 186328 163044 186340
rect 163096 186328 163102 186380
rect 173894 186328 173900 186380
rect 173952 186368 173958 186380
rect 174078 186368 174084 186380
rect 173952 186340 174084 186368
rect 173952 186328 173958 186340
rect 174078 186328 174084 186340
rect 174136 186328 174142 186380
rect 252646 186328 252652 186380
rect 252704 186368 252710 186380
rect 252830 186368 252836 186380
rect 252704 186340 252836 186368
rect 252704 186328 252710 186340
rect 252830 186328 252836 186340
rect 252888 186328 252894 186380
rect 284294 186328 284300 186380
rect 284352 186368 284358 186380
rect 284478 186368 284484 186380
rect 284352 186340 284484 186368
rect 284352 186328 284358 186340
rect 284478 186328 284484 186340
rect 284536 186328 284542 186380
rect 307846 186328 307852 186380
rect 307904 186368 307910 186380
rect 308030 186368 308036 186380
rect 307904 186340 308036 186368
rect 307904 186328 307910 186340
rect 308030 186328 308036 186340
rect 308088 186328 308094 186380
rect 346118 186328 346124 186380
rect 346176 186368 346182 186380
rect 346302 186368 346308 186380
rect 346176 186340 346308 186368
rect 346176 186328 346182 186340
rect 346302 186328 346308 186340
rect 346360 186328 346366 186380
rect 357158 186328 357164 186380
rect 357216 186368 357222 186380
rect 357342 186368 357348 186380
rect 357216 186340 357348 186368
rect 357216 186328 357222 186340
rect 357342 186328 357348 186340
rect 357400 186328 357406 186380
rect 423125 186371 423183 186377
rect 423125 186337 423137 186371
rect 423171 186368 423183 186371
rect 423214 186368 423220 186380
rect 423171 186340 423220 186368
rect 423171 186337 423183 186340
rect 423125 186331 423183 186337
rect 423214 186328 423220 186340
rect 423272 186328 423278 186380
rect 378870 183608 378876 183660
rect 378928 183648 378934 183660
rect 379054 183648 379060 183660
rect 378928 183620 379060 183648
rect 378928 183608 378934 183620
rect 379054 183608 379060 183620
rect 379112 183608 379118 183660
rect 384574 183608 384580 183660
rect 384632 183648 384638 183660
rect 384666 183648 384672 183660
rect 384632 183620 384672 183648
rect 384632 183608 384638 183620
rect 384666 183608 384672 183620
rect 384724 183608 384730 183660
rect 150713 183583 150771 183589
rect 150713 183549 150725 183583
rect 150759 183580 150771 183583
rect 150802 183580 150808 183592
rect 150759 183552 150808 183580
rect 150759 183549 150771 183552
rect 150713 183543 150771 183549
rect 150802 183540 150808 183552
rect 150860 183540 150866 183592
rect 151814 183540 151820 183592
rect 151872 183580 151878 183592
rect 151998 183580 152004 183592
rect 151872 183552 152004 183580
rect 151872 183540 151878 183552
rect 151998 183540 152004 183552
rect 152056 183540 152062 183592
rect 218238 183540 218244 183592
rect 218296 183580 218302 183592
rect 218422 183580 218428 183592
rect 218296 183552 218428 183580
rect 218296 183540 218302 183552
rect 218422 183540 218428 183552
rect 218480 183540 218486 183592
rect 238478 183540 238484 183592
rect 238536 183580 238542 183592
rect 238662 183580 238668 183592
rect 238536 183552 238668 183580
rect 238536 183540 238542 183552
rect 238662 183540 238668 183552
rect 238720 183540 238726 183592
rect 248138 183540 248144 183592
rect 248196 183580 248202 183592
rect 248322 183580 248328 183592
rect 248196 183552 248328 183580
rect 248196 183540 248202 183552
rect 248322 183540 248328 183552
rect 248380 183540 248386 183592
rect 423122 183580 423128 183592
rect 423083 183552 423128 183580
rect 423122 183540 423128 183552
rect 423180 183540 423186 183592
rect 424594 183540 424600 183592
rect 424652 183580 424658 183592
rect 424686 183580 424692 183592
rect 424652 183552 424692 183580
rect 424652 183540 424658 183552
rect 424686 183540 424692 183552
rect 424744 183540 424750 183592
rect 190730 183512 190736 183524
rect 190691 183484 190736 183512
rect 190730 183472 190736 183484
rect 190788 183472 190794 183524
rect 219526 183512 219532 183524
rect 219487 183484 219532 183512
rect 219526 183472 219532 183484
rect 219584 183472 219590 183524
rect 192018 183444 192024 183456
rect 191979 183416 192024 183444
rect 192018 183404 192024 183416
rect 192076 183404 192082 183456
rect 218238 183444 218244 183456
rect 218199 183416 218244 183444
rect 218238 183404 218244 183416
rect 218296 183404 218302 183456
rect 150713 182155 150771 182161
rect 150713 182121 150725 182155
rect 150759 182152 150771 182155
rect 150802 182152 150808 182164
rect 150759 182124 150808 182152
rect 150759 182121 150771 182124
rect 150713 182115 150771 182121
rect 150802 182112 150808 182124
rect 150860 182112 150866 182164
rect 151998 182112 152004 182164
rect 152056 182152 152062 182164
rect 152182 182152 152188 182164
rect 152056 182124 152188 182152
rect 152056 182112 152062 182124
rect 152182 182112 152188 182124
rect 152240 182112 152246 182164
rect 238481 182155 238539 182161
rect 238481 182121 238493 182155
rect 238527 182152 238539 182155
rect 238662 182152 238668 182164
rect 238527 182124 238668 182152
rect 238527 182121 238539 182124
rect 238481 182115 238539 182121
rect 238662 182112 238668 182124
rect 238720 182112 238726 182164
rect 248138 182112 248144 182164
rect 248196 182152 248202 182164
rect 248322 182152 248328 182164
rect 248196 182124 248328 182152
rect 248196 182112 248202 182124
rect 248322 182112 248328 182124
rect 248380 182112 248386 182164
rect 374270 182112 374276 182164
rect 374328 182152 374334 182164
rect 374454 182152 374460 182164
rect 374328 182124 374460 182152
rect 374328 182112 374334 182124
rect 374454 182112 374460 182124
rect 374512 182112 374518 182164
rect 379054 182112 379060 182164
rect 379112 182152 379118 182164
rect 379330 182152 379336 182164
rect 379112 182124 379336 182152
rect 379112 182112 379118 182124
rect 379330 182112 379336 182124
rect 379388 182112 379394 182164
rect 384574 182152 384580 182164
rect 384535 182124 384580 182152
rect 384574 182112 384580 182124
rect 384632 182112 384638 182164
rect 423122 182112 423128 182164
rect 423180 182152 423186 182164
rect 423214 182152 423220 182164
rect 423180 182124 423220 182152
rect 423180 182112 423186 182124
rect 423214 182112 423220 182124
rect 423272 182112 423278 182164
rect 424502 182152 424508 182164
rect 424463 182124 424508 182152
rect 424502 182112 424508 182124
rect 424560 182112 424566 182164
rect 449158 182112 449164 182164
rect 449216 182152 449222 182164
rect 580166 182152 580172 182164
rect 449216 182124 580172 182152
rect 449216 182112 449222 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 218241 180047 218299 180053
rect 218241 180013 218253 180047
rect 218287 180044 218299 180047
rect 218330 180044 218336 180056
rect 218287 180016 218336 180044
rect 218287 180013 218299 180016
rect 218241 180007 218299 180013
rect 218330 180004 218336 180016
rect 218388 180004 218394 180056
rect 219529 180047 219587 180053
rect 219529 180013 219541 180047
rect 219575 180044 219587 180047
rect 219618 180044 219624 180056
rect 219575 180016 219624 180044
rect 219575 180013 219587 180016
rect 219529 180007 219587 180013
rect 219618 180004 219624 180016
rect 219676 180004 219682 180056
rect 2774 179460 2780 179512
rect 2832 179500 2838 179512
rect 4890 179500 4896 179512
rect 2832 179472 4896 179500
rect 2832 179460 2838 179472
rect 4890 179460 4896 179472
rect 4948 179460 4954 179512
rect 196250 179432 196256 179444
rect 196211 179404 196256 179432
rect 196250 179392 196256 179404
rect 196308 179392 196314 179444
rect 194778 179364 194784 179376
rect 194739 179336 194784 179364
rect 194778 179324 194784 179336
rect 194836 179324 194842 179376
rect 216582 178984 216588 179036
rect 216640 179024 216646 179036
rect 216858 179024 216864 179036
rect 216640 178996 216864 179024
rect 216640 178984 216646 178996
rect 216858 178984 216864 178996
rect 216916 178984 216922 179036
rect 162946 176672 162952 176724
rect 163004 176672 163010 176724
rect 156138 176604 156144 176656
rect 156196 176604 156202 176656
rect 156156 176520 156184 176604
rect 162964 176576 162992 176672
rect 384574 176644 384580 176656
rect 384535 176616 384580 176644
rect 384574 176604 384580 176616
rect 384632 176604 384638 176656
rect 163038 176576 163044 176588
rect 162964 176548 163044 176576
rect 163038 176536 163044 176548
rect 163096 176536 163102 176588
rect 156138 176468 156144 176520
rect 156196 176468 156202 176520
rect 154850 173952 154856 174004
rect 154908 173992 154914 174004
rect 154942 173992 154948 174004
rect 154908 173964 154948 173992
rect 154908 173952 154914 173964
rect 154942 173952 154948 173964
rect 155000 173952 155006 174004
rect 226610 173992 226616 174004
rect 226536 173964 226616 173992
rect 168650 173884 168656 173936
rect 168708 173924 168714 173936
rect 168834 173924 168840 173936
rect 168708 173896 168840 173924
rect 168708 173884 168714 173896
rect 168834 173884 168840 173896
rect 168892 173884 168898 173936
rect 169754 173884 169760 173936
rect 169812 173924 169818 173936
rect 170030 173924 170036 173936
rect 169812 173896 170036 173924
rect 169812 173884 169818 173896
rect 170030 173884 170036 173896
rect 170088 173884 170094 173936
rect 174078 173884 174084 173936
rect 174136 173924 174142 173936
rect 174262 173924 174268 173936
rect 174136 173896 174268 173924
rect 174136 173884 174142 173896
rect 174262 173884 174268 173896
rect 174320 173884 174326 173936
rect 178218 173884 178224 173936
rect 178276 173924 178282 173936
rect 178402 173924 178408 173936
rect 178276 173896 178408 173924
rect 178276 173884 178282 173896
rect 178402 173884 178408 173896
rect 178460 173884 178466 173936
rect 190730 173924 190736 173936
rect 190691 173896 190736 173924
rect 190730 173884 190736 173896
rect 190788 173884 190794 173936
rect 192018 173924 192024 173936
rect 191979 173896 192024 173924
rect 192018 173884 192024 173896
rect 192076 173884 192082 173936
rect 205910 173884 205916 173936
rect 205968 173924 205974 173936
rect 206094 173924 206100 173936
rect 205968 173896 206100 173924
rect 205968 173884 205974 173896
rect 206094 173884 206100 173896
rect 206152 173884 206158 173936
rect 207014 173884 207020 173936
rect 207072 173924 207078 173936
rect 207198 173924 207204 173936
rect 207072 173896 207204 173924
rect 207072 173884 207078 173896
rect 207198 173884 207204 173896
rect 207256 173884 207262 173936
rect 208486 173884 208492 173936
rect 208544 173924 208550 173936
rect 208578 173924 208584 173936
rect 208544 173896 208584 173924
rect 208544 173884 208550 173896
rect 208578 173884 208584 173896
rect 208636 173884 208642 173936
rect 211246 173884 211252 173936
rect 211304 173924 211310 173936
rect 211338 173924 211344 173936
rect 211304 173896 211344 173924
rect 211304 173884 211310 173896
rect 211338 173884 211344 173896
rect 211396 173884 211402 173936
rect 222470 173884 222476 173936
rect 222528 173924 222534 173936
rect 222654 173924 222660 173936
rect 222528 173896 222660 173924
rect 222528 173884 222534 173896
rect 222654 173884 222660 173896
rect 222712 173884 222718 173936
rect 226536 173868 226564 173964
rect 226610 173952 226616 173964
rect 226668 173952 226674 174004
rect 229278 173884 229284 173936
rect 229336 173924 229342 173936
rect 229462 173924 229468 173936
rect 229336 173896 229468 173924
rect 229336 173884 229342 173896
rect 229462 173884 229468 173896
rect 229520 173884 229526 173936
rect 236270 173884 236276 173936
rect 236328 173924 236334 173936
rect 236454 173924 236460 173936
rect 236328 173896 236460 173924
rect 236328 173884 236334 173896
rect 236454 173884 236460 173896
rect 236512 173884 236518 173936
rect 237558 173884 237564 173936
rect 237616 173924 237622 173936
rect 237742 173924 237748 173936
rect 237616 173896 237748 173924
rect 237616 173884 237622 173896
rect 237742 173884 237748 173896
rect 237800 173884 237806 173936
rect 239030 173884 239036 173936
rect 239088 173924 239094 173936
rect 239214 173924 239220 173936
rect 239088 173896 239220 173924
rect 239088 173884 239094 173896
rect 239214 173884 239220 173896
rect 239272 173884 239278 173936
rect 245930 173884 245936 173936
rect 245988 173924 245994 173936
rect 246114 173924 246120 173936
rect 245988 173896 246120 173924
rect 245988 173884 245994 173896
rect 246114 173884 246120 173896
rect 246172 173884 246178 173936
rect 247034 173884 247040 173936
rect 247092 173924 247098 173936
rect 247310 173924 247316 173936
rect 247092 173896 247316 173924
rect 247092 173884 247098 173896
rect 247310 173884 247316 173896
rect 247368 173884 247374 173936
rect 252554 173884 252560 173936
rect 252612 173924 252618 173936
rect 252830 173924 252836 173936
rect 252612 173896 252836 173924
rect 252612 173884 252618 173896
rect 252830 173884 252836 173896
rect 252888 173884 252894 173936
rect 258074 173884 258080 173936
rect 258132 173924 258138 173936
rect 258350 173924 258356 173936
rect 258132 173896 258356 173924
rect 258132 173884 258138 173896
rect 258350 173884 258356 173896
rect 258408 173884 258414 173936
rect 263594 173884 263600 173936
rect 263652 173924 263658 173936
rect 263778 173924 263784 173936
rect 263652 173896 263784 173924
rect 263652 173884 263658 173896
rect 263778 173884 263784 173896
rect 263836 173884 263842 173936
rect 271874 173884 271880 173936
rect 271932 173924 271938 173936
rect 272058 173924 272064 173936
rect 271932 173896 272064 173924
rect 271932 173884 271938 173896
rect 272058 173884 272064 173896
rect 272116 173884 272122 173936
rect 284478 173884 284484 173936
rect 284536 173924 284542 173936
rect 284662 173924 284668 173936
rect 284536 173896 284668 173924
rect 284536 173884 284542 173896
rect 284662 173884 284668 173896
rect 284720 173884 284726 173936
rect 308030 173884 308036 173936
rect 308088 173924 308094 173936
rect 308214 173924 308220 173936
rect 308088 173896 308220 173924
rect 308088 173884 308094 173896
rect 308214 173884 308220 173896
rect 308272 173884 308278 173936
rect 346026 173884 346032 173936
rect 346084 173924 346090 173936
rect 346302 173924 346308 173936
rect 346084 173896 346308 173924
rect 346084 173884 346090 173896
rect 346302 173884 346308 173896
rect 346360 173884 346366 173936
rect 357066 173884 357072 173936
rect 357124 173924 357130 173936
rect 357342 173924 357348 173936
rect 357124 173896 357348 173924
rect 357124 173884 357130 173896
rect 357342 173884 357348 173896
rect 357400 173884 357406 173936
rect 403802 173884 403808 173936
rect 403860 173924 403866 173936
rect 403986 173924 403992 173936
rect 403860 173896 403992 173924
rect 403860 173884 403866 173896
rect 403986 173884 403992 173896
rect 404044 173884 404050 173936
rect 226518 173816 226524 173868
rect 226576 173816 226582 173868
rect 424505 173859 424563 173865
rect 424505 173825 424517 173859
rect 424551 173856 424563 173859
rect 424686 173856 424692 173868
rect 424551 173828 424692 173856
rect 424551 173825 424563 173828
rect 424505 173819 424563 173825
rect 424686 173816 424692 173828
rect 424744 173816 424750 173868
rect 150710 173720 150716 173732
rect 150671 173692 150716 173720
rect 150710 173680 150716 173692
rect 150768 173680 150774 173732
rect 238478 172564 238484 172576
rect 238439 172536 238484 172564
rect 238478 172524 238484 172536
rect 238536 172524 238542 172576
rect 423217 172499 423275 172505
rect 423217 172465 423229 172499
rect 423263 172496 423275 172499
rect 423306 172496 423312 172508
rect 423263 172468 423312 172496
rect 423263 172465 423275 172468
rect 423217 172459 423275 172465
rect 423306 172456 423312 172468
rect 423364 172456 423370 172508
rect 424686 172456 424692 172508
rect 424744 172496 424750 172508
rect 424962 172496 424968 172508
rect 424744 172468 424968 172496
rect 424744 172456 424750 172468
rect 424962 172456 424968 172468
rect 425020 172456 425026 172508
rect 219529 171071 219587 171077
rect 219529 171037 219541 171071
rect 219575 171068 219587 171071
rect 219618 171068 219624 171080
rect 219575 171040 219624 171068
rect 219575 171037 219587 171040
rect 219529 171031 219587 171037
rect 219618 171028 219624 171040
rect 219676 171028 219682 171080
rect 194778 169776 194784 169788
rect 194739 169748 194784 169776
rect 194778 169736 194784 169748
rect 194836 169736 194842 169788
rect 194778 168348 194784 168360
rect 194739 168320 194784 168348
rect 194778 168308 194784 168320
rect 194836 168308 194842 168360
rect 162854 167016 162860 167068
rect 162912 167056 162918 167068
rect 163038 167056 163044 167068
rect 162912 167028 163044 167056
rect 162912 167016 162918 167028
rect 163038 167016 163044 167028
rect 163096 167016 163102 167068
rect 173894 167016 173900 167068
rect 173952 167056 173958 167068
rect 174078 167056 174084 167068
rect 173952 167028 174084 167056
rect 173952 167016 173958 167028
rect 174078 167016 174084 167028
rect 174136 167016 174142 167068
rect 252646 167016 252652 167068
rect 252704 167056 252710 167068
rect 252830 167056 252836 167068
rect 252704 167028 252836 167056
rect 252704 167016 252710 167028
rect 252830 167016 252836 167028
rect 252888 167016 252894 167068
rect 284294 167016 284300 167068
rect 284352 167056 284358 167068
rect 284478 167056 284484 167068
rect 284352 167028 284484 167056
rect 284352 167016 284358 167028
rect 284478 167016 284484 167028
rect 284536 167016 284542 167068
rect 307846 167016 307852 167068
rect 307904 167056 307910 167068
rect 308030 167056 308036 167068
rect 307904 167028 308036 167056
rect 307904 167016 307910 167028
rect 308030 167016 308036 167028
rect 308088 167016 308094 167068
rect 346118 167016 346124 167068
rect 346176 167056 346182 167068
rect 346302 167056 346308 167068
rect 346176 167028 346308 167056
rect 346176 167016 346182 167028
rect 346302 167016 346308 167028
rect 346360 167016 346366 167068
rect 357158 167016 357164 167068
rect 357216 167056 357222 167068
rect 357342 167056 357348 167068
rect 357216 167028 357348 167056
rect 357216 167016 357222 167028
rect 357342 167016 357348 167028
rect 357400 167016 357406 167068
rect 265066 166948 265072 167000
rect 265124 166948 265130 167000
rect 270586 166948 270592 167000
rect 270644 166948 270650 167000
rect 265084 166864 265112 166948
rect 270604 166864 270632 166948
rect 265066 166812 265072 166864
rect 265124 166812 265130 166864
rect 270586 166812 270592 166864
rect 270644 166812 270650 166864
rect 151998 164228 152004 164280
rect 152056 164268 152062 164280
rect 152182 164268 152188 164280
rect 152056 164240 152188 164268
rect 152056 164228 152062 164240
rect 152182 164228 152188 164240
rect 152240 164228 152246 164280
rect 238478 164228 238484 164280
rect 238536 164268 238542 164280
rect 238662 164268 238668 164280
rect 238536 164240 238668 164268
rect 238536 164228 238542 164240
rect 238662 164228 238668 164240
rect 238720 164228 238726 164280
rect 379146 164228 379152 164280
rect 379204 164268 379210 164280
rect 379330 164268 379336 164280
rect 379204 164240 379336 164268
rect 379204 164228 379210 164240
rect 379330 164228 379336 164240
rect 379388 164228 379394 164280
rect 156138 164200 156144 164212
rect 156099 164172 156144 164200
rect 156138 164160 156144 164172
rect 156196 164160 156202 164212
rect 169938 164160 169944 164212
rect 169996 164200 170002 164212
rect 170030 164200 170036 164212
rect 169996 164172 170036 164200
rect 169996 164160 170002 164172
rect 170030 164160 170036 164172
rect 170088 164160 170094 164212
rect 173986 164200 173992 164212
rect 173947 164172 173992 164200
rect 173986 164160 173992 164172
rect 174044 164160 174050 164212
rect 178218 164160 178224 164212
rect 178276 164200 178282 164212
rect 178402 164200 178408 164212
rect 178276 164172 178408 164200
rect 178276 164160 178282 164172
rect 178402 164160 178408 164172
rect 178460 164160 178466 164212
rect 236270 164200 236276 164212
rect 236231 164172 236276 164200
rect 236270 164160 236276 164172
rect 236328 164160 236334 164212
rect 237558 164200 237564 164212
rect 237519 164172 237564 164200
rect 237558 164160 237564 164172
rect 237616 164160 237622 164212
rect 239030 164160 239036 164212
rect 239088 164200 239094 164212
rect 239122 164200 239128 164212
rect 239088 164172 239128 164200
rect 239088 164160 239094 164172
rect 239122 164160 239128 164172
rect 239180 164160 239186 164212
rect 247034 164160 247040 164212
rect 247092 164200 247098 164212
rect 247218 164200 247224 164212
rect 247092 164172 247224 164200
rect 247092 164160 247098 164172
rect 247218 164160 247224 164172
rect 247276 164160 247282 164212
rect 252738 164200 252744 164212
rect 252699 164172 252744 164200
rect 252738 164160 252744 164172
rect 252796 164160 252802 164212
rect 258074 164160 258080 164212
rect 258132 164200 258138 164212
rect 258258 164200 258264 164212
rect 258132 164172 258264 164200
rect 258132 164160 258138 164172
rect 258258 164160 258264 164172
rect 258316 164160 258322 164212
rect 284386 164200 284392 164212
rect 284347 164172 284392 164200
rect 284386 164160 284392 164172
rect 284444 164160 284450 164212
rect 307938 164200 307944 164212
rect 307899 164172 307944 164200
rect 307938 164160 307944 164172
rect 307996 164160 308002 164212
rect 346210 164200 346216 164212
rect 346171 164172 346216 164200
rect 346210 164160 346216 164172
rect 346268 164160 346274 164212
rect 357250 164200 357256 164212
rect 357211 164172 357256 164200
rect 357250 164160 357256 164172
rect 357308 164160 357314 164212
rect 403526 164160 403532 164212
rect 403584 164200 403590 164212
rect 403710 164200 403716 164212
rect 403584 164172 403716 164200
rect 403584 164160 403590 164172
rect 403710 164160 403716 164172
rect 403768 164160 403774 164212
rect 196250 162868 196256 162920
rect 196308 162868 196314 162920
rect 423214 162908 423220 162920
rect 423175 162880 423220 162908
rect 423214 162868 423220 162880
rect 423272 162868 423278 162920
rect 190454 162800 190460 162852
rect 190512 162840 190518 162852
rect 190638 162840 190644 162852
rect 190512 162812 190644 162840
rect 190512 162800 190518 162812
rect 190638 162800 190644 162812
rect 190696 162800 190702 162852
rect 196268 162784 196296 162868
rect 198274 162800 198280 162852
rect 198332 162840 198338 162852
rect 198366 162840 198372 162852
rect 198332 162812 198372 162840
rect 198332 162800 198338 162812
rect 198366 162800 198372 162812
rect 198424 162800 198430 162852
rect 206002 162840 206008 162852
rect 205963 162812 206008 162840
rect 206002 162800 206008 162812
rect 206060 162800 206066 162852
rect 238386 162800 238392 162852
rect 238444 162840 238450 162852
rect 238662 162840 238668 162852
rect 238444 162812 238668 162840
rect 238444 162800 238450 162812
rect 238662 162800 238668 162812
rect 238720 162800 238726 162852
rect 248322 162840 248328 162852
rect 248283 162812 248328 162840
rect 248322 162800 248328 162812
rect 248380 162800 248386 162852
rect 265066 162800 265072 162852
rect 265124 162840 265130 162852
rect 265250 162840 265256 162852
rect 265124 162812 265256 162840
rect 265124 162800 265130 162812
rect 265250 162800 265256 162812
rect 265308 162800 265314 162852
rect 270586 162800 270592 162852
rect 270644 162840 270650 162852
rect 270770 162840 270776 162852
rect 270644 162812 270776 162840
rect 270644 162800 270650 162812
rect 270770 162800 270776 162812
rect 270828 162800 270834 162852
rect 374270 162840 374276 162852
rect 374231 162812 374276 162840
rect 374270 162800 374276 162812
rect 374328 162800 374334 162852
rect 379054 162840 379060 162852
rect 379015 162812 379060 162840
rect 379054 162800 379060 162812
rect 379112 162800 379118 162852
rect 384574 162840 384580 162852
rect 384535 162812 384580 162840
rect 384574 162800 384580 162812
rect 384632 162800 384638 162852
rect 424686 162840 424692 162852
rect 424647 162812 424692 162840
rect 424686 162800 424692 162812
rect 424744 162800 424750 162852
rect 196250 162732 196256 162784
rect 196308 162732 196314 162784
rect 219526 162432 219532 162444
rect 219487 162404 219532 162432
rect 219526 162392 219532 162404
rect 219584 162392 219590 162444
rect 216766 161412 216772 161424
rect 216727 161384 216772 161412
rect 216766 161372 216772 161384
rect 216824 161372 216830 161424
rect 217962 161372 217968 161424
rect 218020 161412 218026 161424
rect 218238 161412 218244 161424
rect 218020 161384 218244 161412
rect 218020 161372 218026 161384
rect 218238 161372 218244 161384
rect 218296 161372 218302 161424
rect 219526 160052 219532 160064
rect 219487 160024 219532 160052
rect 219526 160012 219532 160024
rect 219584 160012 219590 160064
rect 194781 158763 194839 158769
rect 194781 158729 194793 158763
rect 194827 158760 194839 158763
rect 194870 158760 194876 158772
rect 194827 158732 194876 158760
rect 194827 158729 194839 158732
rect 194781 158723 194839 158729
rect 194870 158720 194876 158732
rect 194928 158720 194934 158772
rect 198277 158695 198335 158701
rect 198277 158661 198289 158695
rect 198323 158692 198335 158695
rect 198366 158692 198372 158704
rect 198323 158664 198372 158692
rect 198323 158661 198335 158664
rect 198277 158655 198335 158661
rect 198366 158652 198372 158664
rect 198424 158652 198430 158704
rect 577958 158652 577964 158704
rect 578016 158692 578022 158704
rect 580074 158692 580080 158704
rect 578016 158664 580080 158692
rect 578016 158652 578022 158664
rect 580074 158652 580080 158664
rect 580132 158652 580138 158704
rect 207106 157428 207112 157480
rect 207164 157428 207170 157480
rect 208486 157428 208492 157480
rect 208544 157428 208550 157480
rect 162946 157360 162952 157412
rect 163004 157360 163010 157412
rect 162964 157264 162992 157360
rect 207124 157344 207152 157428
rect 208504 157344 208532 157428
rect 211246 157360 211252 157412
rect 211304 157360 211310 157412
rect 423214 157360 423220 157412
rect 423272 157360 423278 157412
rect 173986 157332 173992 157344
rect 173947 157304 173992 157332
rect 173986 157292 173992 157304
rect 174044 157292 174050 157344
rect 206002 157332 206008 157344
rect 205963 157304 206008 157332
rect 206002 157292 206008 157304
rect 206060 157292 206066 157344
rect 207106 157292 207112 157344
rect 207164 157292 207170 157344
rect 208486 157292 208492 157344
rect 208544 157292 208550 157344
rect 211264 157276 211292 157360
rect 252738 157332 252744 157344
rect 252699 157304 252744 157332
rect 252738 157292 252744 157304
rect 252796 157292 252802 157344
rect 284386 157332 284392 157344
rect 284347 157304 284392 157332
rect 284386 157292 284392 157304
rect 284444 157292 284450 157344
rect 307938 157332 307944 157344
rect 307899 157304 307944 157332
rect 307938 157292 307944 157304
rect 307996 157292 308002 157344
rect 346210 157332 346216 157344
rect 346171 157304 346216 157332
rect 346210 157292 346216 157304
rect 346268 157292 346274 157344
rect 357250 157332 357256 157344
rect 357211 157304 357256 157332
rect 357250 157292 357256 157304
rect 357308 157292 357314 157344
rect 379054 157332 379060 157344
rect 379015 157304 379060 157332
rect 379054 157292 379060 157304
rect 379112 157292 379118 157344
rect 163038 157264 163044 157276
rect 162964 157236 163044 157264
rect 163038 157224 163044 157236
rect 163096 157224 163102 157276
rect 211246 157224 211252 157276
rect 211304 157224 211310 157276
rect 236270 157264 236276 157276
rect 236231 157236 236276 157264
rect 236270 157224 236276 157236
rect 236328 157224 236334 157276
rect 237558 157264 237564 157276
rect 237519 157236 237564 157264
rect 237558 157224 237564 157236
rect 237616 157224 237622 157276
rect 423232 157264 423260 157360
rect 424686 157332 424692 157344
rect 424647 157304 424692 157332
rect 424686 157292 424692 157304
rect 424744 157292 424750 157344
rect 423306 157264 423312 157276
rect 423232 157236 423312 157264
rect 423306 157224 423312 157236
rect 423364 157224 423370 157276
rect 156138 154612 156144 154624
rect 156099 154584 156144 154612
rect 156138 154572 156144 154584
rect 156196 154572 156202 154624
rect 229186 154572 229192 154624
rect 229244 154612 229250 154624
rect 229278 154612 229284 154624
rect 229244 154584 229284 154612
rect 229244 154572 229250 154584
rect 229278 154572 229284 154584
rect 229336 154572 229342 154624
rect 222470 154504 222476 154556
rect 222528 154544 222534 154556
rect 222654 154544 222660 154556
rect 222528 154516 222660 154544
rect 222528 154504 222534 154516
rect 222654 154504 222660 154516
rect 222712 154504 222718 154556
rect 223758 154504 223764 154556
rect 223816 154544 223822 154556
rect 223942 154544 223948 154556
rect 223816 154516 223948 154544
rect 223816 154504 223822 154516
rect 223942 154504 223948 154516
rect 224000 154504 224006 154556
rect 226518 154504 226524 154556
rect 226576 154544 226582 154556
rect 226610 154544 226616 154556
rect 226576 154516 226616 154544
rect 226576 154504 226582 154516
rect 226610 154504 226616 154516
rect 226668 154504 226674 154556
rect 239030 154504 239036 154556
rect 239088 154504 239094 154556
rect 263778 154544 263784 154556
rect 263739 154516 263784 154544
rect 263778 154504 263784 154516
rect 263836 154504 263842 154556
rect 271874 154504 271880 154556
rect 271932 154544 271938 154556
rect 272058 154544 272064 154556
rect 271932 154516 272064 154544
rect 271932 154504 271938 154516
rect 272058 154504 272064 154516
rect 272116 154504 272122 154556
rect 239048 154476 239076 154504
rect 239122 154476 239128 154488
rect 239048 154448 239128 154476
rect 239122 154436 239128 154448
rect 239180 154436 239186 154488
rect 248322 153252 248328 153264
rect 248283 153224 248328 153252
rect 248322 153212 248328 153224
rect 248380 153212 248386 153264
rect 374270 153252 374276 153264
rect 374231 153224 374276 153252
rect 374270 153212 374276 153224
rect 374328 153212 374334 153264
rect 384574 153252 384580 153264
rect 384535 153224 384580 153252
rect 384574 153212 384580 153224
rect 384632 153212 384638 153264
rect 423217 153187 423275 153193
rect 423217 153153 423229 153187
rect 423263 153184 423275 153187
rect 423306 153184 423312 153196
rect 423263 153156 423312 153184
rect 423263 153153 423275 153156
rect 423217 153147 423275 153153
rect 423306 153144 423312 153156
rect 423364 153144 423370 153196
rect 424686 153144 424692 153196
rect 424744 153184 424750 153196
rect 424778 153184 424784 153196
rect 424744 153156 424784 153184
rect 424744 153144 424750 153156
rect 424778 153144 424784 153156
rect 424836 153144 424842 153196
rect 216769 151827 216827 151833
rect 216769 151793 216781 151827
rect 216815 151824 216827 151827
rect 216858 151824 216864 151836
rect 216815 151796 216864 151824
rect 216815 151793 216827 151796
rect 216769 151787 216827 151793
rect 216858 151784 216864 151796
rect 216916 151784 216922 151836
rect 3326 151716 3332 151768
rect 3384 151756 3390 151768
rect 19978 151756 19984 151768
rect 3384 151728 19984 151756
rect 3384 151716 3390 151728
rect 19978 151716 19984 151728
rect 20036 151716 20042 151768
rect 219529 150467 219587 150473
rect 219529 150433 219541 150467
rect 219575 150464 219587 150467
rect 219618 150464 219624 150476
rect 219575 150436 219624 150464
rect 219575 150433 219587 150436
rect 219529 150427 219587 150433
rect 219618 150424 219624 150436
rect 219676 150424 219682 150476
rect 194689 150399 194747 150405
rect 194689 150365 194701 150399
rect 194735 150396 194747 150399
rect 194778 150396 194784 150408
rect 194735 150368 194784 150396
rect 194735 150365 194747 150368
rect 194689 150359 194747 150365
rect 194778 150356 194784 150368
rect 194836 150356 194842 150408
rect 198274 149104 198280 149116
rect 198235 149076 198280 149104
rect 198274 149064 198280 149076
rect 198332 149064 198338 149116
rect 263778 148356 263784 148368
rect 263739 148328 263784 148356
rect 263778 148316 263784 148328
rect 263836 148316 263842 148368
rect 162854 147636 162860 147688
rect 162912 147676 162918 147688
rect 163038 147676 163044 147688
rect 162912 147648 163044 147676
rect 162912 147636 162918 147648
rect 163038 147636 163044 147648
rect 163096 147636 163102 147688
rect 173894 147636 173900 147688
rect 173952 147676 173958 147688
rect 174078 147676 174084 147688
rect 173952 147648 174084 147676
rect 173952 147636 173958 147648
rect 174078 147636 174084 147648
rect 174136 147636 174142 147688
rect 252646 147636 252652 147688
rect 252704 147676 252710 147688
rect 252830 147676 252836 147688
rect 252704 147648 252836 147676
rect 252704 147636 252710 147648
rect 252830 147636 252836 147648
rect 252888 147636 252894 147688
rect 284294 147636 284300 147688
rect 284352 147676 284358 147688
rect 284478 147676 284484 147688
rect 284352 147648 284484 147676
rect 284352 147636 284358 147648
rect 284478 147636 284484 147648
rect 284536 147636 284542 147688
rect 307846 147636 307852 147688
rect 307904 147676 307910 147688
rect 308030 147676 308036 147688
rect 307904 147648 308036 147676
rect 307904 147636 307910 147648
rect 308030 147636 308036 147648
rect 308088 147636 308094 147688
rect 346118 147636 346124 147688
rect 346176 147676 346182 147688
rect 346302 147676 346308 147688
rect 346176 147648 346308 147676
rect 346176 147636 346182 147648
rect 346302 147636 346308 147648
rect 346360 147636 346366 147688
rect 357158 147636 357164 147688
rect 357216 147676 357222 147688
rect 357342 147676 357348 147688
rect 357216 147648 357348 147676
rect 357216 147636 357222 147648
rect 357342 147636 357348 147648
rect 357400 147636 357406 147688
rect 238570 144916 238576 144968
rect 238628 144956 238634 144968
rect 238662 144956 238668 144968
rect 238628 144928 238668 144956
rect 238628 144916 238634 144928
rect 238662 144916 238668 144928
rect 238720 144916 238726 144968
rect 379146 144916 379152 144968
rect 379204 144916 379210 144968
rect 173986 144888 173992 144900
rect 173947 144860 173992 144888
rect 173986 144848 173992 144860
rect 174044 144848 174050 144900
rect 178218 144848 178224 144900
rect 178276 144888 178282 144900
rect 178402 144888 178408 144900
rect 178276 144860 178408 144888
rect 178276 144848 178282 144860
rect 178402 144848 178408 144860
rect 178460 144848 178466 144900
rect 190638 144848 190644 144900
rect 190696 144848 190702 144900
rect 191834 144848 191840 144900
rect 191892 144888 191898 144900
rect 191926 144888 191932 144900
rect 191892 144860 191932 144888
rect 191892 144848 191898 144860
rect 191926 144848 191932 144860
rect 191984 144848 191990 144900
rect 205910 144848 205916 144900
rect 205968 144888 205974 144900
rect 206002 144888 206008 144900
rect 205968 144860 206008 144888
rect 205968 144848 205974 144860
rect 206002 144848 206008 144860
rect 206060 144848 206066 144900
rect 207106 144848 207112 144900
rect 207164 144888 207170 144900
rect 207198 144888 207204 144900
rect 207164 144860 207204 144888
rect 207164 144848 207170 144860
rect 207198 144848 207204 144860
rect 207256 144848 207262 144900
rect 208486 144848 208492 144900
rect 208544 144888 208550 144900
rect 208670 144888 208676 144900
rect 208544 144860 208676 144888
rect 208544 144848 208550 144860
rect 208670 144848 208676 144860
rect 208728 144848 208734 144900
rect 211246 144848 211252 144900
rect 211304 144888 211310 144900
rect 211430 144888 211436 144900
rect 211304 144860 211436 144888
rect 211304 144848 211310 144860
rect 211430 144848 211436 144860
rect 211488 144848 211494 144900
rect 234890 144848 234896 144900
rect 234948 144888 234954 144900
rect 234982 144888 234988 144900
rect 234948 144860 234988 144888
rect 234948 144848 234954 144860
rect 234982 144848 234988 144860
rect 235040 144848 235046 144900
rect 236270 144848 236276 144900
rect 236328 144888 236334 144900
rect 236362 144888 236368 144900
rect 236328 144860 236368 144888
rect 236328 144848 236334 144860
rect 236362 144848 236368 144860
rect 236420 144848 236426 144900
rect 237558 144848 237564 144900
rect 237616 144888 237622 144900
rect 237650 144888 237656 144900
rect 237616 144860 237656 144888
rect 237616 144848 237622 144860
rect 237650 144848 237656 144860
rect 237708 144848 237714 144900
rect 239030 144848 239036 144900
rect 239088 144888 239094 144900
rect 239122 144888 239128 144900
rect 239088 144860 239128 144888
rect 239088 144848 239094 144860
rect 239122 144848 239128 144860
rect 239180 144848 239186 144900
rect 252738 144888 252744 144900
rect 252699 144860 252744 144888
rect 252738 144848 252744 144860
rect 252796 144848 252802 144900
rect 284386 144888 284392 144900
rect 284347 144860 284392 144888
rect 284386 144848 284392 144860
rect 284444 144848 284450 144900
rect 303890 144848 303896 144900
rect 303948 144888 303954 144900
rect 303982 144888 303988 144900
rect 303948 144860 303988 144888
rect 303948 144848 303954 144860
rect 303982 144848 303988 144860
rect 304040 144848 304046 144900
rect 307938 144888 307944 144900
rect 307899 144860 307944 144888
rect 307938 144848 307944 144860
rect 307996 144848 308002 144900
rect 346210 144888 346216 144900
rect 346171 144860 346216 144888
rect 346210 144848 346216 144860
rect 346268 144848 346274 144900
rect 357250 144888 357256 144900
rect 357211 144860 357256 144888
rect 357250 144848 357256 144860
rect 357308 144848 357314 144900
rect 190656 144820 190684 144848
rect 379164 144832 379192 144916
rect 190730 144820 190736 144832
rect 190656 144792 190736 144820
rect 190730 144780 190736 144792
rect 190788 144780 190794 144832
rect 379146 144780 379152 144832
rect 379204 144780 379210 144832
rect 384574 144780 384580 144832
rect 384632 144820 384638 144832
rect 384850 144820 384856 144832
rect 384632 144792 384856 144820
rect 384632 144780 384638 144792
rect 384850 144780 384856 144792
rect 384908 144780 384914 144832
rect 423214 143596 423220 143608
rect 423175 143568 423220 143596
rect 423214 143556 423220 143568
rect 423272 143556 423278 143608
rect 162946 143528 162952 143540
rect 162907 143500 162952 143528
rect 162946 143488 162952 143500
rect 163004 143488 163010 143540
rect 189258 143528 189264 143540
rect 189219 143500 189264 143528
rect 189258 143488 189264 143500
rect 189316 143488 189322 143540
rect 190362 143488 190368 143540
rect 190420 143528 190426 143540
rect 190730 143528 190736 143540
rect 190420 143500 190736 143528
rect 190420 143488 190426 143500
rect 190730 143488 190736 143500
rect 190788 143488 190794 143540
rect 205910 143488 205916 143540
rect 205968 143528 205974 143540
rect 206094 143528 206100 143540
rect 205968 143500 206100 143528
rect 205968 143488 205974 143500
rect 206094 143488 206100 143500
rect 206152 143488 206158 143540
rect 238662 143528 238668 143540
rect 238623 143500 238668 143528
rect 238662 143488 238668 143500
rect 238720 143488 238726 143540
rect 245746 143488 245752 143540
rect 245804 143488 245810 143540
rect 248322 143528 248328 143540
rect 248283 143500 248328 143528
rect 248322 143488 248328 143500
rect 248380 143488 248386 143540
rect 374270 143528 374276 143540
rect 374231 143500 374276 143528
rect 374270 143488 374276 143500
rect 374328 143488 374334 143540
rect 424686 143528 424692 143540
rect 424647 143500 424692 143528
rect 424686 143488 424692 143500
rect 424744 143488 424750 143540
rect 245764 143460 245792 143488
rect 245930 143460 245936 143472
rect 245764 143432 245936 143460
rect 245930 143420 245936 143432
rect 245988 143420 245994 143472
rect 196250 142236 196256 142248
rect 196176 142208 196256 142236
rect 196176 142112 196204 142208
rect 196250 142196 196256 142208
rect 196308 142196 196314 142248
rect 217962 142128 217968 142180
rect 218020 142168 218026 142180
rect 218422 142168 218428 142180
rect 218020 142140 218428 142168
rect 218020 142128 218026 142140
rect 218422 142128 218428 142140
rect 218480 142128 218486 142180
rect 151998 142060 152004 142112
rect 152056 142100 152062 142112
rect 152182 142100 152188 142112
rect 152056 142072 152188 142100
rect 152056 142060 152062 142072
rect 152182 142060 152188 142072
rect 152240 142060 152246 142112
rect 196158 142060 196164 142112
rect 196216 142060 196222 142112
rect 263778 142100 263784 142112
rect 263739 142072 263784 142100
rect 263778 142060 263784 142072
rect 263836 142060 263842 142112
rect 379146 142100 379152 142112
rect 379107 142072 379152 142100
rect 379146 142060 379152 142072
rect 379204 142060 379210 142112
rect 194686 140808 194692 140820
rect 194647 140780 194692 140808
rect 194686 140768 194692 140780
rect 194744 140768 194750 140820
rect 150710 140700 150716 140752
rect 150768 140740 150774 140752
rect 150805 140743 150863 140749
rect 150805 140740 150817 140743
rect 150768 140712 150817 140740
rect 150768 140700 150774 140712
rect 150805 140709 150817 140712
rect 150851 140709 150863 140743
rect 152182 140740 152188 140752
rect 152143 140712 152188 140740
rect 150805 140703 150863 140709
rect 152182 140700 152188 140712
rect 152240 140700 152246 140752
rect 198274 138048 198280 138100
rect 198332 138048 198338 138100
rect 403618 138088 403624 138100
rect 403544 138060 403624 138088
rect 198292 137964 198320 138048
rect 247218 137980 247224 138032
rect 247276 137980 247282 138032
rect 162946 137952 162952 137964
rect 162907 137924 162952 137952
rect 162946 137912 162952 137924
rect 163004 137912 163010 137964
rect 173986 137952 173992 137964
rect 173947 137924 173992 137952
rect 173986 137912 173992 137924
rect 174044 137912 174050 137964
rect 198274 137912 198280 137964
rect 198332 137912 198338 137964
rect 247236 137952 247264 137980
rect 403544 137964 403572 138060
rect 403618 138048 403624 138060
rect 403676 138048 403682 138100
rect 423214 137980 423220 138032
rect 423272 137980 423278 138032
rect 247310 137952 247316 137964
rect 247236 137924 247316 137952
rect 247310 137912 247316 137924
rect 247368 137912 247374 137964
rect 252738 137952 252744 137964
rect 252699 137924 252744 137952
rect 252738 137912 252744 137924
rect 252796 137912 252802 137964
rect 284386 137952 284392 137964
rect 284347 137924 284392 137952
rect 284386 137912 284392 137924
rect 284444 137912 284450 137964
rect 307938 137952 307944 137964
rect 307899 137924 307944 137952
rect 307938 137912 307944 137924
rect 307996 137912 308002 137964
rect 346210 137952 346216 137964
rect 346171 137924 346216 137952
rect 346210 137912 346216 137924
rect 346268 137912 346274 137964
rect 357250 137952 357256 137964
rect 357211 137924 357256 137952
rect 357250 137912 357256 137924
rect 357308 137912 357314 137964
rect 403526 137912 403532 137964
rect 403584 137912 403590 137964
rect 423232 137952 423260 137980
rect 423306 137952 423312 137964
rect 423232 137924 423312 137952
rect 423306 137912 423312 137924
rect 423364 137912 423370 137964
rect 424686 137952 424692 137964
rect 424647 137924 424692 137952
rect 424686 137912 424692 137924
rect 424744 137912 424750 137964
rect 216769 135235 216827 135241
rect 216769 135201 216781 135235
rect 216815 135232 216827 135235
rect 216858 135232 216864 135244
rect 216815 135204 216864 135232
rect 216815 135201 216827 135204
rect 216769 135195 216827 135201
rect 216858 135192 216864 135204
rect 216916 135192 216922 135244
rect 234798 135192 234804 135244
rect 234856 135232 234862 135244
rect 234982 135232 234988 135244
rect 234856 135204 234988 135232
rect 234856 135192 234862 135204
rect 234982 135192 234988 135204
rect 235040 135192 235046 135244
rect 271874 135192 271880 135244
rect 271932 135232 271938 135244
rect 272058 135232 272064 135244
rect 271932 135204 272064 135232
rect 271932 135192 271938 135204
rect 272058 135192 272064 135204
rect 272116 135192 272122 135244
rect 403250 135192 403256 135244
rect 403308 135232 403314 135244
rect 403526 135232 403532 135244
rect 403308 135204 403532 135232
rect 403308 135192 403314 135204
rect 403526 135192 403532 135204
rect 403584 135192 403590 135244
rect 577866 135192 577872 135244
rect 577924 135232 577930 135244
rect 580626 135232 580632 135244
rect 577924 135204 580632 135232
rect 577924 135192 577930 135204
rect 580626 135192 580632 135204
rect 580684 135192 580690 135244
rect 168742 133968 168748 134020
rect 168800 134008 168806 134020
rect 168834 134008 168840 134020
rect 168800 133980 168840 134008
rect 168800 133968 168806 133980
rect 168834 133968 168840 133980
rect 168892 133968 168898 134020
rect 189258 133940 189264 133952
rect 189219 133912 189264 133940
rect 189258 133900 189264 133912
rect 189316 133900 189322 133952
rect 248322 133940 248328 133952
rect 248283 133912 248328 133940
rect 248322 133900 248328 133912
rect 248380 133900 248386 133952
rect 374270 133940 374276 133952
rect 374231 133912 374276 133940
rect 374270 133900 374276 133912
rect 374328 133900 374334 133952
rect 153378 133872 153384 133884
rect 153339 133844 153384 133872
rect 153378 133832 153384 133844
rect 153436 133832 153442 133884
rect 156138 133872 156144 133884
rect 156099 133844 156144 133872
rect 156138 133832 156144 133844
rect 156196 133832 156202 133884
rect 168834 133872 168840 133884
rect 168795 133844 168840 133872
rect 168834 133832 168840 133844
rect 168892 133832 168898 133884
rect 190454 133832 190460 133884
rect 190512 133872 190518 133884
rect 190638 133872 190644 133884
rect 190512 133844 190644 133872
rect 190512 133832 190518 133844
rect 190638 133832 190644 133844
rect 190696 133832 190702 133884
rect 234801 133875 234859 133881
rect 234801 133841 234813 133875
rect 234847 133872 234859 133875
rect 234982 133872 234988 133884
rect 234847 133844 234988 133872
rect 234847 133841 234859 133844
rect 234801 133835 234859 133841
rect 234982 133832 234988 133844
rect 235040 133832 235046 133884
rect 245749 133875 245807 133881
rect 245749 133841 245761 133875
rect 245795 133872 245807 133875
rect 245930 133872 245936 133884
rect 245795 133844 245936 133872
rect 245795 133841 245807 133844
rect 245749 133835 245807 133841
rect 245930 133832 245936 133844
rect 245988 133832 245994 133884
rect 384666 133872 384672 133884
rect 384627 133844 384672 133872
rect 384666 133832 384672 133844
rect 384724 133832 384730 133884
rect 424689 133875 424747 133881
rect 424689 133841 424701 133875
rect 424735 133872 424747 133875
rect 424778 133872 424784 133884
rect 424735 133844 424784 133872
rect 424735 133841 424747 133844
rect 424689 133835 424747 133841
rect 424778 133832 424784 133844
rect 424836 133832 424842 133884
rect 263778 132512 263784 132524
rect 263739 132484 263784 132512
rect 263778 132472 263784 132484
rect 263836 132472 263842 132524
rect 379149 132515 379207 132521
rect 379149 132481 379161 132515
rect 379195 132512 379207 132515
rect 379238 132512 379244 132524
rect 379195 132484 379244 132512
rect 379195 132481 379207 132484
rect 379149 132475 379207 132481
rect 379238 132472 379244 132484
rect 379296 132472 379302 132524
rect 192018 132444 192024 132456
rect 191979 132416 192024 132444
rect 192018 132404 192024 132416
rect 192076 132404 192082 132456
rect 379149 132379 379207 132385
rect 379149 132345 379161 132379
rect 379195 132376 379207 132379
rect 379238 132376 379244 132388
rect 379195 132348 379244 132376
rect 379195 132345 379207 132348
rect 379149 132339 379207 132345
rect 379238 132336 379244 132348
rect 379296 132336 379302 132388
rect 150802 131112 150808 131164
rect 150860 131152 150866 131164
rect 152182 131152 152188 131164
rect 150860 131124 150905 131152
rect 152143 131124 152188 131152
rect 150860 131112 150866 131124
rect 152182 131112 152188 131124
rect 152240 131112 152246 131164
rect 216766 129724 216772 129736
rect 216727 129696 216772 129724
rect 216766 129684 216772 129696
rect 216824 129684 216830 129736
rect 423306 129004 423312 129056
rect 423364 129044 423370 129056
rect 423490 129044 423496 129056
rect 423364 129016 423496 129044
rect 423364 129004 423370 129016
rect 423490 129004 423496 129016
rect 423548 129004 423554 129056
rect 218330 128432 218336 128444
rect 218256 128404 218336 128432
rect 162854 128324 162860 128376
rect 162912 128364 162918 128376
rect 163038 128364 163044 128376
rect 162912 128336 163044 128364
rect 162912 128324 162918 128336
rect 163038 128324 163044 128336
rect 163096 128324 163102 128376
rect 173894 128324 173900 128376
rect 173952 128364 173958 128376
rect 174078 128364 174084 128376
rect 173952 128336 174084 128364
rect 173952 128324 173958 128336
rect 174078 128324 174084 128336
rect 174136 128324 174142 128376
rect 218256 128308 218284 128404
rect 218330 128392 218336 128404
rect 218388 128392 218394 128444
rect 252646 128324 252652 128376
rect 252704 128364 252710 128376
rect 252830 128364 252836 128376
rect 252704 128336 252836 128364
rect 252704 128324 252710 128336
rect 252830 128324 252836 128336
rect 252888 128324 252894 128376
rect 284294 128324 284300 128376
rect 284352 128364 284358 128376
rect 284478 128364 284484 128376
rect 284352 128336 284484 128364
rect 284352 128324 284358 128336
rect 284478 128324 284484 128336
rect 284536 128324 284542 128376
rect 307846 128324 307852 128376
rect 307904 128364 307910 128376
rect 308030 128364 308036 128376
rect 307904 128336 308036 128364
rect 307904 128324 307910 128336
rect 308030 128324 308036 128336
rect 308088 128324 308094 128376
rect 346118 128324 346124 128376
rect 346176 128364 346182 128376
rect 346302 128364 346308 128376
rect 346176 128336 346308 128364
rect 346176 128324 346182 128336
rect 346302 128324 346308 128336
rect 346360 128324 346366 128376
rect 357158 128324 357164 128376
rect 357216 128364 357222 128376
rect 357342 128364 357348 128376
rect 357216 128336 357348 128364
rect 357216 128324 357222 128336
rect 357342 128324 357348 128336
rect 357400 128324 357406 128376
rect 218238 128256 218244 128308
rect 218296 128256 218302 128308
rect 384666 127820 384672 127832
rect 384627 127792 384672 127820
rect 384666 127780 384672 127792
rect 384724 127780 384730 127832
rect 238662 125644 238668 125656
rect 238623 125616 238668 125644
rect 238662 125604 238668 125616
rect 238720 125604 238726 125656
rect 173986 125576 173992 125588
rect 173947 125548 173992 125576
rect 173986 125536 173992 125548
rect 174044 125536 174050 125588
rect 178218 125576 178224 125588
rect 178179 125548 178224 125576
rect 178218 125536 178224 125548
rect 178276 125536 178282 125588
rect 205818 125536 205824 125588
rect 205876 125576 205882 125588
rect 206002 125576 206008 125588
rect 205876 125548 206008 125576
rect 205876 125536 205882 125548
rect 206002 125536 206008 125548
rect 206060 125536 206066 125588
rect 208486 125536 208492 125588
rect 208544 125576 208550 125588
rect 208670 125576 208676 125588
rect 208544 125548 208676 125576
rect 208544 125536 208550 125548
rect 208670 125536 208676 125548
rect 208728 125536 208734 125588
rect 211246 125536 211252 125588
rect 211304 125536 211310 125588
rect 216766 125536 216772 125588
rect 216824 125576 216830 125588
rect 216950 125576 216956 125588
rect 216824 125548 216956 125576
rect 216824 125536 216830 125548
rect 216950 125536 216956 125548
rect 217008 125536 217014 125588
rect 218238 125536 218244 125588
rect 218296 125576 218302 125588
rect 218422 125576 218428 125588
rect 218296 125548 218428 125576
rect 218296 125536 218302 125548
rect 218422 125536 218428 125548
rect 218480 125536 218486 125588
rect 219526 125536 219532 125588
rect 219584 125576 219590 125588
rect 219710 125576 219716 125588
rect 219584 125548 219716 125576
rect 219584 125536 219590 125548
rect 219710 125536 219716 125548
rect 219768 125536 219774 125588
rect 238938 125536 238944 125588
rect 238996 125576 239002 125588
rect 239122 125576 239128 125588
rect 238996 125548 239128 125576
rect 238996 125536 239002 125548
rect 239122 125536 239128 125548
rect 239180 125536 239186 125588
rect 252738 125576 252744 125588
rect 252699 125548 252744 125576
rect 252738 125536 252744 125548
rect 252796 125536 252802 125588
rect 284386 125576 284392 125588
rect 284347 125548 284392 125576
rect 284386 125536 284392 125548
rect 284444 125536 284450 125588
rect 303890 125536 303896 125588
rect 303948 125576 303954 125588
rect 303982 125576 303988 125588
rect 303948 125548 303988 125576
rect 303948 125536 303954 125548
rect 303982 125536 303988 125548
rect 304040 125536 304046 125588
rect 307938 125576 307944 125588
rect 307899 125548 307944 125576
rect 307938 125536 307944 125548
rect 307996 125536 308002 125588
rect 346210 125576 346216 125588
rect 346171 125548 346216 125576
rect 346210 125536 346216 125548
rect 346268 125536 346274 125588
rect 357250 125576 357256 125588
rect 357211 125548 357256 125576
rect 357250 125536 357256 125548
rect 357308 125536 357314 125588
rect 211264 125508 211292 125536
rect 211338 125508 211344 125520
rect 211264 125480 211344 125508
rect 211338 125468 211344 125480
rect 211396 125468 211402 125520
rect 234798 124284 234804 124296
rect 234759 124256 234804 124284
rect 234798 124244 234804 124256
rect 234856 124244 234862 124296
rect 424686 124284 424692 124296
rect 424647 124256 424692 124284
rect 424686 124244 424692 124256
rect 424744 124244 424750 124296
rect 153378 124216 153384 124228
rect 153339 124188 153384 124216
rect 153378 124176 153384 124188
rect 153436 124176 153442 124228
rect 156138 124216 156144 124228
rect 156099 124188 156144 124216
rect 156138 124176 156144 124188
rect 156196 124176 156202 124228
rect 168834 124216 168840 124228
rect 168795 124188 168840 124216
rect 168834 124176 168840 124188
rect 168892 124176 168898 124228
rect 245746 124216 245752 124228
rect 245707 124188 245752 124216
rect 245746 124176 245752 124188
rect 245804 124176 245810 124228
rect 162946 124148 162952 124160
rect 162907 124120 162952 124148
rect 162946 124108 162952 124120
rect 163004 124108 163010 124160
rect 189258 124148 189264 124160
rect 189219 124120 189264 124148
rect 189258 124108 189264 124120
rect 189316 124108 189322 124160
rect 190638 124108 190644 124160
rect 190696 124108 190702 124160
rect 192018 124148 192024 124160
rect 191979 124120 192024 124148
rect 192018 124108 192024 124120
rect 192076 124108 192082 124160
rect 234798 124148 234804 124160
rect 234759 124120 234804 124148
rect 234798 124108 234804 124120
rect 234856 124108 234862 124160
rect 238573 124151 238631 124157
rect 238573 124117 238585 124151
rect 238619 124148 238631 124151
rect 238662 124148 238668 124160
rect 238619 124120 238668 124148
rect 238619 124117 238631 124120
rect 238573 124111 238631 124117
rect 238662 124108 238668 124120
rect 238720 124108 238726 124160
rect 248322 124148 248328 124160
rect 248283 124120 248328 124148
rect 248322 124108 248328 124120
rect 248380 124108 248386 124160
rect 374270 124148 374276 124160
rect 374231 124120 374276 124148
rect 374270 124108 374276 124120
rect 374328 124108 374334 124160
rect 384390 124108 384396 124160
rect 384448 124108 384454 124160
rect 384482 124108 384488 124160
rect 384540 124108 384546 124160
rect 424686 124148 424692 124160
rect 424647 124120 424692 124148
rect 424686 124108 424692 124120
rect 424744 124108 424750 124160
rect 190656 124080 190684 124108
rect 190914 124080 190920 124092
rect 190656 124052 190920 124080
rect 190914 124040 190920 124052
rect 190972 124040 190978 124092
rect 384408 123956 384436 124108
rect 384500 124024 384528 124108
rect 384482 123972 384488 124024
rect 384540 123972 384546 124024
rect 384390 123904 384396 123956
rect 384448 123904 384454 123956
rect 151998 122816 152004 122868
rect 152056 122856 152062 122868
rect 152090 122856 152096 122868
rect 152056 122828 152096 122856
rect 152056 122816 152062 122828
rect 152090 122816 152096 122828
rect 152148 122816 152154 122868
rect 196158 122816 196164 122868
rect 196216 122856 196222 122868
rect 196250 122856 196256 122868
rect 196216 122828 196256 122856
rect 196216 122816 196222 122828
rect 196250 122816 196256 122828
rect 196308 122816 196314 122868
rect 379146 122856 379152 122868
rect 379107 122828 379152 122856
rect 379146 122816 379152 122828
rect 379204 122816 379210 122868
rect 263778 122788 263784 122800
rect 263739 122760 263784 122788
rect 263778 122748 263784 122760
rect 263836 122748 263842 122800
rect 264974 122788 264980 122800
rect 264935 122760 264980 122788
rect 264974 122748 264980 122760
rect 265032 122748 265038 122800
rect 423214 122788 423220 122800
rect 423175 122760 423220 122788
rect 423214 122748 423220 122760
rect 423272 122748 423278 122800
rect 151998 121428 152004 121440
rect 151959 121400 152004 121428
rect 151998 121388 152004 121400
rect 152056 121388 152062 121440
rect 208578 120504 208584 120556
rect 208636 120544 208642 120556
rect 208670 120544 208676 120556
rect 208636 120516 208676 120544
rect 208636 120504 208642 120516
rect 208670 120504 208676 120516
rect 208728 120504 208734 120556
rect 156138 118736 156144 118788
rect 156196 118736 156202 118788
rect 222562 118736 222568 118788
rect 222620 118736 222626 118788
rect 223850 118736 223856 118788
rect 223908 118736 223914 118788
rect 156156 118652 156184 118736
rect 222580 118652 222608 118736
rect 223868 118652 223896 118736
rect 247218 118668 247224 118720
rect 247276 118668 247282 118720
rect 403434 118668 403440 118720
rect 403492 118668 403498 118720
rect 156138 118600 156144 118652
rect 156196 118600 156202 118652
rect 173986 118640 173992 118652
rect 173947 118612 173992 118640
rect 173986 118600 173992 118612
rect 174044 118600 174050 118652
rect 222562 118600 222568 118652
rect 222620 118600 222626 118652
rect 223850 118600 223856 118652
rect 223908 118600 223914 118652
rect 247236 118640 247264 118668
rect 247310 118640 247316 118652
rect 247236 118612 247316 118640
rect 247310 118600 247316 118612
rect 247368 118600 247374 118652
rect 252738 118640 252744 118652
rect 252699 118612 252744 118640
rect 252738 118600 252744 118612
rect 252796 118600 252802 118652
rect 284386 118640 284392 118652
rect 284347 118612 284392 118640
rect 284386 118600 284392 118612
rect 284444 118600 284450 118652
rect 307938 118640 307944 118652
rect 307899 118612 307944 118640
rect 307938 118600 307944 118612
rect 307996 118600 308002 118652
rect 346210 118640 346216 118652
rect 346171 118612 346216 118640
rect 346210 118600 346216 118612
rect 346268 118600 346274 118652
rect 357250 118640 357256 118652
rect 357211 118612 357256 118640
rect 357250 118600 357256 118612
rect 357308 118600 357314 118652
rect 403452 118640 403480 118668
rect 403526 118640 403532 118652
rect 403452 118612 403532 118640
rect 403526 118600 403532 118612
rect 403584 118600 403590 118652
rect 150710 116328 150716 116340
rect 150671 116300 150716 116328
rect 150710 116288 150716 116300
rect 150768 116288 150774 116340
rect 178218 115988 178224 116000
rect 178179 115960 178224 115988
rect 178218 115948 178224 115960
rect 178276 115948 178282 116000
rect 236270 115880 236276 115932
rect 236328 115880 236334 115932
rect 237558 115880 237564 115932
rect 237616 115880 237622 115932
rect 403250 115880 403256 115932
rect 403308 115920 403314 115932
rect 403526 115920 403532 115932
rect 403308 115892 403532 115920
rect 403308 115880 403314 115892
rect 403526 115880 403532 115892
rect 403584 115880 403590 115932
rect 168834 115852 168840 115864
rect 168760 115824 168840 115852
rect 168760 115796 168788 115824
rect 168834 115812 168840 115824
rect 168892 115812 168898 115864
rect 236288 115852 236316 115880
rect 236362 115852 236368 115864
rect 236288 115824 236368 115852
rect 236362 115812 236368 115824
rect 236420 115812 236426 115864
rect 237576 115852 237604 115880
rect 237650 115852 237656 115864
rect 237576 115824 237656 115852
rect 237650 115812 237656 115824
rect 237708 115812 237714 115864
rect 168742 115744 168748 115796
rect 168800 115744 168806 115796
rect 153470 114588 153476 114640
rect 153528 114588 153534 114640
rect 216950 114628 216956 114640
rect 216876 114600 216956 114628
rect 153286 114520 153292 114572
rect 153344 114560 153350 114572
rect 153488 114560 153516 114588
rect 216876 114572 216904 114600
rect 216950 114588 216956 114600
rect 217008 114588 217014 114640
rect 153344 114532 153516 114560
rect 162949 114563 163007 114569
rect 153344 114520 153350 114532
rect 162949 114529 162961 114563
rect 162995 114560 163007 114563
rect 163038 114560 163044 114572
rect 162995 114532 163044 114560
rect 162995 114529 163007 114532
rect 162949 114523 163007 114529
rect 163038 114520 163044 114532
rect 163096 114520 163102 114572
rect 189258 114560 189264 114572
rect 189219 114532 189264 114560
rect 189258 114520 189264 114532
rect 189316 114520 189322 114572
rect 216858 114520 216864 114572
rect 216916 114520 216922 114572
rect 234798 114560 234804 114572
rect 234759 114532 234804 114560
rect 234798 114520 234804 114532
rect 234856 114520 234862 114572
rect 238570 114560 238576 114572
rect 238531 114532 238576 114560
rect 238570 114520 238576 114532
rect 238628 114520 238634 114572
rect 248322 114560 248328 114572
rect 248283 114532 248328 114560
rect 248322 114520 248328 114532
rect 248380 114520 248386 114572
rect 374270 114560 374276 114572
rect 374231 114532 374276 114560
rect 374270 114520 374276 114532
rect 374328 114520 374334 114572
rect 384574 114520 384580 114572
rect 384632 114560 384638 114572
rect 384666 114560 384672 114572
rect 384632 114532 384672 114560
rect 384632 114520 384638 114532
rect 384666 114520 384672 114532
rect 384724 114520 384730 114572
rect 424689 114563 424747 114569
rect 424689 114529 424701 114563
rect 424735 114560 424747 114563
rect 424778 114560 424784 114572
rect 424735 114532 424784 114560
rect 424735 114529 424747 114532
rect 424689 114523 424747 114529
rect 424778 114520 424784 114532
rect 424836 114520 424842 114572
rect 168834 114492 168840 114504
rect 168795 114464 168840 114492
rect 168834 114452 168840 114464
rect 168892 114452 168898 114504
rect 207014 114492 207020 114504
rect 206975 114464 207020 114492
rect 207014 114452 207020 114464
rect 207072 114452 207078 114504
rect 271966 114452 271972 114504
rect 272024 114492 272030 114504
rect 272058 114492 272064 114504
rect 272024 114464 272064 114492
rect 272024 114452 272030 114464
rect 272058 114452 272064 114464
rect 272116 114452 272122 114504
rect 153286 114424 153292 114436
rect 153247 114396 153292 114424
rect 153286 114384 153292 114396
rect 153344 114384 153350 114436
rect 384574 114424 384580 114436
rect 384535 114396 384580 114424
rect 384574 114384 384580 114396
rect 384632 114384 384638 114436
rect 263778 114288 263784 114300
rect 263739 114260 263784 114288
rect 263778 114248 263784 114260
rect 263836 114248 263842 114300
rect 191929 113271 191987 113277
rect 191929 113237 191941 113271
rect 191975 113268 191987 113271
rect 192018 113268 192024 113280
rect 191975 113240 192024 113268
rect 191975 113237 191987 113240
rect 191929 113231 191987 113237
rect 192018 113228 192024 113240
rect 192076 113228 192082 113280
rect 194686 113160 194692 113212
rect 194744 113200 194750 113212
rect 194778 113200 194784 113212
rect 194744 113172 194784 113200
rect 194744 113160 194750 113172
rect 194778 113160 194784 113172
rect 194836 113160 194842 113212
rect 196158 113160 196164 113212
rect 196216 113200 196222 113212
rect 196250 113200 196256 113212
rect 196216 113172 196256 113200
rect 196216 113160 196222 113172
rect 196250 113160 196256 113172
rect 196308 113160 196314 113212
rect 264977 113203 265035 113209
rect 264977 113169 264989 113203
rect 265023 113200 265035 113203
rect 265066 113200 265072 113212
rect 265023 113172 265072 113200
rect 265023 113169 265035 113172
rect 264977 113163 265035 113169
rect 265066 113160 265072 113172
rect 265124 113160 265130 113212
rect 423217 113203 423275 113209
rect 423217 113169 423229 113203
rect 423263 113200 423275 113203
rect 423306 113200 423312 113212
rect 423263 113172 423312 113200
rect 423263 113169 423275 113172
rect 423217 113163 423275 113169
rect 423306 113160 423312 113172
rect 423364 113160 423370 113212
rect 151998 111840 152004 111852
rect 151959 111812 152004 111840
rect 151998 111800 152004 111812
rect 152056 111800 152062 111852
rect 191926 111840 191932 111852
rect 191887 111812 191932 111840
rect 191926 111800 191932 111812
rect 191984 111800 191990 111852
rect 577774 111732 577780 111784
rect 577832 111772 577838 111784
rect 580626 111772 580632 111784
rect 577832 111744 580632 111772
rect 577832 111732 577838 111744
rect 580626 111732 580632 111744
rect 580684 111732 580690 111784
rect 245749 109735 245807 109741
rect 245749 109701 245761 109735
rect 245795 109732 245807 109735
rect 245930 109732 245936 109744
rect 245795 109704 245936 109732
rect 245795 109701 245807 109704
rect 245749 109695 245807 109701
rect 245930 109692 245936 109704
rect 245988 109692 245994 109744
rect 423033 109735 423091 109741
rect 423033 109701 423045 109735
rect 423079 109732 423091 109735
rect 423306 109732 423312 109744
rect 423079 109704 423312 109732
rect 423079 109701 423091 109704
rect 423033 109695 423091 109701
rect 423306 109692 423312 109704
rect 423364 109692 423370 109744
rect 218330 109080 218336 109132
rect 218388 109080 218394 109132
rect 219618 109080 219624 109132
rect 219676 109080 219682 109132
rect 162854 109012 162860 109064
rect 162912 109052 162918 109064
rect 163038 109052 163044 109064
rect 162912 109024 163044 109052
rect 162912 109012 162918 109024
rect 163038 109012 163044 109024
rect 163096 109012 163102 109064
rect 173894 109012 173900 109064
rect 173952 109052 173958 109064
rect 174078 109052 174084 109064
rect 173952 109024 174084 109052
rect 173952 109012 173958 109024
rect 174078 109012 174084 109024
rect 174136 109012 174142 109064
rect 218348 108996 218376 109080
rect 219636 108996 219664 109080
rect 252646 109012 252652 109064
rect 252704 109052 252710 109064
rect 252830 109052 252836 109064
rect 252704 109024 252836 109052
rect 252704 109012 252710 109024
rect 252830 109012 252836 109024
rect 252888 109012 252894 109064
rect 284294 109012 284300 109064
rect 284352 109052 284358 109064
rect 284478 109052 284484 109064
rect 284352 109024 284484 109052
rect 284352 109012 284358 109024
rect 284478 109012 284484 109024
rect 284536 109012 284542 109064
rect 307846 109012 307852 109064
rect 307904 109052 307910 109064
rect 308030 109052 308036 109064
rect 307904 109024 308036 109052
rect 307904 109012 307910 109024
rect 308030 109012 308036 109024
rect 308088 109012 308094 109064
rect 346118 109012 346124 109064
rect 346176 109052 346182 109064
rect 346302 109052 346308 109064
rect 346176 109024 346308 109052
rect 346176 109012 346182 109024
rect 346302 109012 346308 109024
rect 346360 109012 346366 109064
rect 357158 109012 357164 109064
rect 357216 109052 357222 109064
rect 357342 109052 357348 109064
rect 357216 109024 357348 109052
rect 357216 109012 357222 109024
rect 357342 109012 357348 109024
rect 357400 109012 357406 109064
rect 218330 108944 218336 108996
rect 218388 108944 218394 108996
rect 219618 108944 219624 108996
rect 219676 108944 219682 108996
rect 424689 107083 424747 107089
rect 424689 107049 424701 107083
rect 424735 107080 424747 107083
rect 424778 107080 424784 107092
rect 424735 107052 424784 107080
rect 424735 107049 424747 107052
rect 424689 107043 424747 107049
rect 424778 107040 424784 107052
rect 424836 107040 424842 107092
rect 208397 106335 208455 106341
rect 208397 106301 208409 106335
rect 208443 106332 208455 106335
rect 208578 106332 208584 106344
rect 208443 106304 208584 106332
rect 208443 106301 208455 106304
rect 208397 106295 208455 106301
rect 208578 106292 208584 106304
rect 208636 106292 208642 106344
rect 211338 106292 211344 106344
rect 211396 106292 211402 106344
rect 238570 106292 238576 106344
rect 238628 106332 238634 106344
rect 238662 106332 238668 106344
rect 238628 106304 238668 106332
rect 238628 106292 238634 106304
rect 238662 106292 238668 106304
rect 238720 106292 238726 106344
rect 168834 106264 168840 106276
rect 168795 106236 168840 106264
rect 168834 106224 168840 106236
rect 168892 106224 168898 106276
rect 173986 106264 173992 106276
rect 173947 106236 173992 106264
rect 173986 106224 173992 106236
rect 174044 106224 174050 106276
rect 178218 106264 178224 106276
rect 178179 106236 178224 106264
rect 178218 106224 178224 106236
rect 178276 106224 178282 106276
rect 190638 106264 190644 106276
rect 190599 106236 190644 106264
rect 190638 106224 190644 106236
rect 190696 106224 190702 106276
rect 154758 106196 154764 106208
rect 154719 106168 154764 106196
rect 154758 106156 154764 106168
rect 154816 106156 154822 106208
rect 211356 106140 211384 106292
rect 222470 106224 222476 106276
rect 222528 106264 222534 106276
rect 222562 106264 222568 106276
rect 222528 106236 222568 106264
rect 222528 106224 222534 106236
rect 222562 106224 222568 106236
rect 222620 106224 222626 106276
rect 223758 106224 223764 106276
rect 223816 106264 223822 106276
rect 223850 106264 223856 106276
rect 223816 106236 223856 106264
rect 223816 106224 223822 106236
rect 223850 106224 223856 106236
rect 223908 106224 223914 106276
rect 252738 106264 252744 106276
rect 252699 106236 252744 106264
rect 252738 106224 252744 106236
rect 252796 106224 252802 106276
rect 284386 106264 284392 106276
rect 284347 106236 284392 106264
rect 284386 106224 284392 106236
rect 284444 106224 284450 106276
rect 307938 106264 307944 106276
rect 307899 106236 307944 106264
rect 307938 106224 307944 106236
rect 307996 106224 308002 106276
rect 346210 106264 346216 106276
rect 346171 106236 346216 106264
rect 346210 106224 346216 106236
rect 346268 106224 346274 106276
rect 357250 106264 357256 106276
rect 357211 106236 357256 106264
rect 357250 106224 357256 106236
rect 357308 106224 357314 106276
rect 211338 106088 211344 106140
rect 211396 106088 211402 106140
rect 153289 104907 153347 104913
rect 153289 104873 153301 104907
rect 153335 104904 153347 104907
rect 153378 104904 153384 104916
rect 153335 104876 153384 104904
rect 153335 104873 153347 104876
rect 153289 104867 153347 104873
rect 153378 104864 153384 104876
rect 153436 104864 153442 104916
rect 189166 104864 189172 104916
rect 189224 104904 189230 104916
rect 189258 104904 189264 104916
rect 189224 104876 189264 104904
rect 189224 104864 189230 104876
rect 189258 104864 189264 104876
rect 189316 104864 189322 104916
rect 205818 104864 205824 104916
rect 205876 104904 205882 104916
rect 206002 104904 206008 104916
rect 205876 104876 206008 104904
rect 205876 104864 205882 104876
rect 206002 104864 206008 104876
rect 206060 104864 206066 104916
rect 207017 104907 207075 104913
rect 207017 104873 207029 104907
rect 207063 104904 207075 104907
rect 207106 104904 207112 104916
rect 207063 104876 207112 104904
rect 207063 104873 207075 104876
rect 207017 104867 207075 104873
rect 207106 104864 207112 104876
rect 207164 104864 207170 104916
rect 208394 104904 208400 104916
rect 208355 104876 208400 104904
rect 208394 104864 208400 104876
rect 208452 104864 208458 104916
rect 245746 104904 245752 104916
rect 245707 104876 245752 104904
rect 245746 104864 245752 104876
rect 245804 104864 245810 104916
rect 384577 104907 384635 104913
rect 384577 104873 384589 104907
rect 384623 104904 384635 104907
rect 384850 104904 384856 104916
rect 384623 104876 384856 104904
rect 384623 104873 384635 104876
rect 384577 104867 384635 104873
rect 384850 104864 384856 104876
rect 384908 104864 384914 104916
rect 423030 104904 423036 104916
rect 422991 104876 423036 104904
rect 423030 104864 423036 104876
rect 423088 104864 423094 104916
rect 168834 104836 168840 104848
rect 168795 104808 168840 104836
rect 168834 104796 168840 104808
rect 168892 104796 168898 104848
rect 222470 104796 222476 104848
rect 222528 104796 222534 104848
rect 223758 104836 223764 104848
rect 223719 104808 223764 104836
rect 223758 104796 223764 104808
rect 223816 104796 223822 104848
rect 238662 104836 238668 104848
rect 238623 104808 238668 104836
rect 238662 104796 238668 104808
rect 238720 104796 238726 104848
rect 248322 104836 248328 104848
rect 248283 104808 248328 104836
rect 248322 104796 248328 104808
rect 248380 104796 248386 104848
rect 263778 104836 263784 104848
rect 263739 104808 263784 104836
rect 263778 104796 263784 104808
rect 263836 104796 263842 104848
rect 374270 104836 374276 104848
rect 374231 104808 374276 104836
rect 374270 104796 374276 104808
rect 374328 104796 374334 104848
rect 222488 104768 222516 104796
rect 222562 104768 222568 104780
rect 222488 104740 222568 104768
rect 222562 104728 222568 104740
rect 222620 104728 222626 104780
rect 150713 103547 150771 103553
rect 150713 103513 150725 103547
rect 150759 103544 150771 103547
rect 150802 103544 150808 103556
rect 150759 103516 150808 103544
rect 150759 103513 150771 103516
rect 150713 103507 150771 103513
rect 150802 103504 150808 103516
rect 150860 103504 150866 103556
rect 206002 103476 206008 103488
rect 205963 103448 206008 103476
rect 206002 103436 206008 103448
rect 206060 103436 206066 103488
rect 208394 103476 208400 103488
rect 208355 103448 208400 103476
rect 208394 103436 208400 103448
rect 208452 103436 208458 103488
rect 270494 103476 270500 103488
rect 270455 103448 270500 103476
rect 270494 103436 270500 103448
rect 270552 103436 270558 103488
rect 272058 103476 272064 103488
rect 272019 103448 272064 103476
rect 272058 103436 272064 103448
rect 272116 103436 272122 103488
rect 191742 102144 191748 102196
rect 191800 102184 191806 102196
rect 192202 102184 192208 102196
rect 191800 102156 192208 102184
rect 191800 102144 191806 102156
rect 192202 102144 192208 102156
rect 192260 102144 192266 102196
rect 151998 102116 152004 102128
rect 151959 102088 152004 102116
rect 151998 102076 152004 102088
rect 152056 102076 152062 102128
rect 190638 101368 190644 101380
rect 190599 101340 190644 101368
rect 190638 101328 190644 101340
rect 190696 101328 190702 101380
rect 379146 100076 379152 100088
rect 379107 100048 379152 100076
rect 379146 100036 379152 100048
rect 379204 100036 379210 100088
rect 153378 99424 153384 99476
rect 153436 99424 153442 99476
rect 156138 99424 156144 99476
rect 156196 99424 156202 99476
rect 214098 99424 214104 99476
rect 214156 99424 214162 99476
rect 153396 99340 153424 99424
rect 156156 99340 156184 99424
rect 162946 99356 162952 99408
rect 163004 99356 163010 99408
rect 153378 99288 153384 99340
rect 153436 99288 153442 99340
rect 156138 99288 156144 99340
rect 156196 99288 156202 99340
rect 162964 99328 162992 99356
rect 214116 99340 214144 99424
rect 247218 99356 247224 99408
rect 247276 99356 247282 99408
rect 403434 99356 403440 99408
rect 403492 99356 403498 99408
rect 163038 99328 163044 99340
rect 162964 99300 163044 99328
rect 163038 99288 163044 99300
rect 163096 99288 163102 99340
rect 173986 99328 173992 99340
rect 173947 99300 173992 99328
rect 173986 99288 173992 99300
rect 174044 99288 174050 99340
rect 214098 99288 214104 99340
rect 214156 99288 214162 99340
rect 247236 99328 247264 99356
rect 247310 99328 247316 99340
rect 247236 99300 247316 99328
rect 247310 99288 247316 99300
rect 247368 99288 247374 99340
rect 252738 99328 252744 99340
rect 252699 99300 252744 99328
rect 252738 99288 252744 99300
rect 252796 99288 252802 99340
rect 284386 99328 284392 99340
rect 284347 99300 284392 99328
rect 284386 99288 284392 99300
rect 284444 99288 284450 99340
rect 307938 99328 307944 99340
rect 307899 99300 307944 99328
rect 307938 99288 307944 99300
rect 307996 99288 308002 99340
rect 346210 99328 346216 99340
rect 346171 99300 346216 99328
rect 346210 99288 346216 99300
rect 346268 99288 346274 99340
rect 357250 99328 357256 99340
rect 357211 99300 357256 99328
rect 357250 99288 357256 99300
rect 357308 99288 357314 99340
rect 403452 99328 403480 99356
rect 403526 99328 403532 99340
rect 403452 99300 403532 99328
rect 403526 99288 403532 99300
rect 403584 99288 403590 99340
rect 424686 99328 424692 99340
rect 424647 99300 424692 99328
rect 424686 99288 424692 99300
rect 424744 99288 424750 99340
rect 198274 98676 198280 98728
rect 198332 98676 198338 98728
rect 198292 98592 198320 98676
rect 198274 98540 198280 98592
rect 198332 98540 198338 98592
rect 263778 96880 263784 96892
rect 263739 96852 263784 96880
rect 263778 96840 263784 96852
rect 263836 96840 263842 96892
rect 154758 96744 154764 96756
rect 154719 96716 154764 96744
rect 154758 96704 154764 96716
rect 154816 96704 154822 96756
rect 178218 96676 178224 96688
rect 178179 96648 178224 96676
rect 178218 96636 178224 96648
rect 178276 96636 178282 96688
rect 154758 96568 154764 96620
rect 154816 96608 154822 96620
rect 154942 96608 154948 96620
rect 154816 96580 154948 96608
rect 154816 96568 154822 96580
rect 154942 96568 154948 96580
rect 155000 96568 155006 96620
rect 162854 96568 162860 96620
rect 162912 96608 162918 96620
rect 163038 96608 163044 96620
rect 162912 96580 163044 96608
rect 162912 96568 162918 96580
rect 163038 96568 163044 96580
rect 163096 96568 163102 96620
rect 303614 96568 303620 96620
rect 303672 96608 303678 96620
rect 303706 96608 303712 96620
rect 303672 96580 303712 96608
rect 303672 96568 303678 96580
rect 303706 96568 303712 96580
rect 303764 96568 303770 96620
rect 384666 96568 384672 96620
rect 384724 96608 384730 96620
rect 384850 96608 384856 96620
rect 384724 96580 384856 96608
rect 384724 96568 384730 96580
rect 384850 96568 384856 96580
rect 384908 96568 384914 96620
rect 403250 96568 403256 96620
rect 403308 96608 403314 96620
rect 403526 96608 403532 96620
rect 403308 96580 403532 96608
rect 403308 96568 403314 96580
rect 403526 96568 403532 96580
rect 403584 96568 403590 96620
rect 423030 96568 423036 96620
rect 423088 96608 423094 96620
rect 423122 96608 423128 96620
rect 423088 96580 423128 96608
rect 423088 96568 423094 96580
rect 423122 96568 423128 96580
rect 423180 96568 423186 96620
rect 168834 95248 168840 95260
rect 168795 95220 168840 95248
rect 168834 95208 168840 95220
rect 168892 95208 168898 95260
rect 207106 95208 207112 95260
rect 207164 95208 207170 95260
rect 223761 95251 223819 95257
rect 223761 95217 223773 95251
rect 223807 95248 223819 95251
rect 224034 95248 224040 95260
rect 223807 95220 224040 95248
rect 223807 95217 223819 95220
rect 223761 95211 223819 95217
rect 224034 95208 224040 95220
rect 224092 95208 224098 95260
rect 238662 95248 238668 95260
rect 238623 95220 238668 95248
rect 238662 95208 238668 95220
rect 238720 95208 238726 95260
rect 248322 95248 248328 95260
rect 248283 95220 248328 95248
rect 248322 95208 248328 95220
rect 248380 95208 248386 95260
rect 374270 95248 374276 95260
rect 374231 95220 374276 95248
rect 374270 95208 374276 95220
rect 374328 95208 374334 95260
rect 188982 95180 188988 95192
rect 188943 95152 188988 95180
rect 188982 95140 188988 95152
rect 189040 95140 189046 95192
rect 207124 95112 207152 95208
rect 211338 95180 211344 95192
rect 211299 95152 211344 95180
rect 211338 95140 211344 95152
rect 211396 95140 211402 95192
rect 216858 95180 216864 95192
rect 216819 95152 216864 95180
rect 216858 95140 216864 95152
rect 216916 95140 216922 95192
rect 218330 95180 218336 95192
rect 218291 95152 218336 95180
rect 218330 95140 218336 95152
rect 218388 95140 218394 95192
rect 219618 95180 219624 95192
rect 219579 95152 219624 95180
rect 219618 95140 219624 95152
rect 219676 95140 219682 95192
rect 207198 95112 207204 95124
rect 207124 95084 207204 95112
rect 207198 95072 207204 95084
rect 207256 95072 207262 95124
rect 208397 95115 208455 95121
rect 208397 95081 208409 95115
rect 208443 95112 208455 95115
rect 208762 95112 208768 95124
rect 208443 95084 208768 95112
rect 208443 95081 208455 95084
rect 208397 95075 208455 95081
rect 208762 95072 208768 95084
rect 208820 95072 208826 95124
rect 206002 93888 206008 93900
rect 205963 93860 206008 93888
rect 206002 93848 206008 93860
rect 206060 93848 206066 93900
rect 270497 93891 270555 93897
rect 270497 93857 270509 93891
rect 270543 93888 270555 93891
rect 270586 93888 270592 93900
rect 270543 93860 270592 93888
rect 270543 93857 270555 93860
rect 270497 93851 270555 93857
rect 270586 93848 270592 93860
rect 270644 93848 270650 93900
rect 272058 93888 272064 93900
rect 272019 93860 272064 93888
rect 272058 93848 272064 93860
rect 272116 93848 272122 93900
rect 226610 93820 226616 93832
rect 226571 93792 226616 93820
rect 226610 93780 226616 93792
rect 226668 93780 226674 93832
rect 151998 92528 152004 92540
rect 151959 92500 152004 92528
rect 151998 92488 152004 92500
rect 152056 92488 152062 92540
rect 192018 92488 192024 92540
rect 192076 92528 192082 92540
rect 192110 92528 192116 92540
rect 192076 92500 192116 92528
rect 192076 92488 192082 92500
rect 192110 92488 192116 92500
rect 192168 92488 192174 92540
rect 226610 92528 226616 92540
rect 226571 92500 226616 92528
rect 226610 92488 226616 92500
rect 226668 92488 226674 92540
rect 150710 92420 150716 92472
rect 150768 92460 150774 92472
rect 150986 92460 150992 92472
rect 150768 92432 150992 92460
rect 150768 92420 150774 92432
rect 150986 92420 150992 92432
rect 151044 92420 151050 92472
rect 168466 91740 168472 91792
rect 168524 91780 168530 91792
rect 168834 91780 168840 91792
rect 168524 91752 168840 91780
rect 168524 91740 168530 91752
rect 168834 91740 168840 91752
rect 168892 91740 168898 91792
rect 190638 91740 190644 91792
rect 190696 91780 190702 91792
rect 190822 91780 190828 91792
rect 190696 91752 190828 91780
rect 190696 91740 190702 91752
rect 190822 91740 190828 91752
rect 190880 91740 190886 91792
rect 245749 90423 245807 90429
rect 245749 90389 245761 90423
rect 245795 90420 245807 90423
rect 245930 90420 245936 90432
rect 245795 90392 245936 90420
rect 245795 90389 245807 90392
rect 245749 90383 245807 90389
rect 245930 90380 245936 90392
rect 245988 90380 245994 90432
rect 173894 89700 173900 89752
rect 173952 89740 173958 89752
rect 174078 89740 174084 89752
rect 173952 89712 174084 89740
rect 173952 89700 173958 89712
rect 174078 89700 174084 89712
rect 174136 89700 174142 89752
rect 252646 89700 252652 89752
rect 252704 89740 252710 89752
rect 252830 89740 252836 89752
rect 252704 89712 252836 89740
rect 252704 89700 252710 89712
rect 252830 89700 252836 89712
rect 252888 89700 252894 89752
rect 264974 89700 264980 89752
rect 265032 89700 265038 89752
rect 284294 89700 284300 89752
rect 284352 89740 284358 89752
rect 284478 89740 284484 89752
rect 284352 89712 284484 89740
rect 284352 89700 284358 89712
rect 284478 89700 284484 89712
rect 284536 89700 284542 89752
rect 307846 89700 307852 89752
rect 307904 89740 307910 89752
rect 308030 89740 308036 89752
rect 307904 89712 308036 89740
rect 307904 89700 307910 89712
rect 308030 89700 308036 89712
rect 308088 89700 308094 89752
rect 346118 89700 346124 89752
rect 346176 89740 346182 89752
rect 346302 89740 346308 89752
rect 346176 89712 346308 89740
rect 346176 89700 346182 89712
rect 346302 89700 346308 89712
rect 346360 89700 346366 89752
rect 357158 89700 357164 89752
rect 357216 89740 357222 89752
rect 357342 89740 357348 89752
rect 357216 89712 357348 89740
rect 357216 89700 357222 89712
rect 357342 89700 357348 89712
rect 357400 89700 357406 89752
rect 264992 89672 265020 89700
rect 265066 89672 265072 89684
rect 264992 89644 265072 89672
rect 265066 89632 265072 89644
rect 265124 89632 265130 89684
rect 379146 89400 379152 89412
rect 379107 89372 379152 89400
rect 379146 89360 379152 89372
rect 379204 89360 379210 89412
rect 189074 86980 189080 87032
rect 189132 86980 189138 87032
rect 206002 87020 206008 87032
rect 205963 86992 206008 87020
rect 206002 86980 206008 86992
rect 206060 86980 206066 87032
rect 229186 86980 229192 87032
rect 229244 87020 229250 87032
rect 229278 87020 229284 87032
rect 229244 86992 229284 87020
rect 229244 86980 229250 86992
rect 229278 86980 229284 86992
rect 229336 86980 229342 87032
rect 236178 86980 236184 87032
rect 236236 87020 236242 87032
rect 236270 87020 236276 87032
rect 236236 86992 236276 87020
rect 236236 86980 236242 86992
rect 236270 86980 236276 86992
rect 236328 86980 236334 87032
rect 169757 86955 169815 86961
rect 169757 86921 169769 86955
rect 169803 86952 169815 86955
rect 169846 86952 169852 86964
rect 169803 86924 169852 86952
rect 169803 86921 169815 86924
rect 169757 86915 169815 86921
rect 169846 86912 169852 86924
rect 169904 86912 169910 86964
rect 173986 86952 173992 86964
rect 173947 86924 173992 86952
rect 173986 86912 173992 86924
rect 174044 86912 174050 86964
rect 178218 86952 178224 86964
rect 178179 86924 178224 86952
rect 178218 86912 178224 86924
rect 178276 86912 178282 86964
rect 189092 86896 189120 86980
rect 190638 86952 190644 86964
rect 190599 86924 190644 86952
rect 190638 86912 190644 86924
rect 190696 86912 190702 86964
rect 191926 86952 191932 86964
rect 191887 86924 191932 86952
rect 191926 86912 191932 86924
rect 191984 86912 191990 86964
rect 222470 86912 222476 86964
rect 222528 86952 222534 86964
rect 222562 86952 222568 86964
rect 222528 86924 222568 86952
rect 222528 86912 222534 86924
rect 222562 86912 222568 86924
rect 222620 86912 222626 86964
rect 223758 86912 223764 86964
rect 223816 86952 223822 86964
rect 223850 86952 223856 86964
rect 223816 86924 223856 86952
rect 223816 86912 223822 86924
rect 223850 86912 223856 86924
rect 223908 86912 223914 86964
rect 247037 86955 247095 86961
rect 247037 86921 247049 86955
rect 247083 86952 247095 86955
rect 247126 86952 247132 86964
rect 247083 86924 247132 86952
rect 247083 86921 247095 86924
rect 247037 86915 247095 86921
rect 247126 86912 247132 86924
rect 247184 86912 247190 86964
rect 252738 86952 252744 86964
rect 252699 86924 252744 86952
rect 252738 86912 252744 86924
rect 252796 86912 252802 86964
rect 258077 86955 258135 86961
rect 258077 86921 258089 86955
rect 258123 86952 258135 86955
rect 258166 86952 258172 86964
rect 258123 86924 258172 86952
rect 258123 86921 258135 86924
rect 258077 86915 258135 86921
rect 258166 86912 258172 86924
rect 258224 86912 258230 86964
rect 284386 86952 284392 86964
rect 284347 86924 284392 86952
rect 284386 86912 284392 86924
rect 284444 86912 284450 86964
rect 307938 86952 307944 86964
rect 307899 86924 307944 86952
rect 307938 86912 307944 86924
rect 307996 86912 308002 86964
rect 346210 86952 346216 86964
rect 346171 86924 346216 86952
rect 346210 86912 346216 86924
rect 346268 86912 346274 86964
rect 357250 86952 357256 86964
rect 357211 86924 357256 86952
rect 357250 86912 357256 86924
rect 357308 86912 357314 86964
rect 423214 86912 423220 86964
rect 423272 86952 423278 86964
rect 423398 86952 423404 86964
rect 423272 86924 423404 86952
rect 423272 86912 423278 86924
rect 423398 86912 423404 86924
rect 423456 86912 423462 86964
rect 424686 86952 424692 86964
rect 424647 86924 424692 86952
rect 424686 86912 424692 86924
rect 424744 86912 424750 86964
rect 189074 86844 189080 86896
rect 189132 86844 189138 86896
rect 188985 85595 189043 85601
rect 188985 85561 188997 85595
rect 189031 85592 189043 85595
rect 189166 85592 189172 85604
rect 189031 85564 189172 85592
rect 189031 85561 189043 85564
rect 188985 85555 189043 85561
rect 189166 85552 189172 85564
rect 189224 85552 189230 85604
rect 194686 85552 194692 85604
rect 194744 85592 194750 85604
rect 194778 85592 194784 85604
rect 194744 85564 194784 85592
rect 194744 85552 194750 85564
rect 194778 85552 194784 85564
rect 194836 85552 194842 85604
rect 206002 85592 206008 85604
rect 205963 85564 206008 85592
rect 206002 85552 206008 85564
rect 206060 85552 206066 85604
rect 207014 85552 207020 85604
rect 207072 85592 207078 85604
rect 207198 85592 207204 85604
rect 207072 85564 207204 85592
rect 207072 85552 207078 85564
rect 207198 85552 207204 85564
rect 207256 85552 207262 85604
rect 211338 85592 211344 85604
rect 211299 85564 211344 85592
rect 211338 85552 211344 85564
rect 211396 85552 211402 85604
rect 216858 85592 216864 85604
rect 216819 85564 216864 85592
rect 216858 85552 216864 85564
rect 216916 85552 216922 85604
rect 218330 85592 218336 85604
rect 218291 85564 218336 85592
rect 218330 85552 218336 85564
rect 218388 85552 218394 85604
rect 219618 85592 219624 85604
rect 219579 85564 219624 85592
rect 219618 85552 219624 85564
rect 219676 85552 219682 85604
rect 162946 85524 162952 85536
rect 162907 85496 162952 85524
rect 162946 85484 162952 85496
rect 163004 85484 163010 85536
rect 223758 85524 223764 85536
rect 223719 85496 223764 85524
rect 223758 85484 223764 85496
rect 223816 85484 223822 85536
rect 229186 85484 229192 85536
rect 229244 85484 229250 85536
rect 238662 85524 238668 85536
rect 238623 85496 238668 85524
rect 238662 85484 238668 85496
rect 238720 85484 238726 85536
rect 248322 85524 248328 85536
rect 248283 85496 248328 85524
rect 248322 85484 248328 85496
rect 248380 85484 248386 85536
rect 270494 85524 270500 85536
rect 270455 85496 270500 85524
rect 270494 85484 270500 85496
rect 270552 85484 270558 85536
rect 272058 85524 272064 85536
rect 272019 85496 272064 85524
rect 272058 85484 272064 85496
rect 272116 85484 272122 85536
rect 374270 85524 374276 85536
rect 374231 85496 374276 85524
rect 374270 85484 374276 85496
rect 374328 85484 374334 85536
rect 229204 85456 229232 85484
rect 229370 85456 229376 85468
rect 229204 85428 229376 85456
rect 229370 85416 229376 85428
rect 229428 85416 229434 85468
rect 194778 84124 194784 84176
rect 194836 84164 194842 84176
rect 194873 84167 194931 84173
rect 194873 84164 194885 84167
rect 194836 84136 194885 84164
rect 194836 84124 194842 84136
rect 194873 84133 194885 84136
rect 194919 84133 194931 84167
rect 207014 84164 207020 84176
rect 206975 84136 207020 84164
rect 194873 84127 194931 84133
rect 207014 84124 207020 84136
rect 207072 84124 207078 84176
rect 208489 84167 208547 84173
rect 208489 84133 208501 84167
rect 208535 84164 208547 84167
rect 208578 84164 208584 84176
rect 208535 84136 208584 84164
rect 208535 84133 208547 84136
rect 208489 84127 208547 84133
rect 208578 84124 208584 84136
rect 208636 84124 208642 84176
rect 245749 83215 245807 83221
rect 245749 83181 245761 83215
rect 245795 83212 245807 83215
rect 246206 83212 246212 83224
rect 245795 83184 246212 83212
rect 245795 83181 245807 83184
rect 245749 83175 245807 83181
rect 246206 83172 246212 83184
rect 246264 83172 246270 83224
rect 151998 82804 152004 82816
rect 151959 82776 152004 82804
rect 151998 82764 152004 82776
rect 152056 82764 152062 82816
rect 226521 82807 226579 82813
rect 226521 82773 226533 82807
rect 226567 82804 226579 82807
rect 226610 82804 226616 82816
rect 226567 82776 226616 82804
rect 226567 82773 226579 82776
rect 226521 82767 226579 82773
rect 226610 82764 226616 82776
rect 226668 82764 226674 82816
rect 190638 80696 190644 80708
rect 190599 80668 190644 80696
rect 190638 80656 190644 80668
rect 190696 80656 190702 80708
rect 403434 80044 403440 80096
rect 403492 80044 403498 80096
rect 403452 79948 403480 80044
rect 403526 79948 403532 79960
rect 403452 79920 403532 79948
rect 403526 79908 403532 79920
rect 403584 79908 403590 79960
rect 168466 77324 168472 77376
rect 168524 77364 168530 77376
rect 168650 77364 168656 77376
rect 168524 77336 168656 77364
rect 168524 77324 168530 77336
rect 168650 77324 168656 77336
rect 168708 77324 168714 77376
rect 169754 77296 169760 77308
rect 169715 77268 169760 77296
rect 169754 77256 169760 77268
rect 169812 77256 169818 77308
rect 173989 77299 174047 77305
rect 173989 77265 174001 77299
rect 174035 77296 174047 77299
rect 174078 77296 174084 77308
rect 174035 77268 174084 77296
rect 174035 77265 174047 77268
rect 173989 77259 174047 77265
rect 174078 77256 174084 77268
rect 174136 77256 174142 77308
rect 178218 77296 178224 77308
rect 178179 77268 178224 77296
rect 178218 77256 178224 77268
rect 178276 77256 178282 77308
rect 234706 77256 234712 77308
rect 234764 77296 234770 77308
rect 234798 77296 234804 77308
rect 234764 77268 234804 77296
rect 234764 77256 234770 77268
rect 234798 77256 234804 77268
rect 234856 77256 234862 77308
rect 236178 77256 236184 77308
rect 236236 77296 236242 77308
rect 236270 77296 236276 77308
rect 236236 77268 236276 77296
rect 236236 77256 236242 77268
rect 236270 77256 236276 77268
rect 236328 77256 236334 77308
rect 237466 77256 237472 77308
rect 237524 77296 237530 77308
rect 237558 77296 237564 77308
rect 237524 77268 237564 77296
rect 237524 77256 237530 77268
rect 237558 77256 237564 77268
rect 237616 77256 237622 77308
rect 247034 77296 247040 77308
rect 246995 77268 247040 77296
rect 247034 77256 247040 77268
rect 247092 77256 247098 77308
rect 252741 77299 252799 77305
rect 252741 77265 252753 77299
rect 252787 77296 252799 77299
rect 252830 77296 252836 77308
rect 252787 77268 252836 77296
rect 252787 77265 252799 77268
rect 252741 77259 252799 77265
rect 252830 77256 252836 77268
rect 252888 77256 252894 77308
rect 258074 77296 258080 77308
rect 258035 77268 258080 77296
rect 258074 77256 258080 77268
rect 258132 77256 258138 77308
rect 265066 77256 265072 77308
rect 265124 77256 265130 77308
rect 284389 77299 284447 77305
rect 284389 77265 284401 77299
rect 284435 77296 284447 77299
rect 284478 77296 284484 77308
rect 284435 77268 284484 77296
rect 284435 77265 284447 77268
rect 284389 77259 284447 77265
rect 284478 77256 284484 77268
rect 284536 77256 284542 77308
rect 307941 77299 307999 77305
rect 307941 77265 307953 77299
rect 307987 77296 307999 77299
rect 308030 77296 308036 77308
rect 307987 77268 308036 77296
rect 307987 77265 307999 77268
rect 307941 77259 307999 77265
rect 308030 77256 308036 77268
rect 308088 77256 308094 77308
rect 346213 77299 346271 77305
rect 346213 77265 346225 77299
rect 346259 77296 346271 77299
rect 346302 77296 346308 77308
rect 346259 77268 346308 77296
rect 346259 77265 346271 77268
rect 346213 77259 346271 77265
rect 346302 77256 346308 77268
rect 346360 77256 346366 77308
rect 357253 77299 357311 77305
rect 357253 77265 357265 77299
rect 357299 77296 357311 77299
rect 357342 77296 357348 77308
rect 357299 77268 357348 77296
rect 357299 77265 357311 77268
rect 357253 77259 357311 77265
rect 357342 77256 357348 77268
rect 357400 77256 357406 77308
rect 424689 77299 424747 77305
rect 424689 77265 424701 77299
rect 424735 77296 424747 77299
rect 424778 77296 424784 77308
rect 424735 77268 424784 77296
rect 424735 77265 424747 77268
rect 424689 77259 424747 77265
rect 424778 77256 424784 77268
rect 424836 77256 424842 77308
rect 154758 77228 154764 77240
rect 154719 77200 154764 77228
rect 154758 77188 154764 77200
rect 154816 77188 154822 77240
rect 265084 77172 265112 77256
rect 303890 77228 303896 77240
rect 303851 77200 303896 77228
rect 303890 77188 303896 77200
rect 303948 77188 303954 77240
rect 577682 77188 577688 77240
rect 577740 77228 577746 77240
rect 579614 77228 579620 77240
rect 577740 77200 579620 77228
rect 577740 77188 577746 77200
rect 579614 77188 579620 77200
rect 579672 77188 579678 77240
rect 265066 77120 265072 77172
rect 265124 77120 265130 77172
rect 357253 77163 357311 77169
rect 357253 77129 357265 77163
rect 357299 77160 357311 77163
rect 357342 77160 357348 77172
rect 357299 77132 357348 77160
rect 357299 77129 357311 77132
rect 357253 77123 357311 77129
rect 357342 77120 357348 77132
rect 357400 77120 357406 77172
rect 198274 76004 198280 76016
rect 198200 75976 198280 76004
rect 198200 75948 198228 75976
rect 198274 75964 198280 75976
rect 198332 75964 198338 76016
rect 162949 75939 163007 75945
rect 162949 75905 162961 75939
rect 162995 75936 163007 75939
rect 163222 75936 163228 75948
rect 162995 75908 163228 75936
rect 162995 75905 163007 75908
rect 162949 75899 163007 75905
rect 163222 75896 163228 75908
rect 163280 75896 163286 75948
rect 191929 75939 191987 75945
rect 191929 75905 191941 75939
rect 191975 75936 191987 75939
rect 192018 75936 192024 75948
rect 191975 75908 192024 75936
rect 191975 75905 191987 75908
rect 191929 75899 191987 75905
rect 192018 75896 192024 75908
rect 192076 75896 192082 75948
rect 198182 75896 198188 75948
rect 198240 75896 198246 75948
rect 238662 75936 238668 75948
rect 238623 75908 238668 75936
rect 238662 75896 238668 75908
rect 238720 75896 238726 75948
rect 248322 75936 248328 75948
rect 248283 75908 248328 75936
rect 248322 75896 248328 75908
rect 248380 75896 248386 75948
rect 270497 75939 270555 75945
rect 270497 75905 270509 75939
rect 270543 75936 270555 75939
rect 270586 75936 270592 75948
rect 270543 75908 270592 75936
rect 270543 75905 270555 75908
rect 270497 75899 270555 75905
rect 270586 75896 270592 75908
rect 270644 75896 270650 75948
rect 272058 75936 272064 75948
rect 272019 75908 272064 75936
rect 272058 75896 272064 75908
rect 272116 75896 272122 75948
rect 374270 75936 374276 75948
rect 374231 75908 374276 75936
rect 374270 75896 374276 75908
rect 374328 75896 374334 75948
rect 196250 75828 196256 75880
rect 196308 75868 196314 75880
rect 196342 75868 196348 75880
rect 196308 75840 196348 75868
rect 196308 75828 196314 75840
rect 196342 75828 196348 75840
rect 196400 75828 196406 75880
rect 384666 75868 384672 75880
rect 384627 75840 384672 75868
rect 384666 75828 384672 75840
rect 384724 75828 384730 75880
rect 194778 74536 194784 74588
rect 194836 74576 194842 74588
rect 194873 74579 194931 74585
rect 194873 74576 194885 74579
rect 194836 74548 194885 74576
rect 194836 74536 194842 74548
rect 194873 74545 194885 74548
rect 194919 74545 194931 74579
rect 223758 74576 223764 74588
rect 223719 74548 223764 74576
rect 194873 74539 194931 74545
rect 223758 74536 223764 74548
rect 223816 74536 223822 74588
rect 198182 74468 198188 74520
rect 198240 74508 198246 74520
rect 198274 74508 198280 74520
rect 198240 74480 198280 74508
rect 198240 74468 198246 74480
rect 198274 74468 198280 74480
rect 198332 74468 198338 74520
rect 211246 74508 211252 74520
rect 211207 74480 211252 74508
rect 211246 74468 211252 74480
rect 211304 74468 211310 74520
rect 246025 74511 246083 74517
rect 246025 74477 246037 74511
rect 246071 74508 246083 74511
rect 246206 74508 246212 74520
rect 246071 74480 246212 74508
rect 246071 74477 246083 74480
rect 246025 74471 246083 74477
rect 246206 74468 246212 74480
rect 246264 74468 246270 74520
rect 151998 73216 152004 73228
rect 151959 73188 152004 73216
rect 151998 73176 152004 73188
rect 152056 73176 152062 73228
rect 219618 70564 219624 70576
rect 219544 70536 219624 70564
rect 190638 70496 190644 70508
rect 190599 70468 190644 70496
rect 190638 70456 190644 70468
rect 190696 70456 190702 70508
rect 192018 70496 192024 70508
rect 191944 70468 192024 70496
rect 191944 70372 191972 70468
rect 192018 70456 192024 70468
rect 192076 70456 192082 70508
rect 194778 70496 194784 70508
rect 194704 70468 194784 70496
rect 194704 70372 194732 70468
rect 194778 70456 194784 70468
rect 194836 70456 194842 70508
rect 216858 70496 216864 70508
rect 216784 70468 216864 70496
rect 216784 70372 216812 70468
rect 216858 70456 216864 70468
rect 216916 70456 216922 70508
rect 219544 70372 219572 70536
rect 219618 70524 219624 70536
rect 219676 70524 219682 70576
rect 346118 70388 346124 70440
rect 346176 70428 346182 70440
rect 346176 70400 346256 70428
rect 346176 70388 346182 70400
rect 346228 70372 346256 70400
rect 191926 70320 191932 70372
rect 191984 70320 191990 70372
rect 194686 70320 194692 70372
rect 194744 70320 194750 70372
rect 216766 70320 216772 70372
rect 216824 70320 216830 70372
rect 219526 70320 219532 70372
rect 219584 70320 219590 70372
rect 346210 70320 346216 70372
rect 346268 70320 346274 70372
rect 150710 70292 150716 70304
rect 150671 70264 150716 70292
rect 150710 70252 150716 70264
rect 150768 70252 150774 70304
rect 303890 70224 303896 70236
rect 303851 70196 303896 70224
rect 303890 70184 303896 70196
rect 303948 70184 303954 70236
rect 248322 67736 248328 67788
rect 248380 67736 248386 67788
rect 265066 67736 265072 67788
rect 265124 67736 265130 67788
rect 162946 67668 162952 67720
rect 163004 67708 163010 67720
rect 163222 67708 163228 67720
rect 163004 67680 163228 67708
rect 163004 67668 163010 67680
rect 163222 67668 163228 67680
rect 163280 67668 163286 67720
rect 248340 67652 248368 67736
rect 252741 67711 252799 67717
rect 252741 67677 252753 67711
rect 252787 67708 252799 67711
rect 252830 67708 252836 67720
rect 252787 67680 252836 67708
rect 252787 67677 252799 67680
rect 252741 67671 252799 67677
rect 252830 67668 252836 67680
rect 252888 67668 252894 67720
rect 265084 67652 265112 67736
rect 307938 67668 307944 67720
rect 307996 67708 308002 67720
rect 308030 67708 308036 67720
rect 307996 67680 308036 67708
rect 307996 67668 308002 67680
rect 308030 67668 308036 67680
rect 308088 67668 308094 67720
rect 154758 67640 154764 67652
rect 154719 67612 154764 67640
rect 154758 67600 154764 67612
rect 154816 67600 154822 67652
rect 173986 67600 173992 67652
rect 174044 67640 174050 67652
rect 174078 67640 174084 67652
rect 174044 67612 174084 67640
rect 174044 67600 174050 67612
rect 174078 67600 174084 67612
rect 174136 67600 174142 67652
rect 222470 67600 222476 67652
rect 222528 67640 222534 67652
rect 222562 67640 222568 67652
rect 222528 67612 222568 67640
rect 222528 67600 222534 67612
rect 222562 67600 222568 67612
rect 222620 67600 222626 67652
rect 248322 67600 248328 67652
rect 248380 67600 248386 67652
rect 265066 67600 265072 67652
rect 265124 67600 265130 67652
rect 357250 67640 357256 67652
rect 357211 67612 357256 67640
rect 357250 67600 357256 67612
rect 357308 67600 357314 67652
rect 423214 67600 423220 67652
rect 423272 67640 423278 67652
rect 423306 67640 423312 67652
rect 423272 67612 423312 67640
rect 423272 67600 423278 67612
rect 423306 67600 423312 67612
rect 423364 67600 423370 67652
rect 236270 67532 236276 67584
rect 236328 67572 236334 67584
rect 236362 67572 236368 67584
rect 236328 67544 236368 67572
rect 236328 67532 236334 67544
rect 236362 67532 236368 67544
rect 236420 67532 236426 67584
rect 237558 67532 237564 67584
rect 237616 67572 237622 67584
rect 237650 67572 237656 67584
rect 237616 67544 237656 67572
rect 237616 67532 237622 67544
rect 237650 67532 237656 67544
rect 237708 67532 237714 67584
rect 307662 67532 307668 67584
rect 307720 67572 307726 67584
rect 307938 67572 307944 67584
rect 307720 67544 307944 67572
rect 307720 67532 307726 67544
rect 307938 67532 307944 67544
rect 307996 67532 308002 67584
rect 424686 67572 424692 67584
rect 424647 67544 424692 67572
rect 424686 67532 424692 67544
rect 424744 67532 424750 67584
rect 208486 66348 208492 66360
rect 208447 66320 208492 66348
rect 208486 66308 208492 66320
rect 208544 66308 208550 66360
rect 190638 66280 190644 66292
rect 190599 66252 190644 66280
rect 190638 66240 190644 66252
rect 190696 66240 190702 66292
rect 207017 66283 207075 66289
rect 207017 66249 207029 66283
rect 207063 66280 207075 66283
rect 207106 66280 207112 66292
rect 207063 66252 207112 66280
rect 207063 66249 207075 66252
rect 207017 66243 207075 66249
rect 207106 66240 207112 66252
rect 207164 66240 207170 66292
rect 252738 66280 252744 66292
rect 252699 66252 252744 66280
rect 252738 66240 252744 66252
rect 252796 66240 252802 66292
rect 284386 66240 284392 66292
rect 284444 66280 284450 66292
rect 284478 66280 284484 66292
rect 284444 66252 284484 66280
rect 284444 66240 284450 66252
rect 284478 66240 284484 66252
rect 284536 66240 284542 66292
rect 384669 66283 384727 66289
rect 384669 66249 384681 66283
rect 384715 66280 384727 66283
rect 384758 66280 384764 66292
rect 384715 66252 384764 66280
rect 384715 66249 384727 66252
rect 384669 66243 384727 66249
rect 384758 66240 384764 66252
rect 384816 66240 384822 66292
rect 162857 66215 162915 66221
rect 162857 66181 162869 66215
rect 162903 66212 162915 66215
rect 162946 66212 162952 66224
rect 162903 66184 162952 66212
rect 162903 66181 162915 66184
rect 162857 66175 162915 66181
rect 162946 66172 162952 66184
rect 163004 66172 163010 66224
rect 168469 66215 168527 66221
rect 168469 66181 168481 66215
rect 168515 66212 168527 66215
rect 168558 66212 168564 66224
rect 168515 66184 168564 66212
rect 168515 66181 168527 66184
rect 168469 66175 168527 66181
rect 168558 66172 168564 66184
rect 168616 66172 168622 66224
rect 191926 66172 191932 66224
rect 191984 66212 191990 66224
rect 192110 66212 192116 66224
rect 191984 66184 192116 66212
rect 191984 66172 191990 66184
rect 192110 66172 192116 66184
rect 192168 66172 192174 66224
rect 219526 66212 219532 66224
rect 219487 66184 219532 66212
rect 219526 66172 219532 66184
rect 219584 66172 219590 66224
rect 238662 66212 238668 66224
rect 238623 66184 238668 66212
rect 238662 66172 238668 66184
rect 238720 66172 238726 66224
rect 248322 66212 248328 66224
rect 248283 66184 248328 66212
rect 248322 66172 248328 66184
rect 248380 66172 248386 66224
rect 263689 66215 263747 66221
rect 263689 66181 263701 66215
rect 263735 66212 263747 66215
rect 263778 66212 263784 66224
rect 263735 66184 263784 66212
rect 263735 66181 263747 66184
rect 263689 66175 263747 66181
rect 263778 66172 263784 66184
rect 263836 66172 263842 66224
rect 265066 66212 265072 66224
rect 265027 66184 265072 66212
rect 265066 66172 265072 66184
rect 265124 66172 265130 66224
rect 374270 66212 374276 66224
rect 374231 66184 374276 66212
rect 374270 66172 374276 66184
rect 374328 66172 374334 66224
rect 379146 66212 379152 66224
rect 379107 66184 379152 66212
rect 379146 66172 379152 66184
rect 379204 66172 379210 66224
rect 211249 64991 211307 64997
rect 211249 64957 211261 64991
rect 211295 64988 211307 64991
rect 211338 64988 211344 65000
rect 211295 64960 211344 64988
rect 211295 64957 211307 64960
rect 211249 64951 211307 64957
rect 211338 64948 211344 64960
rect 211396 64948 211402 65000
rect 246022 64920 246028 64932
rect 245983 64892 246028 64920
rect 246022 64880 246028 64892
rect 246080 64880 246086 64932
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 21358 64852 21364 64864
rect 3384 64824 21364 64852
rect 3384 64812 3390 64824
rect 21358 64812 21364 64824
rect 21416 64812 21422 64864
rect 150710 64852 150716 64864
rect 150671 64824 150716 64852
rect 150710 64812 150716 64824
rect 150768 64812 150774 64864
rect 189166 64852 189172 64864
rect 189127 64824 189172 64852
rect 189166 64812 189172 64824
rect 189224 64812 189230 64864
rect 207106 64852 207112 64864
rect 207067 64824 207112 64852
rect 207106 64812 207112 64824
rect 207164 64812 207170 64864
rect 208486 64852 208492 64864
rect 208447 64824 208492 64852
rect 208486 64812 208492 64824
rect 208544 64812 208550 64864
rect 211338 64852 211344 64864
rect 211299 64824 211344 64852
rect 211338 64812 211344 64824
rect 211396 64812 211402 64864
rect 218238 64852 218244 64864
rect 218199 64824 218244 64852
rect 218238 64812 218244 64824
rect 218296 64812 218302 64864
rect 223669 64855 223727 64861
rect 223669 64821 223681 64855
rect 223715 64852 223727 64855
rect 223758 64852 223764 64864
rect 223715 64824 223764 64852
rect 223715 64821 223727 64824
rect 223669 64815 223727 64821
rect 223758 64812 223764 64824
rect 223816 64812 223822 64864
rect 577590 64676 577596 64728
rect 577648 64716 577654 64728
rect 580350 64716 580356 64728
rect 577648 64688 580356 64716
rect 577648 64676 577654 64688
rect 580350 64676 580356 64688
rect 580408 64676 580414 64728
rect 190638 64648 190644 64660
rect 190599 64620 190644 64648
rect 190638 64608 190644 64620
rect 190696 64608 190702 64660
rect 198182 63492 198188 63504
rect 198143 63464 198188 63492
rect 198182 63452 198188 63464
rect 198240 63452 198246 63504
rect 177942 62772 177948 62824
rect 178000 62812 178006 62824
rect 178218 62812 178224 62824
rect 178000 62784 178224 62812
rect 178000 62772 178006 62784
rect 178218 62772 178224 62784
rect 178276 62772 178282 62824
rect 403434 62092 403440 62144
rect 403492 62132 403498 62144
rect 403526 62132 403532 62144
rect 403492 62104 403532 62132
rect 403492 62092 403498 62104
rect 403526 62092 403532 62104
rect 403584 62092 403590 62144
rect 284386 60800 284392 60852
rect 284444 60800 284450 60852
rect 284404 60716 284432 60800
rect 169846 60664 169852 60716
rect 169904 60704 169910 60716
rect 170030 60704 170036 60716
rect 169904 60676 170036 60704
rect 169904 60664 169910 60676
rect 170030 60664 170036 60676
rect 170088 60664 170094 60716
rect 258166 60664 258172 60716
rect 258224 60704 258230 60716
rect 258350 60704 258356 60716
rect 258224 60676 258356 60704
rect 258224 60664 258230 60676
rect 258350 60664 258356 60676
rect 258408 60664 258414 60716
rect 265066 60704 265072 60716
rect 265027 60676 265072 60704
rect 265066 60664 265072 60676
rect 265124 60664 265130 60716
rect 278866 60664 278872 60716
rect 278924 60664 278930 60716
rect 284386 60664 284392 60716
rect 284444 60664 284450 60716
rect 278884 60636 278912 60664
rect 278958 60636 278964 60648
rect 278884 60608 278964 60636
rect 278958 60596 278964 60608
rect 279016 60596 279022 60648
rect 252462 58012 252468 58064
rect 252520 58012 252526 58064
rect 423214 58012 423220 58064
rect 423272 58052 423278 58064
rect 423490 58052 423496 58064
rect 423272 58024 423496 58052
rect 423272 58012 423278 58024
rect 423490 58012 423496 58024
rect 423548 58012 423554 58064
rect 214098 57944 214104 57996
rect 214156 57984 214162 57996
rect 214190 57984 214196 57996
rect 214156 57956 214196 57984
rect 214156 57944 214162 57956
rect 214190 57944 214196 57956
rect 214248 57944 214254 57996
rect 229278 57944 229284 57996
rect 229336 57984 229342 57996
rect 229370 57984 229376 57996
rect 229336 57956 229376 57984
rect 229336 57944 229342 57956
rect 229370 57944 229376 57956
rect 229428 57944 229434 57996
rect 252480 57928 252508 58012
rect 303614 57944 303620 57996
rect 303672 57984 303678 57996
rect 303890 57984 303896 57996
rect 303672 57956 303896 57984
rect 303672 57944 303678 57956
rect 303890 57944 303896 57956
rect 303948 57944 303954 57996
rect 424689 57987 424747 57993
rect 424689 57953 424701 57987
rect 424735 57984 424747 57987
rect 424778 57984 424784 57996
rect 424735 57956 424784 57984
rect 424735 57953 424747 57956
rect 424689 57947 424747 57953
rect 424778 57944 424784 57956
rect 424836 57944 424842 57996
rect 154758 57916 154764 57928
rect 154719 57888 154764 57916
rect 154758 57876 154764 57888
rect 154816 57876 154822 57928
rect 173989 57919 174047 57925
rect 173989 57885 174001 57919
rect 174035 57916 174047 57919
rect 174078 57916 174084 57928
rect 174035 57888 174084 57916
rect 174035 57885 174047 57888
rect 173989 57879 174047 57885
rect 174078 57876 174084 57888
rect 174136 57876 174142 57928
rect 178218 57916 178224 57928
rect 178179 57888 178224 57916
rect 178218 57876 178224 57888
rect 178276 57876 178282 57928
rect 252462 57876 252468 57928
rect 252520 57876 252526 57928
rect 258169 57919 258227 57925
rect 258169 57885 258181 57919
rect 258215 57916 258227 57919
rect 258350 57916 258356 57928
rect 258215 57888 258356 57916
rect 258215 57885 258227 57888
rect 258169 57879 258227 57885
rect 258350 57876 258356 57888
rect 258408 57876 258414 57928
rect 307846 57916 307852 57928
rect 307807 57888 307852 57916
rect 307846 57876 307852 57888
rect 307904 57876 307910 57928
rect 357253 57919 357311 57925
rect 357253 57885 357265 57919
rect 357299 57916 357311 57919
rect 357342 57916 357348 57928
rect 357299 57888 357348 57916
rect 357299 57885 357311 57888
rect 357253 57879 357311 57885
rect 357342 57876 357348 57888
rect 357400 57876 357406 57928
rect 252370 56992 252376 57044
rect 252428 57032 252434 57044
rect 252830 57032 252836 57044
rect 252428 57004 252836 57032
rect 252428 56992 252434 57004
rect 252830 56992 252836 57004
rect 252888 56992 252894 57044
rect 246022 56692 246028 56704
rect 245856 56664 246028 56692
rect 162854 56584 162860 56636
rect 162912 56624 162918 56636
rect 168466 56624 168472 56636
rect 162912 56596 162957 56624
rect 168427 56596 168472 56624
rect 162912 56584 162918 56596
rect 168466 56584 168472 56596
rect 168524 56584 168530 56636
rect 190641 56627 190699 56633
rect 190641 56593 190653 56627
rect 190687 56624 190699 56627
rect 190730 56624 190736 56636
rect 190687 56596 190736 56624
rect 190687 56593 190699 56596
rect 190641 56587 190699 56593
rect 190730 56584 190736 56596
rect 190788 56584 190794 56636
rect 245856 56568 245884 56664
rect 246022 56652 246028 56664
rect 246080 56652 246086 56704
rect 379146 56692 379152 56704
rect 379107 56664 379152 56692
rect 379146 56652 379152 56664
rect 379204 56652 379210 56704
rect 247126 56584 247132 56636
rect 247184 56624 247190 56636
rect 247310 56624 247316 56636
rect 247184 56596 247316 56624
rect 247184 56584 247190 56596
rect 247310 56584 247316 56596
rect 247368 56584 247374 56636
rect 248322 56624 248328 56636
rect 248283 56596 248328 56624
rect 248322 56584 248328 56596
rect 248380 56584 248386 56636
rect 374270 56624 374276 56636
rect 374231 56596 374276 56624
rect 374270 56584 374276 56596
rect 374328 56584 374334 56636
rect 216858 56516 216864 56568
rect 216916 56556 216922 56568
rect 216950 56556 216956 56568
rect 216916 56528 216956 56556
rect 216916 56516 216922 56528
rect 216950 56516 216956 56528
rect 217008 56516 217014 56568
rect 245838 56516 245844 56568
rect 245896 56516 245902 56568
rect 379146 56556 379152 56568
rect 379107 56528 379152 56556
rect 379146 56516 379152 56528
rect 379204 56516 379210 56568
rect 207106 56352 207112 56364
rect 207067 56324 207112 56352
rect 207106 56312 207112 56324
rect 207164 56312 207170 56364
rect 192021 55335 192079 55341
rect 192021 55301 192033 55335
rect 192067 55332 192079 55335
rect 192110 55332 192116 55344
rect 192067 55304 192116 55332
rect 192067 55301 192079 55304
rect 192021 55295 192079 55301
rect 192110 55292 192116 55304
rect 192168 55292 192174 55344
rect 194686 55264 194692 55276
rect 194647 55236 194692 55264
rect 194686 55224 194692 55236
rect 194744 55224 194750 55276
rect 208486 55264 208492 55276
rect 208447 55236 208492 55264
rect 208486 55224 208492 55236
rect 208544 55224 208550 55276
rect 211341 55267 211399 55273
rect 211341 55233 211353 55267
rect 211387 55264 211399 55267
rect 211522 55264 211528 55276
rect 211387 55236 211528 55264
rect 211387 55233 211399 55236
rect 211341 55227 211399 55233
rect 211522 55224 211528 55236
rect 211580 55224 211586 55276
rect 223666 55264 223672 55276
rect 223627 55236 223672 55264
rect 223666 55224 223672 55236
rect 223724 55224 223730 55276
rect 226521 55267 226579 55273
rect 226521 55233 226533 55267
rect 226567 55264 226579 55267
rect 226702 55264 226708 55276
rect 226567 55236 226708 55264
rect 226567 55233 226579 55236
rect 226521 55227 226579 55233
rect 226702 55224 226708 55236
rect 226760 55224 226766 55276
rect 216950 55196 216956 55208
rect 216911 55168 216956 55196
rect 216950 55156 216956 55168
rect 217008 55156 217014 55208
rect 192018 53836 192024 53848
rect 191979 53808 192024 53836
rect 192018 53796 192024 53808
rect 192076 53796 192082 53848
rect 194686 53836 194692 53848
rect 194647 53808 194692 53836
rect 194686 53796 194692 53808
rect 194744 53796 194750 53848
rect 198182 53836 198188 53848
rect 198143 53808 198188 53836
rect 198182 53796 198188 53808
rect 198240 53796 198246 53848
rect 403618 52436 403624 52488
rect 403676 52476 403682 52488
rect 403710 52476 403716 52488
rect 403676 52448 403716 52476
rect 403676 52436 403682 52448
rect 403710 52436 403716 52448
rect 403768 52436 403774 52488
rect 179506 51144 179512 51196
rect 179564 51144 179570 51196
rect 270586 51184 270592 51196
rect 270547 51156 270592 51184
rect 270586 51144 270592 51156
rect 270644 51144 270650 51196
rect 179524 51060 179552 51144
rect 196250 51116 196256 51128
rect 196176 51088 196256 51116
rect 196176 51060 196204 51088
rect 196250 51076 196256 51088
rect 196308 51076 196314 51128
rect 271877 51119 271935 51125
rect 271877 51085 271889 51119
rect 271923 51116 271935 51119
rect 272058 51116 272064 51128
rect 271923 51088 272064 51116
rect 271923 51085 271935 51088
rect 271877 51079 271935 51085
rect 272058 51076 272064 51088
rect 272116 51076 272122 51128
rect 284386 51116 284392 51128
rect 284312 51088 284392 51116
rect 284312 51060 284340 51088
rect 284386 51076 284392 51088
rect 284444 51076 284450 51128
rect 179506 51008 179512 51060
rect 179564 51008 179570 51060
rect 196158 51008 196164 51060
rect 196216 51008 196222 51060
rect 252370 51008 252376 51060
rect 252428 51048 252434 51060
rect 252738 51048 252744 51060
rect 252428 51020 252744 51048
rect 252428 51008 252434 51020
rect 252738 51008 252744 51020
rect 252796 51008 252802 51060
rect 284294 51008 284300 51060
rect 284352 51008 284358 51060
rect 154758 48396 154764 48408
rect 154719 48368 154764 48396
rect 154758 48356 154764 48368
rect 154816 48356 154822 48408
rect 173986 48328 173992 48340
rect 173947 48300 173992 48328
rect 173986 48288 173992 48300
rect 174044 48288 174050 48340
rect 178221 48331 178279 48337
rect 178221 48297 178233 48331
rect 178267 48328 178279 48331
rect 178310 48328 178316 48340
rect 178267 48300 178316 48328
rect 178267 48297 178279 48300
rect 178221 48291 178279 48297
rect 178310 48288 178316 48300
rect 178368 48288 178374 48340
rect 190638 48288 190644 48340
rect 190696 48328 190702 48340
rect 190730 48328 190736 48340
rect 190696 48300 190736 48328
rect 190696 48288 190702 48300
rect 190730 48288 190736 48300
rect 190788 48288 190794 48340
rect 238662 48328 238668 48340
rect 238623 48300 238668 48328
rect 238662 48288 238668 48300
rect 238720 48288 238726 48340
rect 258166 48328 258172 48340
rect 258127 48300 258172 48328
rect 258166 48288 258172 48300
rect 258224 48288 258230 48340
rect 263686 48328 263692 48340
rect 263647 48300 263692 48328
rect 263686 48288 263692 48300
rect 263744 48288 263750 48340
rect 270586 48328 270592 48340
rect 270547 48300 270592 48328
rect 270586 48288 270592 48300
rect 270644 48288 270650 48340
rect 271874 48328 271880 48340
rect 271835 48300 271880 48328
rect 271874 48288 271880 48300
rect 271932 48288 271938 48340
rect 307849 48331 307907 48337
rect 307849 48297 307861 48331
rect 307895 48328 307907 48331
rect 307938 48328 307944 48340
rect 307895 48300 307944 48328
rect 307895 48297 307907 48300
rect 307849 48291 307907 48297
rect 307938 48288 307944 48300
rect 307996 48288 308002 48340
rect 346210 48288 346216 48340
rect 346268 48328 346274 48340
rect 346302 48328 346308 48340
rect 346268 48300 346308 48328
rect 346268 48288 346274 48300
rect 346302 48288 346308 48300
rect 346360 48288 346366 48340
rect 357250 48328 357256 48340
rect 357211 48300 357256 48328
rect 357250 48288 357256 48300
rect 357308 48288 357314 48340
rect 384758 48288 384764 48340
rect 384816 48328 384822 48340
rect 384850 48328 384856 48340
rect 384816 48300 384856 48328
rect 384816 48288 384822 48300
rect 384850 48288 384856 48300
rect 384908 48288 384914 48340
rect 403710 48288 403716 48340
rect 403768 48328 403774 48340
rect 403802 48328 403808 48340
rect 403768 48300 403808 48328
rect 403768 48288 403774 48300
rect 403802 48288 403808 48300
rect 403860 48288 403866 48340
rect 154758 48260 154764 48272
rect 154719 48232 154764 48260
rect 154758 48220 154764 48232
rect 154816 48220 154822 48272
rect 225046 48220 225052 48272
rect 225104 48260 225110 48272
rect 225138 48260 225144 48272
rect 225104 48232 225144 48260
rect 225104 48220 225110 48232
rect 225138 48220 225144 48232
rect 225196 48220 225202 48272
rect 234801 48263 234859 48269
rect 234801 48229 234813 48263
rect 234847 48260 234859 48263
rect 234890 48260 234896 48272
rect 234847 48232 234896 48260
rect 234847 48229 234859 48232
rect 234801 48223 234859 48229
rect 234890 48220 234896 48232
rect 234948 48220 234954 48272
rect 236270 48220 236276 48272
rect 236328 48260 236334 48272
rect 236362 48260 236368 48272
rect 236328 48232 236368 48260
rect 236328 48220 236334 48232
rect 236362 48220 236368 48232
rect 236420 48220 236426 48272
rect 237558 48220 237564 48272
rect 237616 48260 237622 48272
rect 237650 48260 237656 48272
rect 237616 48232 237656 48260
rect 237616 48220 237622 48232
rect 237650 48220 237656 48232
rect 237708 48220 237714 48272
rect 284294 48220 284300 48272
rect 284352 48260 284358 48272
rect 284481 48263 284539 48269
rect 284481 48260 284493 48263
rect 284352 48232 284493 48260
rect 284352 48220 284358 48232
rect 284481 48229 284493 48232
rect 284527 48229 284539 48263
rect 424686 48260 424692 48272
rect 424647 48232 424692 48260
rect 284481 48223 284539 48229
rect 424686 48220 424692 48232
rect 424744 48220 424750 48272
rect 211249 47311 211307 47317
rect 211249 47277 211261 47311
rect 211295 47308 211307 47311
rect 211522 47308 211528 47320
rect 211295 47280 211528 47308
rect 211295 47277 211307 47280
rect 211249 47271 211307 47277
rect 211522 47268 211528 47280
rect 211580 47268 211586 47320
rect 189169 46971 189227 46977
rect 189169 46937 189181 46971
rect 189215 46968 189227 46971
rect 189350 46968 189356 46980
rect 189215 46940 189356 46968
rect 189215 46937 189227 46940
rect 189169 46931 189227 46937
rect 189350 46928 189356 46940
rect 189408 46928 189414 46980
rect 218238 46968 218244 46980
rect 218199 46940 218244 46968
rect 218238 46928 218244 46940
rect 218296 46928 218302 46980
rect 219526 46968 219532 46980
rect 219487 46940 219532 46968
rect 219526 46928 219532 46940
rect 219584 46928 219590 46980
rect 379149 46971 379207 46977
rect 379149 46937 379161 46971
rect 379195 46968 379207 46971
rect 379238 46968 379244 46980
rect 379195 46940 379244 46968
rect 379195 46937 379207 46940
rect 379149 46931 379207 46937
rect 379238 46928 379244 46940
rect 379296 46928 379302 46980
rect 168558 46900 168564 46912
rect 168519 46872 168564 46900
rect 168558 46860 168564 46872
rect 168616 46860 168622 46912
rect 169846 46900 169852 46912
rect 169807 46872 169852 46900
rect 169846 46860 169852 46872
rect 169904 46860 169910 46912
rect 207106 46900 207112 46912
rect 207067 46872 207112 46900
rect 207106 46860 207112 46872
rect 207164 46860 207170 46912
rect 214006 46860 214012 46912
rect 214064 46900 214070 46912
rect 214101 46903 214159 46909
rect 214101 46900 214113 46903
rect 214064 46872 214113 46900
rect 214064 46860 214070 46872
rect 214101 46869 214113 46872
rect 214147 46869 214159 46903
rect 214101 46863 214159 46869
rect 238573 46903 238631 46909
rect 238573 46869 238585 46903
rect 238619 46900 238631 46903
rect 238662 46900 238668 46912
rect 238619 46872 238668 46900
rect 238619 46869 238631 46872
rect 238573 46863 238631 46869
rect 238662 46860 238668 46872
rect 238720 46860 238726 46912
rect 245838 46860 245844 46912
rect 245896 46860 245902 46912
rect 247126 46860 247132 46912
rect 247184 46900 247190 46912
rect 247402 46900 247408 46912
rect 247184 46872 247408 46900
rect 247184 46860 247190 46872
rect 247402 46860 247408 46872
rect 247460 46860 247466 46912
rect 248322 46900 248328 46912
rect 248283 46872 248328 46900
rect 248322 46860 248328 46872
rect 248380 46860 248386 46912
rect 374270 46900 374276 46912
rect 374231 46872 374276 46900
rect 374270 46860 374276 46872
rect 374328 46860 374334 46912
rect 245746 46792 245752 46844
rect 245804 46832 245810 46844
rect 245856 46832 245884 46860
rect 245804 46804 245884 46832
rect 245804 46792 245810 46804
rect 194686 45772 194692 45824
rect 194744 45812 194750 45824
rect 194744 45784 194824 45812
rect 194744 45772 194750 45784
rect 150526 45636 150532 45688
rect 150584 45676 150590 45688
rect 150710 45676 150716 45688
rect 150584 45648 150716 45676
rect 150584 45636 150590 45648
rect 150710 45636 150716 45648
rect 150768 45636 150774 45688
rect 194796 45620 194824 45784
rect 194778 45568 194784 45620
rect 194836 45568 194842 45620
rect 211246 45608 211252 45620
rect 211207 45580 211252 45608
rect 211246 45568 211252 45580
rect 211304 45568 211310 45620
rect 216950 45608 216956 45620
rect 216911 45580 216956 45608
rect 216950 45568 216956 45580
rect 217008 45568 217014 45620
rect 196158 45500 196164 45552
rect 196216 45540 196222 45552
rect 196342 45540 196348 45552
rect 196216 45512 196348 45540
rect 196216 45500 196222 45512
rect 196342 45500 196348 45512
rect 196400 45500 196406 45552
rect 218238 45500 218244 45552
rect 218296 45540 218302 45552
rect 218330 45540 218336 45552
rect 218296 45512 218336 45540
rect 218296 45500 218302 45512
rect 218330 45500 218336 45512
rect 218388 45500 218394 45552
rect 219437 45543 219495 45549
rect 219437 45509 219449 45543
rect 219483 45540 219495 45543
rect 219526 45540 219532 45552
rect 219483 45512 219532 45540
rect 219483 45509 219495 45512
rect 219437 45503 219495 45509
rect 219526 45500 219532 45512
rect 219584 45500 219590 45552
rect 245746 45540 245752 45552
rect 245707 45512 245752 45540
rect 245746 45500 245752 45512
rect 245804 45500 245810 45552
rect 247402 45540 247408 45552
rect 247363 45512 247408 45540
rect 247402 45500 247408 45512
rect 247460 45500 247466 45552
rect 154761 43707 154819 43713
rect 154761 43673 154773 43707
rect 154807 43704 154819 43707
rect 155034 43704 155040 43716
rect 154807 43676 155040 43704
rect 154807 43673 154819 43676
rect 154761 43667 154819 43673
rect 155034 43664 155040 43676
rect 155092 43664 155098 43716
rect 208578 42072 208584 42084
rect 208539 42044 208584 42072
rect 208578 42032 208584 42044
rect 208636 42032 208642 42084
rect 222470 42072 222476 42084
rect 222431 42044 222476 42072
rect 222470 42032 222476 42044
rect 222528 42032 222534 42084
rect 223758 42072 223764 42084
rect 223719 42044 223764 42072
rect 223758 42032 223764 42044
rect 223816 42032 223822 42084
rect 178126 41352 178132 41404
rect 178184 41392 178190 41404
rect 178310 41392 178316 41404
rect 178184 41364 178316 41392
rect 178184 41352 178190 41364
rect 178310 41352 178316 41364
rect 178368 41352 178374 41404
rect 284478 41392 284484 41404
rect 284439 41364 284484 41392
rect 284478 41352 284484 41364
rect 284536 41352 284542 41404
rect 340690 40196 340696 40248
rect 340748 40236 340754 40248
rect 340966 40236 340972 40248
rect 340748 40208 340972 40236
rect 340748 40196 340754 40208
rect 340966 40196 340972 40208
rect 341024 40196 341030 40248
rect 201494 40128 201500 40180
rect 201552 40168 201558 40180
rect 219342 40168 219348 40180
rect 201552 40140 219348 40168
rect 201552 40128 201558 40140
rect 219342 40128 219348 40140
rect 219400 40128 219406 40180
rect 321278 40128 321284 40180
rect 321336 40168 321342 40180
rect 321554 40168 321560 40180
rect 321336 40140 321560 40168
rect 321336 40128 321342 40140
rect 321554 40128 321560 40140
rect 321612 40128 321618 40180
rect 359918 40128 359924 40180
rect 359976 40168 359982 40180
rect 360194 40168 360200 40180
rect 359976 40140 360200 40168
rect 359976 40128 359982 40140
rect 360194 40128 360200 40140
rect 360252 40128 360258 40180
rect 444374 40060 444380 40112
rect 444432 40100 444438 40112
rect 447226 40100 447232 40112
rect 444432 40072 447232 40100
rect 444432 40060 444438 40072
rect 447226 40060 447232 40072
rect 447284 40060 447290 40112
rect 476022 40060 476028 40112
rect 476080 40100 476086 40112
rect 482922 40100 482928 40112
rect 476080 40072 482928 40100
rect 476080 40060 476086 40072
rect 482922 40060 482928 40072
rect 482980 40060 482986 40112
rect 258258 38768 258264 38820
rect 258316 38768 258322 38820
rect 258276 38684 258304 38768
rect 423306 38700 423312 38752
rect 423364 38740 423370 38752
rect 423490 38740 423496 38752
rect 423364 38712 423496 38740
rect 423364 38700 423370 38712
rect 423490 38700 423496 38712
rect 423548 38700 423554 38752
rect 189258 38632 189264 38684
rect 189316 38672 189322 38684
rect 189350 38672 189356 38684
rect 189316 38644 189356 38672
rect 189316 38632 189322 38644
rect 189350 38632 189356 38644
rect 189408 38632 189414 38684
rect 190638 38632 190644 38684
rect 190696 38672 190702 38684
rect 190730 38672 190736 38684
rect 190696 38644 190736 38672
rect 190696 38632 190702 38644
rect 190730 38632 190736 38644
rect 190788 38632 190794 38684
rect 234798 38672 234804 38684
rect 234759 38644 234804 38672
rect 234798 38632 234804 38644
rect 234856 38632 234862 38684
rect 252646 38632 252652 38684
rect 252704 38672 252710 38684
rect 252830 38672 252836 38684
rect 252704 38644 252836 38672
rect 252704 38632 252710 38644
rect 252830 38632 252836 38644
rect 252888 38632 252894 38684
rect 258258 38632 258264 38684
rect 258316 38632 258322 38684
rect 264974 38632 264980 38684
rect 265032 38672 265038 38684
rect 265066 38672 265072 38684
rect 265032 38644 265072 38672
rect 265032 38632 265038 38644
rect 265066 38632 265072 38644
rect 265124 38632 265130 38684
rect 384666 38632 384672 38684
rect 384724 38672 384730 38684
rect 384758 38672 384764 38684
rect 384724 38644 384764 38672
rect 384724 38632 384730 38644
rect 384758 38632 384764 38644
rect 384816 38632 384822 38684
rect 424689 38675 424747 38681
rect 424689 38641 424701 38675
rect 424735 38672 424747 38675
rect 424778 38672 424784 38684
rect 424735 38644 424784 38672
rect 424735 38641 424747 38644
rect 424689 38635 424747 38641
rect 424778 38632 424784 38644
rect 424836 38632 424842 38684
rect 284389 38607 284447 38613
rect 284389 38573 284401 38607
rect 284435 38604 284447 38607
rect 284478 38604 284484 38616
rect 284435 38576 284484 38604
rect 284435 38573 284447 38576
rect 284389 38567 284447 38573
rect 284478 38564 284484 38576
rect 284536 38564 284542 38616
rect 307941 38607 307999 38613
rect 307941 38573 307953 38607
rect 307987 38604 307999 38607
rect 308030 38604 308036 38616
rect 307987 38576 308036 38604
rect 307987 38573 307999 38576
rect 307941 38567 307999 38573
rect 308030 38564 308036 38576
rect 308088 38564 308094 38616
rect 357253 38607 357311 38613
rect 357253 38573 357265 38607
rect 357299 38604 357311 38607
rect 357342 38604 357348 38616
rect 357299 38576 357348 38604
rect 357299 38573 357311 38576
rect 357253 38567 357311 38573
rect 357342 38564 357348 38576
rect 357400 38564 357406 38616
rect 403802 38604 403808 38616
rect 403763 38576 403808 38604
rect 403802 38564 403808 38576
rect 403860 38564 403866 38616
rect 168561 37315 168619 37321
rect 168561 37281 168573 37315
rect 168607 37312 168619 37315
rect 168650 37312 168656 37324
rect 168607 37284 168656 37312
rect 168607 37281 168619 37284
rect 168561 37275 168619 37281
rect 168650 37272 168656 37284
rect 168708 37272 168714 37324
rect 169849 37315 169907 37321
rect 169849 37281 169861 37315
rect 169895 37312 169907 37315
rect 169938 37312 169944 37324
rect 169895 37284 169944 37312
rect 169895 37281 169907 37284
rect 169849 37275 169907 37281
rect 169938 37272 169944 37284
rect 169996 37272 170002 37324
rect 207109 37315 207167 37321
rect 207109 37281 207121 37315
rect 207155 37281 207167 37315
rect 207109 37275 207167 37281
rect 238573 37315 238631 37321
rect 238573 37281 238585 37315
rect 238619 37312 238631 37315
rect 238662 37312 238668 37324
rect 238619 37284 238668 37312
rect 238619 37281 238631 37284
rect 238573 37275 238631 37281
rect 190641 37247 190699 37253
rect 190641 37213 190653 37247
rect 190687 37244 190699 37247
rect 190730 37244 190736 37256
rect 190687 37216 190736 37244
rect 190687 37213 190699 37216
rect 190641 37207 190699 37213
rect 190730 37204 190736 37216
rect 190788 37204 190794 37256
rect 207124 37176 207152 37275
rect 238662 37272 238668 37284
rect 238720 37272 238726 37324
rect 248322 37312 248328 37324
rect 248283 37284 248328 37312
rect 248322 37272 248328 37284
rect 248380 37272 248386 37324
rect 374270 37312 374276 37324
rect 374231 37284 374276 37312
rect 374270 37272 374276 37284
rect 374328 37272 374334 37324
rect 379146 37272 379152 37324
rect 379204 37312 379210 37324
rect 379238 37312 379244 37324
rect 379204 37284 379244 37312
rect 379204 37272 379210 37284
rect 379238 37272 379244 37284
rect 379296 37272 379302 37324
rect 219437 37247 219495 37253
rect 219437 37213 219449 37247
rect 219483 37244 219495 37247
rect 219526 37244 219532 37256
rect 219483 37216 219532 37244
rect 219483 37213 219495 37216
rect 219437 37207 219495 37213
rect 219526 37204 219532 37216
rect 219584 37204 219590 37256
rect 247402 37244 247408 37256
rect 247363 37216 247408 37244
rect 247402 37204 247408 37216
rect 247460 37204 247466 37256
rect 207201 37179 207259 37185
rect 207201 37176 207213 37179
rect 207124 37148 207213 37176
rect 207201 37145 207213 37148
rect 207247 37145 207259 37179
rect 207201 37139 207259 37145
rect 194502 34484 194508 34536
rect 194560 34524 194566 34536
rect 194686 34524 194692 34536
rect 194560 34496 194692 34524
rect 194560 34484 194566 34496
rect 194686 34484 194692 34496
rect 194744 34484 194750 34536
rect 173989 33847 174047 33853
rect 173989 33813 174001 33847
rect 174035 33844 174047 33847
rect 174078 33844 174084 33856
rect 174035 33816 174084 33844
rect 174035 33813 174047 33816
rect 173989 33807 174047 33813
rect 174078 33804 174084 33816
rect 174136 33804 174142 33856
rect 213914 32376 213920 32428
rect 213972 32416 213978 32428
rect 214101 32419 214159 32425
rect 214101 32416 214113 32419
rect 213972 32388 214113 32416
rect 213972 32376 213978 32388
rect 214101 32385 214113 32388
rect 214147 32385 214159 32419
rect 214101 32379 214159 32385
rect 270586 31872 270592 31884
rect 270547 31844 270592 31872
rect 270586 31832 270592 31844
rect 270644 31832 270650 31884
rect 273346 31872 273352 31884
rect 273307 31844 273352 31872
rect 273346 31832 273352 31844
rect 273404 31832 273410 31884
rect 168650 31764 168656 31816
rect 168708 31764 168714 31816
rect 169938 31764 169944 31816
rect 169996 31764 170002 31816
rect 346118 31764 346124 31816
rect 346176 31764 346182 31816
rect 379330 31804 379336 31816
rect 379256 31776 379336 31804
rect 168668 31668 168696 31764
rect 169956 31680 169984 31764
rect 168742 31668 168748 31680
rect 168668 31640 168748 31668
rect 168742 31628 168748 31640
rect 168800 31628 168806 31680
rect 169938 31628 169944 31680
rect 169996 31628 170002 31680
rect 346136 31668 346164 31764
rect 357250 31736 357256 31748
rect 357211 31708 357256 31736
rect 357250 31696 357256 31708
rect 357308 31696 357314 31748
rect 379256 31680 379284 31776
rect 379330 31764 379336 31776
rect 379388 31764 379394 31816
rect 423306 31764 423312 31816
rect 423364 31764 423370 31816
rect 424778 31764 424784 31816
rect 424836 31804 424842 31816
rect 424962 31804 424968 31816
rect 424836 31776 424968 31804
rect 424836 31764 424842 31776
rect 424962 31764 424968 31776
rect 425020 31764 425026 31816
rect 384666 31696 384672 31748
rect 384724 31736 384730 31748
rect 384850 31736 384856 31748
rect 384724 31708 384856 31736
rect 384724 31696 384730 31708
rect 384850 31696 384856 31708
rect 384908 31696 384914 31748
rect 393958 31696 393964 31748
rect 394016 31736 394022 31748
rect 394142 31736 394148 31748
rect 394016 31708 394148 31736
rect 394016 31696 394022 31708
rect 394142 31696 394148 31708
rect 394200 31696 394206 31748
rect 346210 31668 346216 31680
rect 346136 31640 346216 31668
rect 346210 31628 346216 31640
rect 346268 31628 346274 31680
rect 379238 31628 379244 31680
rect 379296 31628 379302 31680
rect 423324 31668 423352 31764
rect 423398 31668 423404 31680
rect 423324 31640 423404 31668
rect 423398 31628 423404 31640
rect 423456 31628 423462 31680
rect 247402 31328 247408 31340
rect 247363 31300 247408 31328
rect 247402 31288 247408 31300
rect 247460 31288 247466 31340
rect 178310 31220 178316 31272
rect 178368 31220 178374 31272
rect 178328 31136 178356 31220
rect 178310 31084 178316 31136
rect 178368 31084 178374 31136
rect 577498 30268 577504 30320
rect 577556 30308 577562 30320
rect 579614 30308 579620 30320
rect 577556 30280 579620 30308
rect 577556 30268 577562 30280
rect 579614 30268 579620 30280
rect 579672 30268 579678 30320
rect 179598 29084 179604 29096
rect 179524 29056 179604 29084
rect 179524 29028 179552 29056
rect 179598 29044 179604 29056
rect 179656 29044 179662 29096
rect 236270 29084 236276 29096
rect 236196 29056 236276 29084
rect 236196 29028 236224 29056
rect 236270 29044 236276 29056
rect 236328 29044 236334 29096
rect 264974 29044 264980 29096
rect 265032 29084 265038 29096
rect 265066 29084 265072 29096
rect 265032 29056 265072 29084
rect 265032 29044 265038 29056
rect 265066 29044 265072 29056
rect 265124 29044 265130 29096
rect 173986 29016 173992 29028
rect 173947 28988 173992 29016
rect 173986 28976 173992 28988
rect 174044 28976 174050 29028
rect 179506 28976 179512 29028
rect 179564 28976 179570 29028
rect 205726 28976 205732 29028
rect 205784 29016 205790 29028
rect 205818 29016 205824 29028
rect 205784 28988 205824 29016
rect 205784 28976 205790 28988
rect 205818 28976 205824 28988
rect 205876 28976 205882 29028
rect 208578 29016 208584 29028
rect 208539 28988 208584 29016
rect 208578 28976 208584 28988
rect 208636 28976 208642 29028
rect 222473 29019 222531 29025
rect 222473 28985 222485 29019
rect 222519 29016 222531 29019
rect 222654 29016 222660 29028
rect 222519 28988 222660 29016
rect 222519 28985 222531 28988
rect 222473 28979 222531 28985
rect 222654 28976 222660 28988
rect 222712 28976 222718 29028
rect 223758 29016 223764 29028
rect 223719 28988 223764 29016
rect 223758 28976 223764 28988
rect 223816 28976 223822 29028
rect 229370 28976 229376 29028
rect 229428 29016 229434 29028
rect 229462 29016 229468 29028
rect 229428 28988 229468 29016
rect 229428 28976 229434 28988
rect 229462 28976 229468 28988
rect 229520 28976 229526 29028
rect 236178 28976 236184 29028
rect 236236 28976 236242 29028
rect 238662 29016 238668 29028
rect 238623 28988 238668 29016
rect 238662 28976 238668 28988
rect 238720 28976 238726 29028
rect 284386 29016 284392 29028
rect 284347 28988 284392 29016
rect 284386 28976 284392 28988
rect 284444 28976 284450 29028
rect 307938 29016 307944 29028
rect 307899 28988 307944 29016
rect 307938 28976 307944 28988
rect 307996 28976 308002 29028
rect 403805 29019 403863 29025
rect 403805 28985 403817 29019
rect 403851 29016 403863 29019
rect 403894 29016 403900 29028
rect 403851 28988 403900 29016
rect 403851 28985 403863 28988
rect 403805 28979 403863 28985
rect 403894 28976 403900 28988
rect 403952 28976 403958 29028
rect 271966 28908 271972 28960
rect 272024 28948 272030 28960
rect 272058 28948 272064 28960
rect 272024 28920 272064 28948
rect 272024 28908 272030 28920
rect 272058 28908 272064 28920
rect 272116 28908 272122 28960
rect 394053 28951 394111 28957
rect 394053 28917 394065 28951
rect 394099 28948 394111 28951
rect 394142 28948 394148 28960
rect 394099 28920 394148 28948
rect 394099 28917 394111 28920
rect 394053 28911 394111 28917
rect 394142 28908 394148 28920
rect 394200 28908 394206 28960
rect 150526 28296 150532 28348
rect 150584 28336 150590 28348
rect 150710 28336 150716 28348
rect 150584 28308 150716 28336
rect 150584 28296 150590 28308
rect 150710 28296 150716 28308
rect 150768 28296 150774 28348
rect 190638 27724 190644 27736
rect 190599 27696 190644 27724
rect 190638 27684 190644 27696
rect 190696 27684 190702 27736
rect 207106 27684 207112 27736
rect 207164 27724 207170 27736
rect 207201 27727 207259 27733
rect 207201 27724 207213 27727
rect 207164 27696 207213 27724
rect 207164 27684 207170 27696
rect 207201 27693 207213 27696
rect 207247 27693 207259 27727
rect 238662 27724 238668 27736
rect 238623 27696 238668 27724
rect 207201 27687 207259 27693
rect 238662 27684 238668 27696
rect 238720 27684 238726 27736
rect 191926 27656 191932 27668
rect 191887 27628 191932 27656
rect 191926 27616 191932 27628
rect 191984 27616 191990 27668
rect 198182 27616 198188 27668
rect 198240 27656 198246 27668
rect 198274 27656 198280 27668
rect 198240 27628 198280 27656
rect 198240 27616 198246 27628
rect 198274 27616 198280 27628
rect 198332 27616 198338 27668
rect 245749 27659 245807 27665
rect 245749 27625 245761 27659
rect 245795 27656 245807 27659
rect 245838 27656 245844 27668
rect 245795 27628 245844 27656
rect 245795 27625 245807 27628
rect 245749 27619 245807 27625
rect 245838 27616 245844 27628
rect 245896 27616 245902 27668
rect 247402 27656 247408 27668
rect 247363 27628 247408 27656
rect 247402 27616 247408 27628
rect 247460 27616 247466 27668
rect 270586 27656 270592 27668
rect 270547 27628 270592 27656
rect 270586 27616 270592 27628
rect 270644 27616 270650 27668
rect 273346 27656 273352 27668
rect 273307 27628 273352 27656
rect 273346 27616 273352 27628
rect 273404 27616 273410 27668
rect 168558 27548 168564 27600
rect 168616 27588 168622 27600
rect 168742 27588 168748 27600
rect 168616 27560 168748 27588
rect 168616 27548 168622 27560
rect 168742 27548 168748 27560
rect 168800 27548 168806 27600
rect 173986 27588 173992 27600
rect 173947 27560 173992 27588
rect 173986 27548 173992 27560
rect 174044 27548 174050 27600
rect 179506 27588 179512 27600
rect 179467 27560 179512 27588
rect 179506 27548 179512 27560
rect 179564 27548 179570 27600
rect 205818 27548 205824 27600
rect 205876 27588 205882 27600
rect 205910 27588 205916 27600
rect 205876 27560 205916 27588
rect 205876 27548 205882 27560
rect 205910 27548 205916 27560
rect 205968 27548 205974 27600
rect 207106 27588 207112 27600
rect 207067 27560 207112 27588
rect 207106 27548 207112 27560
rect 207164 27548 207170 27600
rect 211246 27548 211252 27600
rect 211304 27588 211310 27600
rect 211341 27591 211399 27597
rect 211341 27588 211353 27591
rect 211304 27560 211353 27588
rect 211304 27548 211310 27560
rect 211341 27557 211353 27560
rect 211387 27557 211399 27591
rect 211341 27551 211399 27557
rect 223669 27591 223727 27597
rect 223669 27557 223681 27591
rect 223715 27588 223727 27591
rect 223758 27588 223764 27600
rect 223715 27560 223764 27588
rect 223715 27557 223727 27560
rect 223669 27551 223727 27557
rect 223758 27548 223764 27560
rect 223816 27548 223822 27600
rect 238573 27591 238631 27597
rect 238573 27557 238585 27591
rect 238619 27588 238631 27591
rect 238662 27588 238668 27600
rect 238619 27560 238668 27588
rect 238619 27557 238631 27560
rect 238573 27551 238631 27557
rect 238662 27548 238668 27560
rect 238720 27548 238726 27600
rect 252738 27588 252744 27600
rect 252699 27560 252744 27588
rect 252738 27548 252744 27560
rect 252796 27548 252802 27600
rect 264974 27588 264980 27600
rect 264935 27560 264980 27588
rect 264974 27548 264980 27560
rect 265032 27548 265038 27600
rect 346210 27588 346216 27600
rect 346171 27560 346216 27588
rect 346210 27548 346216 27560
rect 346268 27548 346274 27600
rect 374270 27588 374276 27600
rect 374231 27560 374276 27588
rect 374270 27548 374276 27560
rect 374328 27548 374334 27600
rect 384577 27591 384635 27597
rect 384577 27557 384589 27591
rect 384623 27588 384635 27591
rect 384850 27588 384856 27600
rect 384623 27560 384856 27588
rect 384623 27557 384635 27560
rect 384577 27551 384635 27557
rect 384850 27548 384856 27560
rect 384908 27548 384914 27600
rect 379238 27520 379244 27532
rect 379199 27492 379244 27520
rect 379238 27480 379244 27492
rect 379296 27480 379302 27532
rect 245838 27248 245844 27260
rect 245799 27220 245844 27248
rect 245838 27208 245844 27220
rect 245896 27208 245902 27260
rect 151998 26256 152004 26308
rect 152056 26296 152062 26308
rect 152090 26296 152096 26308
rect 152056 26268 152096 26296
rect 152056 26256 152062 26268
rect 152090 26256 152096 26268
rect 152148 26256 152154 26308
rect 191926 26296 191932 26308
rect 191887 26268 191932 26296
rect 191926 26256 191932 26268
rect 191984 26256 191990 26308
rect 189166 26228 189172 26240
rect 189127 26200 189172 26228
rect 189166 26188 189172 26200
rect 189224 26188 189230 26240
rect 194686 26228 194692 26240
rect 194647 26200 194692 26228
rect 194686 26188 194692 26200
rect 194744 26188 194750 26240
rect 190638 22108 190644 22160
rect 190696 22108 190702 22160
rect 198274 22148 198280 22160
rect 198200 22120 198280 22148
rect 173986 22080 173992 22092
rect 173947 22052 173992 22080
rect 173986 22040 173992 22052
rect 174044 22040 174050 22092
rect 190656 22012 190684 22108
rect 198200 22092 198228 22120
rect 198274 22108 198280 22120
rect 198332 22108 198338 22160
rect 196158 22040 196164 22092
rect 196216 22080 196222 22092
rect 196342 22080 196348 22092
rect 196216 22052 196348 22080
rect 196216 22040 196222 22052
rect 196342 22040 196348 22052
rect 196400 22040 196406 22092
rect 198182 22040 198188 22092
rect 198240 22040 198246 22092
rect 346210 22080 346216 22092
rect 346171 22052 346216 22080
rect 346210 22040 346216 22052
rect 346268 22040 346274 22092
rect 379241 22083 379299 22089
rect 379241 22049 379253 22083
rect 379287 22080 379299 22083
rect 379330 22080 379336 22092
rect 379287 22052 379336 22080
rect 379287 22049 379299 22052
rect 379241 22043 379299 22049
rect 379330 22040 379336 22052
rect 379388 22040 379394 22092
rect 190730 22012 190736 22024
rect 190656 21984 190736 22012
rect 190730 21972 190736 21984
rect 190788 21972 190794 22024
rect 191742 21360 191748 21412
rect 191800 21400 191806 21412
rect 191929 21403 191987 21409
rect 191929 21400 191941 21403
rect 191800 21372 191941 21400
rect 191800 21360 191806 21372
rect 191929 21369 191941 21372
rect 191975 21369 191987 21403
rect 191929 21363 191987 21369
rect 218238 19388 218244 19440
rect 218296 19388 218302 19440
rect 219526 19388 219532 19440
rect 219584 19388 219590 19440
rect 211338 19360 211344 19372
rect 211299 19332 211344 19360
rect 211338 19320 211344 19332
rect 211396 19320 211402 19372
rect 218256 19304 218284 19388
rect 219544 19304 219572 19388
rect 229278 19320 229284 19372
rect 229336 19360 229342 19372
rect 229370 19360 229376 19372
rect 229336 19332 229376 19360
rect 229336 19320 229342 19332
rect 229370 19320 229376 19332
rect 229428 19320 229434 19372
rect 234706 19320 234712 19372
rect 234764 19360 234770 19372
rect 234798 19360 234804 19372
rect 234764 19332 234804 19360
rect 234764 19320 234770 19332
rect 234798 19320 234804 19332
rect 234856 19320 234862 19372
rect 236178 19320 236184 19372
rect 236236 19360 236242 19372
rect 236270 19360 236276 19372
rect 236236 19332 236276 19360
rect 236236 19320 236242 19332
rect 236270 19320 236276 19332
rect 236328 19320 236334 19372
rect 237466 19320 237472 19372
rect 237524 19360 237530 19372
rect 237558 19360 237564 19372
rect 237524 19332 237564 19360
rect 237524 19320 237530 19332
rect 237558 19320 237564 19332
rect 237616 19320 237622 19372
rect 239030 19320 239036 19372
rect 239088 19360 239094 19372
rect 239122 19360 239128 19372
rect 239088 19332 239128 19360
rect 239088 19320 239094 19332
rect 239122 19320 239128 19332
rect 239180 19320 239186 19372
rect 245841 19363 245899 19369
rect 245841 19329 245853 19363
rect 245887 19360 245899 19363
rect 245930 19360 245936 19372
rect 245887 19332 245936 19360
rect 245887 19329 245899 19332
rect 245841 19323 245899 19329
rect 245930 19320 245936 19332
rect 245988 19320 245994 19372
rect 270497 19363 270555 19369
rect 270497 19329 270509 19363
rect 270543 19360 270555 19363
rect 270586 19360 270592 19372
rect 270543 19332 270592 19360
rect 270543 19329 270555 19332
rect 270497 19323 270555 19329
rect 270586 19320 270592 19332
rect 270644 19320 270650 19372
rect 394050 19360 394056 19372
rect 394011 19332 394056 19360
rect 394050 19320 394056 19332
rect 394108 19320 394114 19372
rect 403710 19320 403716 19372
rect 403768 19360 403774 19372
rect 403802 19360 403808 19372
rect 403768 19332 403808 19360
rect 403768 19320 403774 19332
rect 403802 19320 403808 19332
rect 403860 19320 403866 19372
rect 218238 19252 218244 19304
rect 218296 19252 218302 19304
rect 219526 19252 219532 19304
rect 219584 19252 219590 19304
rect 247957 19295 248015 19301
rect 247957 19261 247969 19295
rect 248003 19292 248015 19295
rect 248322 19292 248328 19304
rect 248003 19264 248328 19292
rect 248003 19261 248015 19264
rect 247957 19255 248015 19261
rect 248322 19252 248328 19264
rect 248380 19252 248386 19304
rect 179506 18000 179512 18012
rect 179467 17972 179512 18000
rect 179506 17960 179512 17972
rect 179564 17960 179570 18012
rect 207109 18003 207167 18009
rect 207109 17969 207121 18003
rect 207155 18000 207167 18003
rect 207198 18000 207204 18012
rect 207155 17972 207204 18000
rect 207155 17969 207167 17972
rect 207109 17963 207167 17969
rect 207198 17960 207204 17972
rect 207256 17960 207262 18012
rect 252741 18003 252799 18009
rect 252741 17969 252753 18003
rect 252787 18000 252799 18003
rect 252830 18000 252836 18012
rect 252787 17972 252836 18000
rect 252787 17969 252799 17972
rect 252741 17963 252799 17969
rect 252830 17960 252836 17972
rect 252888 17960 252894 18012
rect 264977 18003 265035 18009
rect 264977 17969 264989 18003
rect 265023 18000 265035 18003
rect 265066 18000 265072 18012
rect 265023 17972 265072 18000
rect 265023 17969 265035 17972
rect 264977 17963 265035 17969
rect 265066 17960 265072 17972
rect 265124 17960 265130 18012
rect 374270 18000 374276 18012
rect 374231 17972 374276 18000
rect 374270 17960 374276 17972
rect 374328 17960 374334 18012
rect 384574 18000 384580 18012
rect 384535 17972 384580 18000
rect 384574 17960 384580 17972
rect 384632 17960 384638 18012
rect 154850 17932 154856 17944
rect 154811 17904 154856 17932
rect 154850 17892 154856 17904
rect 154908 17892 154914 17944
rect 338206 16804 338212 16856
rect 338264 16844 338270 16856
rect 342622 16844 342628 16856
rect 338264 16816 342628 16844
rect 338264 16804 338270 16816
rect 342622 16804 342628 16816
rect 342680 16804 342686 16856
rect 359918 16804 359924 16856
rect 359976 16844 359982 16856
rect 362218 16844 362224 16856
rect 359976 16816 362224 16844
rect 359976 16804 359982 16816
rect 362218 16804 362224 16816
rect 362276 16804 362282 16856
rect 379238 16804 379244 16856
rect 379296 16844 379302 16856
rect 379606 16844 379612 16856
rect 379296 16816 379612 16844
rect 379296 16804 379302 16816
rect 379606 16804 379612 16816
rect 379664 16804 379670 16856
rect 318794 16736 318800 16788
rect 318852 16776 318858 16788
rect 321554 16776 321560 16788
rect 318852 16748 321560 16776
rect 318852 16736 318858 16748
rect 321554 16736 321560 16748
rect 321612 16736 321618 16788
rect 398650 16736 398656 16788
rect 398708 16776 398714 16788
rect 400858 16776 400864 16788
rect 398708 16748 400864 16776
rect 398708 16736 398714 16748
rect 400858 16736 400864 16748
rect 400916 16736 400922 16788
rect 417970 16736 417976 16788
rect 418028 16776 418034 16788
rect 418246 16776 418252 16788
rect 418028 16748 418252 16776
rect 418028 16736 418034 16748
rect 418246 16736 418252 16748
rect 418304 16736 418310 16788
rect 173894 16668 173900 16720
rect 173952 16708 173958 16720
rect 183462 16708 183468 16720
rect 173952 16680 183468 16708
rect 173952 16668 173958 16680
rect 183462 16668 183468 16680
rect 183520 16668 183526 16720
rect 444374 16668 444380 16720
rect 444432 16708 444438 16720
rect 447226 16708 447232 16720
rect 444432 16680 447232 16708
rect 444432 16668 444438 16680
rect 447226 16668 447232 16680
rect 447284 16668 447290 16720
rect 476022 16668 476028 16720
rect 476080 16708 476086 16720
rect 482922 16708 482928 16720
rect 476080 16680 482928 16708
rect 476080 16668 476086 16680
rect 482922 16668 482928 16680
rect 482980 16668 482986 16720
rect 189166 16640 189172 16652
rect 189127 16612 189172 16640
rect 189166 16600 189172 16612
rect 189224 16600 189230 16652
rect 194686 16640 194692 16652
rect 194647 16612 194692 16640
rect 194686 16600 194692 16612
rect 194744 16600 194750 16652
rect 190454 13472 190460 13524
rect 190512 13512 190518 13524
rect 190730 13512 190736 13524
rect 190512 13484 190736 13512
rect 190512 13472 190518 13484
rect 190730 13472 190736 13484
rect 190788 13472 190794 13524
rect 374181 12563 374239 12569
rect 374181 12529 374193 12563
rect 374227 12560 374239 12563
rect 374270 12560 374276 12572
rect 374227 12532 374276 12560
rect 374227 12529 374239 12532
rect 374181 12523 374239 12529
rect 374270 12520 374276 12532
rect 374328 12520 374334 12572
rect 168558 12492 168564 12504
rect 168484 12464 168564 12492
rect 168484 12436 168512 12464
rect 168558 12452 168564 12464
rect 168616 12452 168622 12504
rect 216858 12492 216864 12504
rect 216784 12464 216864 12492
rect 216784 12436 216812 12464
rect 216858 12452 216864 12464
rect 216916 12452 216922 12504
rect 424778 12452 424784 12504
rect 424836 12492 424842 12504
rect 424962 12492 424968 12504
rect 424836 12464 424968 12492
rect 424836 12452 424842 12464
rect 424962 12452 424968 12464
rect 425020 12452 425026 12504
rect 154850 12424 154856 12436
rect 154811 12396 154856 12424
rect 154850 12384 154856 12396
rect 154908 12384 154914 12436
rect 168466 12384 168472 12436
rect 168524 12384 168530 12436
rect 216766 12384 216772 12436
rect 216824 12384 216830 12436
rect 356330 12384 356336 12436
rect 356388 12384 356394 12436
rect 357434 12384 357440 12436
rect 357492 12424 357498 12436
rect 358538 12424 358544 12436
rect 357492 12396 358544 12424
rect 357492 12384 357498 12396
rect 358538 12384 358544 12396
rect 358596 12384 358602 12436
rect 375558 12384 375564 12436
rect 375616 12424 375622 12436
rect 376386 12424 376392 12436
rect 375616 12396 376392 12424
rect 375616 12384 375622 12396
rect 376386 12384 376392 12396
rect 376444 12384 376450 12436
rect 356348 12356 356376 12384
rect 357342 12356 357348 12368
rect 356348 12328 357348 12356
rect 357342 12316 357348 12328
rect 357400 12316 357406 12368
rect 169846 9664 169852 9716
rect 169904 9704 169910 9716
rect 170122 9704 170128 9716
rect 169904 9676 170128 9704
rect 169904 9664 169910 9676
rect 170122 9664 170128 9676
rect 170180 9664 170186 9716
rect 191926 9704 191932 9716
rect 191887 9676 191932 9704
rect 191926 9664 191932 9676
rect 191984 9664 191990 9716
rect 223666 9704 223672 9716
rect 223627 9676 223672 9704
rect 223666 9664 223672 9676
rect 223724 9664 223730 9716
rect 238570 9704 238576 9716
rect 238531 9676 238576 9704
rect 238570 9664 238576 9676
rect 238628 9664 238634 9716
rect 247954 9704 247960 9716
rect 247915 9676 247960 9704
rect 247954 9664 247960 9676
rect 248012 9664 248018 9716
rect 270497 9707 270555 9713
rect 270497 9673 270509 9707
rect 270543 9704 270555 9707
rect 270586 9704 270592 9716
rect 270543 9676 270592 9704
rect 270543 9673 270555 9676
rect 270497 9667 270555 9673
rect 270586 9664 270592 9676
rect 270644 9664 270650 9716
rect 309410 9664 309416 9716
rect 309468 9704 309474 9716
rect 309778 9704 309784 9716
rect 309468 9676 309784 9704
rect 309468 9664 309474 9676
rect 309778 9664 309784 9676
rect 309836 9664 309842 9716
rect 374178 9704 374184 9716
rect 374139 9676 374184 9704
rect 374178 9664 374184 9676
rect 374236 9664 374242 9716
rect 384574 9664 384580 9716
rect 384632 9704 384638 9716
rect 384850 9704 384856 9716
rect 384632 9676 384856 9704
rect 384632 9664 384638 9676
rect 384850 9664 384856 9676
rect 384908 9664 384914 9716
rect 109954 9596 109960 9648
rect 110012 9636 110018 9648
rect 205818 9636 205824 9648
rect 110012 9608 205824 9636
rect 110012 9596 110018 9608
rect 205818 9596 205824 9608
rect 205876 9596 205882 9648
rect 106366 9528 106372 9580
rect 106424 9568 106430 9580
rect 204346 9568 204352 9580
rect 106424 9540 204352 9568
rect 106424 9528 106430 9540
rect 204346 9528 204352 9540
rect 204404 9528 204410 9580
rect 102778 9460 102784 9512
rect 102836 9500 102842 9512
rect 201586 9500 201592 9512
rect 102836 9472 201592 9500
rect 102836 9460 102842 9472
rect 201586 9460 201592 9472
rect 201644 9460 201650 9512
rect 383562 9460 383568 9512
rect 383620 9500 383626 9512
rect 452470 9500 452476 9512
rect 383620 9472 452476 9500
rect 383620 9460 383626 9472
rect 452470 9460 452476 9472
rect 452528 9460 452534 9512
rect 95694 9392 95700 9444
rect 95752 9432 95758 9444
rect 198826 9432 198832 9444
rect 95752 9404 198832 9432
rect 95752 9392 95758 9404
rect 198826 9392 198832 9404
rect 198884 9392 198890 9444
rect 380710 9392 380716 9444
rect 380768 9432 380774 9444
rect 448974 9432 448980 9444
rect 380768 9404 448980 9432
rect 380768 9392 380774 9404
rect 448974 9392 448980 9404
rect 449032 9392 449038 9444
rect 92106 9324 92112 9376
rect 92164 9364 92170 9376
rect 196066 9364 196072 9376
rect 92164 9336 196072 9364
rect 92164 9324 92170 9336
rect 196066 9324 196072 9336
rect 196124 9324 196130 9376
rect 384850 9324 384856 9376
rect 384908 9364 384914 9376
rect 456058 9364 456064 9376
rect 384908 9336 456064 9364
rect 384908 9324 384914 9336
rect 456058 9324 456064 9336
rect 456116 9324 456122 9376
rect 88518 9256 88524 9308
rect 88576 9296 88582 9308
rect 194778 9296 194784 9308
rect 88576 9268 194784 9296
rect 88576 9256 88582 9268
rect 194778 9256 194784 9268
rect 194836 9256 194842 9308
rect 386230 9256 386236 9308
rect 386288 9296 386294 9308
rect 459646 9296 459652 9308
rect 386288 9268 459652 9296
rect 386288 9256 386294 9268
rect 459646 9256 459652 9268
rect 459704 9256 459710 9308
rect 84930 9188 84936 9240
rect 84988 9228 84994 9240
rect 193306 9228 193312 9240
rect 84988 9200 193312 9228
rect 84988 9188 84994 9200
rect 193306 9188 193312 9200
rect 193364 9188 193370 9240
rect 388990 9188 388996 9240
rect 389048 9228 389054 9240
rect 463234 9228 463240 9240
rect 389048 9200 463240 9228
rect 389048 9188 389054 9200
rect 463234 9188 463240 9200
rect 463292 9188 463298 9240
rect 81434 9120 81440 9172
rect 81492 9160 81498 9172
rect 190546 9160 190552 9172
rect 81492 9132 190552 9160
rect 81492 9120 81498 9132
rect 190546 9120 190552 9132
rect 190604 9120 190610 9172
rect 391750 9120 391756 9172
rect 391808 9160 391814 9172
rect 470318 9160 470324 9172
rect 391808 9132 470324 9160
rect 391808 9120 391814 9132
rect 470318 9120 470324 9132
rect 470376 9120 470382 9172
rect 77846 9052 77852 9104
rect 77904 9092 77910 9104
rect 189166 9092 189172 9104
rect 77904 9064 189172 9092
rect 77904 9052 77910 9064
rect 189166 9052 189172 9064
rect 189224 9052 189230 9104
rect 445570 9052 445576 9104
rect 445628 9092 445634 9104
rect 573818 9092 573824 9104
rect 445628 9064 573824 9092
rect 445628 9052 445634 9064
rect 573818 9052 573824 9064
rect 573876 9052 573882 9104
rect 74258 8984 74264 9036
rect 74316 9024 74322 9036
rect 187786 9024 187792 9036
rect 74316 8996 187792 9024
rect 74316 8984 74322 8996
rect 187786 8984 187792 8996
rect 187844 8984 187850 9036
rect 446950 8984 446956 9036
rect 447008 9024 447014 9036
rect 577406 9024 577412 9036
rect 447008 8996 577412 9024
rect 447008 8984 447014 8996
rect 577406 8984 577412 8996
rect 577464 8984 577470 9036
rect 31478 8916 31484 8968
rect 31536 8956 31542 8968
rect 165706 8956 165712 8968
rect 31536 8928 165712 8956
rect 31536 8916 31542 8928
rect 165706 8916 165712 8928
rect 165764 8916 165770 8968
rect 448330 8916 448336 8968
rect 448388 8956 448394 8968
rect 580994 8956 581000 8968
rect 448388 8928 581000 8956
rect 448388 8916 448394 8928
rect 580994 8916 581000 8928
rect 581052 8916 581058 8968
rect 117130 8848 117136 8900
rect 117188 8888 117194 8900
rect 209866 8888 209872 8900
rect 117188 8860 209872 8888
rect 117188 8848 117194 8860
rect 209866 8848 209872 8860
rect 209924 8848 209930 8900
rect 120626 8780 120632 8832
rect 120684 8820 120690 8832
rect 211338 8820 211344 8832
rect 120684 8792 211344 8820
rect 120684 8780 120690 8792
rect 211338 8780 211344 8792
rect 211396 8780 211402 8832
rect 124214 8712 124220 8764
rect 124272 8752 124278 8764
rect 212626 8752 212632 8764
rect 124272 8724 212632 8752
rect 124272 8712 124278 8724
rect 212626 8712 212632 8724
rect 212684 8712 212690 8764
rect 131390 8644 131396 8696
rect 131448 8684 131454 8696
rect 216766 8684 216772 8696
rect 131448 8656 216772 8684
rect 131448 8644 131454 8656
rect 216766 8644 216772 8656
rect 216824 8644 216830 8696
rect 134886 8576 134892 8628
rect 134944 8616 134950 8628
rect 218238 8616 218244 8628
rect 134944 8588 218244 8616
rect 134944 8576 134950 8588
rect 218238 8576 218244 8588
rect 218296 8576 218302 8628
rect 138474 8508 138480 8560
rect 138532 8548 138538 8560
rect 220906 8548 220912 8560
rect 138532 8520 220912 8548
rect 138532 8508 138538 8520
rect 220906 8508 220912 8520
rect 220964 8508 220970 8560
rect 142062 8440 142068 8492
rect 142120 8480 142126 8492
rect 222378 8480 222384 8492
rect 142120 8452 222384 8480
rect 142120 8440 142126 8452
rect 222378 8440 222384 8452
rect 222436 8440 222442 8492
rect 145650 8372 145656 8424
rect 145708 8412 145714 8424
rect 223666 8412 223672 8424
rect 145708 8384 223672 8412
rect 145708 8372 145714 8384
rect 223666 8372 223672 8384
rect 223724 8372 223730 8424
rect 156322 8304 156328 8356
rect 156380 8344 156386 8356
rect 229278 8344 229284 8356
rect 156380 8316 229284 8344
rect 156380 8304 156386 8316
rect 229278 8304 229284 8316
rect 229336 8304 229342 8356
rect 119430 8236 119436 8288
rect 119488 8276 119494 8288
rect 211154 8276 211160 8288
rect 119488 8248 211160 8276
rect 119488 8236 119494 8248
rect 211154 8236 211160 8248
rect 211212 8236 211218 8288
rect 422110 8236 422116 8288
rect 422168 8276 422174 8288
rect 527450 8276 527456 8288
rect 422168 8248 527456 8276
rect 422168 8236 422174 8248
rect 527450 8236 527456 8248
rect 527508 8236 527514 8288
rect 2774 8168 2780 8220
rect 2832 8208 2838 8220
rect 4798 8208 4804 8220
rect 2832 8180 4804 8208
rect 2832 8168 2838 8180
rect 4798 8168 4804 8180
rect 4856 8168 4862 8220
rect 115934 8168 115940 8220
rect 115992 8208 115998 8220
rect 208578 8208 208584 8220
rect 115992 8180 208584 8208
rect 115992 8168 115998 8180
rect 208578 8168 208584 8180
rect 208636 8168 208642 8220
rect 423398 8168 423404 8220
rect 423456 8208 423462 8220
rect 531038 8208 531044 8220
rect 423456 8180 531044 8208
rect 423456 8168 423462 8180
rect 531038 8168 531044 8180
rect 531096 8168 531102 8220
rect 112346 8100 112352 8152
rect 112404 8140 112410 8152
rect 207198 8140 207204 8152
rect 112404 8112 207204 8140
rect 112404 8100 112410 8112
rect 207198 8100 207204 8112
rect 207256 8100 207262 8152
rect 420822 8100 420828 8152
rect 420880 8140 420886 8152
rect 423309 8143 423367 8149
rect 423309 8140 423321 8143
rect 420880 8112 423321 8140
rect 420880 8100 420886 8112
rect 423309 8109 423321 8112
rect 423355 8109 423367 8143
rect 423309 8103 423367 8109
rect 424870 8100 424876 8152
rect 424928 8140 424934 8152
rect 534534 8140 534540 8152
rect 424928 8112 534540 8140
rect 424928 8100 424934 8112
rect 534534 8100 534540 8112
rect 534592 8100 534598 8152
rect 108758 8032 108764 8084
rect 108816 8072 108822 8084
rect 205634 8072 205640 8084
rect 108816 8044 205640 8072
rect 108816 8032 108822 8044
rect 205634 8032 205640 8044
rect 205692 8032 205698 8084
rect 426250 8032 426256 8084
rect 426308 8072 426314 8084
rect 538122 8072 538128 8084
rect 426308 8044 538128 8072
rect 426308 8032 426314 8044
rect 538122 8032 538128 8044
rect 538180 8032 538186 8084
rect 105170 7964 105176 8016
rect 105228 8004 105234 8016
rect 202966 8004 202972 8016
rect 105228 7976 202972 8004
rect 105228 7964 105234 7976
rect 202966 7964 202972 7976
rect 203024 7964 203030 8016
rect 429102 7964 429108 8016
rect 429160 8004 429166 8016
rect 541710 8004 541716 8016
rect 429160 7976 541716 8004
rect 429160 7964 429166 7976
rect 541710 7964 541716 7976
rect 541768 7964 541774 8016
rect 101582 7896 101588 7948
rect 101640 7936 101646 7948
rect 201678 7936 201684 7948
rect 101640 7908 201684 7936
rect 101640 7896 101646 7908
rect 201678 7896 201684 7908
rect 201736 7896 201742 7948
rect 430390 7896 430396 7948
rect 430448 7936 430454 7948
rect 545298 7936 545304 7948
rect 430448 7908 545304 7936
rect 430448 7896 430454 7908
rect 545298 7896 545304 7908
rect 545356 7896 545362 7948
rect 98086 7828 98092 7880
rect 98144 7868 98150 7880
rect 200206 7868 200212 7880
rect 98144 7840 200212 7868
rect 98144 7828 98150 7840
rect 200206 7828 200212 7840
rect 200264 7828 200270 7880
rect 431678 7828 431684 7880
rect 431736 7868 431742 7880
rect 548886 7868 548892 7880
rect 431736 7840 548892 7868
rect 431736 7828 431742 7840
rect 548886 7828 548892 7840
rect 548944 7828 548950 7880
rect 94498 7760 94504 7812
rect 94556 7800 94562 7812
rect 197446 7800 197452 7812
rect 94556 7772 197452 7800
rect 94556 7760 94562 7772
rect 197446 7760 197452 7772
rect 197504 7760 197510 7812
rect 434530 7760 434536 7812
rect 434588 7800 434594 7812
rect 552382 7800 552388 7812
rect 434588 7772 552388 7800
rect 434588 7760 434594 7772
rect 552382 7760 552388 7772
rect 552440 7760 552446 7812
rect 90910 7692 90916 7744
rect 90968 7732 90974 7744
rect 196342 7732 196348 7744
rect 90968 7704 196348 7732
rect 90968 7692 90974 7704
rect 196342 7692 196348 7704
rect 196400 7692 196406 7744
rect 435910 7692 435916 7744
rect 435968 7732 435974 7744
rect 555970 7732 555976 7744
rect 435968 7704 555976 7732
rect 435968 7692 435974 7704
rect 555970 7692 555976 7704
rect 556028 7692 556034 7744
rect 87322 7624 87328 7676
rect 87380 7664 87386 7676
rect 194594 7664 194600 7676
rect 87380 7636 194600 7664
rect 87380 7624 87386 7636
rect 194594 7624 194600 7636
rect 194652 7624 194658 7676
rect 369670 7624 369676 7676
rect 369728 7664 369734 7676
rect 427538 7664 427544 7676
rect 369728 7636 427544 7664
rect 369728 7624 369734 7636
rect 427538 7624 427544 7636
rect 427596 7624 427602 7676
rect 437290 7624 437296 7676
rect 437348 7664 437354 7676
rect 559558 7664 559564 7676
rect 437348 7636 559564 7664
rect 437348 7624 437354 7636
rect 559558 7624 559564 7636
rect 559616 7624 559622 7676
rect 23106 7556 23112 7608
rect 23164 7596 23170 7608
rect 161566 7596 161572 7608
rect 23164 7568 161572 7596
rect 23164 7556 23170 7568
rect 161566 7556 161572 7568
rect 161624 7556 161630 7608
rect 162302 7556 162308 7608
rect 162360 7596 162366 7608
rect 233418 7596 233424 7608
rect 162360 7568 233424 7596
rect 162360 7556 162366 7568
rect 233418 7556 233424 7568
rect 233476 7556 233482 7608
rect 434530 7596 434536 7608
rect 376588 7568 434536 7596
rect 123018 7488 123024 7540
rect 123076 7528 123082 7540
rect 212718 7528 212724 7540
rect 123076 7500 212724 7528
rect 123076 7488 123082 7500
rect 212718 7488 212724 7500
rect 212776 7488 212782 7540
rect 127802 7420 127808 7472
rect 127860 7460 127866 7472
rect 215386 7460 215392 7472
rect 127860 7432 215392 7460
rect 127860 7420 127866 7432
rect 215386 7420 215392 7432
rect 215444 7420 215450 7472
rect 373718 7420 373724 7472
rect 373776 7460 373782 7472
rect 376588 7460 376616 7568
rect 434530 7556 434536 7568
rect 434588 7556 434594 7608
rect 441430 7556 441436 7608
rect 441488 7596 441494 7608
rect 566734 7596 566740 7608
rect 441488 7568 566740 7596
rect 441488 7556 441494 7568
rect 566734 7556 566740 7568
rect 566792 7556 566798 7608
rect 419350 7488 419356 7540
rect 419408 7528 419414 7540
rect 523862 7528 523868 7540
rect 419408 7500 523868 7528
rect 419408 7488 419414 7500
rect 523862 7488 523868 7500
rect 523920 7488 523926 7540
rect 373776 7432 376616 7460
rect 373776 7420 373782 7432
rect 411070 7420 411076 7472
rect 411128 7460 411134 7472
rect 508406 7460 508412 7472
rect 411128 7432 508412 7460
rect 411128 7420 411134 7432
rect 508406 7420 508412 7432
rect 508464 7420 508470 7472
rect 126606 7352 126612 7404
rect 126664 7392 126670 7404
rect 214098 7392 214104 7404
rect 126664 7364 214104 7392
rect 126664 7352 126670 7364
rect 214098 7352 214104 7364
rect 214156 7352 214162 7404
rect 409782 7352 409788 7404
rect 409840 7392 409846 7404
rect 504818 7392 504824 7404
rect 409840 7364 504824 7392
rect 409840 7352 409846 7364
rect 504818 7352 504824 7364
rect 504876 7352 504882 7404
rect 130194 7284 130200 7336
rect 130252 7324 130258 7336
rect 216674 7324 216680 7336
rect 130252 7296 216680 7324
rect 130252 7284 130258 7296
rect 216674 7284 216680 7296
rect 216732 7284 216738 7336
rect 408310 7284 408316 7336
rect 408368 7324 408374 7336
rect 501230 7324 501236 7336
rect 408368 7296 501236 7324
rect 408368 7284 408374 7296
rect 501230 7284 501236 7296
rect 501288 7284 501294 7336
rect 133782 7216 133788 7268
rect 133840 7256 133846 7268
rect 218146 7256 218152 7268
rect 133840 7228 218152 7256
rect 133840 7216 133846 7228
rect 218146 7216 218152 7228
rect 218204 7216 218210 7268
rect 405550 7216 405556 7268
rect 405608 7256 405614 7268
rect 497734 7256 497740 7268
rect 405608 7228 497740 7256
rect 405608 7216 405614 7228
rect 497734 7216 497740 7228
rect 497792 7216 497798 7268
rect 137278 7148 137284 7200
rect 137336 7188 137342 7200
rect 219526 7188 219532 7200
rect 137336 7160 219532 7188
rect 137336 7148 137342 7160
rect 219526 7148 219532 7160
rect 219584 7148 219590 7200
rect 404262 7148 404268 7200
rect 404320 7188 404326 7200
rect 494146 7188 494152 7200
rect 404320 7160 494152 7188
rect 404320 7148 404326 7160
rect 494146 7148 494152 7160
rect 494204 7148 494210 7200
rect 140866 7080 140872 7132
rect 140924 7120 140930 7132
rect 222286 7120 222292 7132
rect 140924 7092 222292 7120
rect 140924 7080 140930 7092
rect 222286 7080 222292 7092
rect 222344 7080 222350 7132
rect 402790 7080 402796 7132
rect 402848 7120 402854 7132
rect 490558 7120 490564 7132
rect 402848 7092 490564 7120
rect 402848 7080 402854 7092
rect 490558 7080 490564 7092
rect 490616 7080 490622 7132
rect 144454 7012 144460 7064
rect 144512 7052 144518 7064
rect 223574 7052 223580 7064
rect 144512 7024 223580 7052
rect 144512 7012 144518 7024
rect 223574 7012 223580 7024
rect 223632 7012 223638 7064
rect 400030 7012 400036 7064
rect 400088 7052 400094 7064
rect 486970 7052 486976 7064
rect 400088 7024 486976 7052
rect 400088 7012 400094 7024
rect 486970 7012 486976 7024
rect 487028 7012 487034 7064
rect 148042 6944 148048 6996
rect 148100 6984 148106 6996
rect 225138 6984 225144 6996
rect 148100 6956 225144 6984
rect 148100 6944 148106 6956
rect 225138 6944 225144 6956
rect 225196 6944 225202 6996
rect 258166 6984 258172 6996
rect 258092 6956 258172 6984
rect 258092 6928 258120 6956
rect 258166 6944 258172 6956
rect 258224 6944 258230 6996
rect 379238 6944 379244 6996
rect 379296 6984 379302 6996
rect 445386 6984 445392 6996
rect 379296 6956 445392 6984
rect 379296 6944 379302 6956
rect 445386 6944 445392 6956
rect 445444 6944 445450 6996
rect 150802 6876 150808 6928
rect 150860 6916 150866 6928
rect 150894 6916 150900 6928
rect 150860 6888 150900 6916
rect 150860 6876 150866 6888
rect 150894 6876 150900 6888
rect 150952 6876 150958 6928
rect 258074 6876 258080 6928
rect 258132 6876 258138 6928
rect 67174 6808 67180 6860
rect 67232 6848 67238 6860
rect 183738 6848 183744 6860
rect 67232 6820 183744 6848
rect 67232 6808 67238 6820
rect 183738 6808 183744 6820
rect 183796 6808 183802 6860
rect 398742 6808 398748 6860
rect 398800 6848 398806 6860
rect 483474 6848 483480 6860
rect 398800 6820 483480 6848
rect 398800 6808 398806 6820
rect 483474 6808 483480 6820
rect 483532 6808 483538 6860
rect 63586 6740 63592 6792
rect 63644 6780 63650 6792
rect 182266 6780 182272 6792
rect 63644 6752 182272 6780
rect 63644 6740 63650 6752
rect 182266 6740 182272 6752
rect 182324 6740 182330 6792
rect 401502 6740 401508 6792
rect 401560 6780 401566 6792
rect 488166 6780 488172 6792
rect 401560 6752 488172 6780
rect 401560 6740 401566 6752
rect 488166 6740 488172 6752
rect 488224 6740 488230 6792
rect 59998 6672 60004 6724
rect 60056 6712 60062 6724
rect 180886 6712 180892 6724
rect 60056 6684 180892 6712
rect 60056 6672 60062 6684
rect 180886 6672 180892 6684
rect 180944 6672 180950 6724
rect 402882 6672 402888 6724
rect 402940 6712 402946 6724
rect 491754 6712 491760 6724
rect 402940 6684 491760 6712
rect 402940 6672 402946 6684
rect 491754 6672 491760 6684
rect 491812 6672 491818 6724
rect 56410 6604 56416 6656
rect 56468 6644 56474 6656
rect 178218 6644 178224 6656
rect 56468 6616 178224 6644
rect 56468 6604 56474 6616
rect 178218 6604 178224 6616
rect 178276 6604 178282 6656
rect 405642 6604 405648 6656
rect 405700 6644 405706 6656
rect 495342 6644 495348 6656
rect 405700 6616 495348 6644
rect 405700 6604 405706 6616
rect 495342 6604 495348 6616
rect 495400 6604 495406 6656
rect 52822 6536 52828 6588
rect 52880 6576 52886 6588
rect 176746 6576 176752 6588
rect 52880 6548 176752 6576
rect 52880 6536 52886 6548
rect 176746 6536 176752 6548
rect 176804 6536 176810 6588
rect 178954 6536 178960 6588
rect 179012 6576 179018 6588
rect 241606 6576 241612 6588
rect 179012 6548 241612 6576
rect 179012 6536 179018 6548
rect 241606 6536 241612 6548
rect 241664 6536 241670 6588
rect 407022 6536 407028 6588
rect 407080 6576 407086 6588
rect 498930 6576 498936 6588
rect 407080 6548 498936 6576
rect 407080 6536 407086 6548
rect 498930 6536 498936 6548
rect 498988 6536 498994 6588
rect 49326 6468 49332 6520
rect 49384 6508 49390 6520
rect 175274 6508 175280 6520
rect 49384 6480 175280 6508
rect 49384 6468 49390 6480
rect 175274 6468 175280 6480
rect 175332 6468 175338 6520
rect 175366 6468 175372 6520
rect 175424 6508 175430 6520
rect 239030 6508 239036 6520
rect 175424 6480 239036 6508
rect 175424 6468 175430 6480
rect 239030 6468 239036 6480
rect 239088 6468 239094 6520
rect 408402 6468 408408 6520
rect 408460 6508 408466 6520
rect 502426 6508 502432 6520
rect 408460 6480 502432 6508
rect 408460 6468 408466 6480
rect 502426 6468 502432 6480
rect 502484 6468 502490 6520
rect 40954 6400 40960 6452
rect 41012 6440 41018 6452
rect 169846 6440 169852 6452
rect 41012 6412 169852 6440
rect 41012 6400 41018 6412
rect 169846 6400 169852 6412
rect 169904 6400 169910 6452
rect 171778 6400 171784 6452
rect 171836 6440 171842 6452
rect 237558 6440 237564 6452
rect 171836 6412 237564 6440
rect 171836 6400 171842 6412
rect 237558 6400 237564 6412
rect 237616 6400 237622 6452
rect 353110 6400 353116 6452
rect 353168 6440 353174 6452
rect 395338 6440 395344 6452
rect 353168 6412 395344 6440
rect 353168 6400 353174 6412
rect 395338 6400 395344 6412
rect 395396 6400 395402 6452
rect 411162 6400 411168 6452
rect 411220 6440 411226 6452
rect 506014 6440 506020 6452
rect 411220 6412 506020 6440
rect 411220 6400 411226 6412
rect 506014 6400 506020 6412
rect 506072 6400 506078 6452
rect 18322 6332 18328 6384
rect 18380 6372 18386 6384
rect 158898 6372 158904 6384
rect 18380 6344 158904 6372
rect 18380 6332 18386 6344
rect 158898 6332 158904 6344
rect 158956 6332 158962 6384
rect 161106 6332 161112 6384
rect 161164 6372 161170 6384
rect 231854 6372 231860 6384
rect 161164 6344 231860 6372
rect 161164 6332 161170 6344
rect 231854 6332 231860 6344
rect 231912 6332 231918 6384
rect 355870 6332 355876 6384
rect 355928 6372 355934 6384
rect 399018 6372 399024 6384
rect 355928 6344 399024 6372
rect 355928 6332 355934 6344
rect 399018 6332 399024 6344
rect 399076 6332 399082 6384
rect 412542 6332 412548 6384
rect 412600 6372 412606 6384
rect 509602 6372 509608 6384
rect 412600 6344 509608 6372
rect 412600 6332 412606 6344
rect 509602 6332 509608 6344
rect 509660 6332 509666 6384
rect 13630 6264 13636 6316
rect 13688 6304 13694 6316
rect 156138 6304 156144 6316
rect 13688 6276 156144 6304
rect 13688 6264 13694 6276
rect 156138 6264 156144 6276
rect 156196 6264 156202 6316
rect 159910 6264 159916 6316
rect 159968 6304 159974 6316
rect 231946 6304 231952 6316
rect 159968 6276 231952 6304
rect 159968 6264 159974 6276
rect 231946 6264 231952 6276
rect 232004 6264 232010 6316
rect 358630 6264 358636 6316
rect 358688 6304 358694 6316
rect 406102 6304 406108 6316
rect 358688 6276 406108 6304
rect 358688 6264 358694 6276
rect 406102 6264 406108 6276
rect 406160 6264 406166 6316
rect 413830 6264 413836 6316
rect 413888 6304 413894 6316
rect 513190 6304 513196 6316
rect 413888 6276 513196 6304
rect 413888 6264 413894 6276
rect 513190 6264 513196 6276
rect 513248 6264 513254 6316
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 153378 6236 153384 6248
rect 8904 6208 153384 6236
rect 8904 6196 8910 6208
rect 153378 6196 153384 6208
rect 153436 6196 153442 6248
rect 157518 6196 157524 6248
rect 157576 6236 157582 6248
rect 230566 6236 230572 6248
rect 157576 6208 230572 6236
rect 157576 6196 157582 6208
rect 230566 6196 230572 6208
rect 230624 6196 230630 6248
rect 362678 6196 362684 6248
rect 362736 6236 362742 6248
rect 413278 6236 413284 6248
rect 362736 6208 413284 6236
rect 362736 6196 362742 6208
rect 413278 6196 413284 6208
rect 413336 6196 413342 6248
rect 416498 6196 416504 6248
rect 416556 6236 416562 6248
rect 516778 6236 516784 6248
rect 416556 6208 516784 6236
rect 416556 6196 416562 6208
rect 516778 6196 516784 6208
rect 516836 6196 516842 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 151906 6168 151912 6180
rect 4120 6140 151912 6168
rect 4120 6128 4126 6140
rect 151906 6128 151912 6140
rect 151964 6128 151970 6180
rect 153930 6128 153936 6180
rect 153988 6168 153994 6180
rect 227806 6168 227812 6180
rect 153988 6140 227812 6168
rect 153988 6128 153994 6140
rect 227806 6128 227812 6140
rect 227864 6128 227870 6180
rect 364150 6128 364156 6180
rect 364208 6168 364214 6180
rect 416866 6168 416872 6180
rect 364208 6140 416872 6168
rect 364208 6128 364214 6140
rect 416866 6128 416872 6140
rect 416924 6128 416930 6180
rect 418062 6128 418068 6180
rect 418120 6168 418126 6180
rect 520274 6168 520280 6180
rect 418120 6140 520280 6168
rect 418120 6128 418126 6140
rect 520274 6128 520280 6140
rect 520332 6128 520338 6180
rect 128998 6060 129004 6112
rect 129056 6100 129062 6112
rect 215294 6100 215300 6112
rect 129056 6072 215300 6100
rect 129056 6060 129062 6072
rect 215294 6060 215300 6072
rect 215352 6060 215358 6112
rect 400122 6060 400128 6112
rect 400180 6100 400186 6112
rect 484578 6100 484584 6112
rect 400180 6072 484584 6100
rect 400180 6060 400186 6072
rect 484578 6060 484584 6072
rect 484636 6060 484642 6112
rect 132586 5992 132592 6044
rect 132644 6032 132650 6044
rect 218054 6032 218060 6044
rect 132644 6004 218060 6032
rect 132644 5992 132650 6004
rect 218054 5992 218060 6004
rect 218112 5992 218118 6044
rect 397362 5992 397368 6044
rect 397420 6032 397426 6044
rect 479886 6032 479892 6044
rect 397420 6004 479892 6032
rect 397420 5992 397426 6004
rect 479886 5992 479892 6004
rect 479944 5992 479950 6044
rect 136082 5924 136088 5976
rect 136140 5964 136146 5976
rect 219434 5964 219440 5976
rect 136140 5936 219440 5964
rect 136140 5924 136146 5936
rect 219434 5924 219440 5936
rect 219492 5924 219498 5976
rect 394602 5924 394608 5976
rect 394660 5964 394666 5976
rect 476298 5964 476304 5976
rect 394660 5936 476304 5964
rect 394660 5924 394666 5936
rect 476298 5924 476304 5936
rect 476356 5924 476362 5976
rect 139670 5856 139676 5908
rect 139728 5896 139734 5908
rect 220814 5896 220820 5908
rect 139728 5868 220820 5896
rect 139728 5856 139734 5868
rect 220814 5856 220820 5868
rect 220872 5856 220878 5908
rect 393222 5856 393228 5908
rect 393280 5896 393286 5908
rect 472710 5896 472716 5908
rect 393280 5868 472716 5896
rect 393280 5856 393286 5868
rect 472710 5856 472716 5868
rect 472768 5856 472774 5908
rect 143258 5788 143264 5840
rect 143316 5828 143322 5840
rect 222194 5828 222200 5840
rect 143316 5800 222200 5828
rect 143316 5788 143322 5800
rect 222194 5788 222200 5800
rect 222252 5788 222258 5840
rect 391842 5788 391848 5840
rect 391900 5828 391906 5840
rect 469122 5828 469128 5840
rect 391900 5800 469128 5828
rect 391900 5788 391906 5800
rect 469122 5788 469128 5800
rect 469180 5788 469186 5840
rect 146846 5720 146852 5772
rect 146904 5760 146910 5772
rect 224954 5760 224960 5772
rect 146904 5732 224960 5760
rect 146904 5720 146910 5732
rect 224954 5720 224960 5732
rect 225012 5720 225018 5772
rect 389082 5720 389088 5772
rect 389140 5760 389146 5772
rect 465626 5760 465632 5772
rect 389140 5732 465632 5760
rect 389140 5720 389146 5732
rect 465626 5720 465632 5732
rect 465684 5720 465690 5772
rect 113177 5695 113235 5701
rect 113177 5661 113189 5695
rect 113223 5692 113235 5695
rect 122745 5695 122803 5701
rect 122745 5692 122757 5695
rect 113223 5664 122757 5692
rect 113223 5661 113235 5664
rect 113177 5655 113235 5661
rect 122745 5661 122757 5664
rect 122791 5661 122803 5695
rect 122745 5655 122803 5661
rect 132497 5695 132555 5701
rect 132497 5661 132509 5695
rect 132543 5692 132555 5695
rect 142065 5695 142123 5701
rect 142065 5692 142077 5695
rect 132543 5664 142077 5692
rect 132543 5661 132555 5664
rect 132497 5655 132555 5661
rect 142065 5661 142077 5664
rect 142111 5661 142123 5695
rect 142065 5655 142123 5661
rect 150434 5652 150440 5704
rect 150492 5692 150498 5704
rect 226518 5692 226524 5704
rect 150492 5664 226524 5692
rect 150492 5652 150498 5664
rect 226518 5652 226524 5664
rect 226576 5652 226582 5704
rect 387702 5652 387708 5704
rect 387760 5692 387766 5704
rect 462038 5692 462044 5704
rect 387760 5664 462044 5692
rect 387760 5652 387766 5664
rect 462038 5652 462044 5664
rect 462096 5652 462102 5704
rect 99282 5584 99288 5636
rect 99340 5624 99346 5636
rect 163498 5624 163504 5636
rect 99340 5596 163504 5624
rect 99340 5584 99346 5596
rect 163498 5584 163504 5596
rect 163556 5584 163562 5636
rect 164694 5584 164700 5636
rect 164752 5624 164758 5636
rect 233326 5624 233332 5636
rect 164752 5596 233332 5624
rect 164752 5584 164758 5596
rect 233326 5584 233332 5596
rect 233384 5584 233390 5636
rect 386322 5584 386328 5636
rect 386380 5624 386386 5636
rect 458450 5624 458456 5636
rect 386380 5596 458456 5624
rect 386380 5584 386386 5596
rect 458450 5584 458456 5596
rect 458508 5584 458514 5636
rect 80149 5559 80207 5565
rect 80149 5525 80161 5559
rect 80195 5556 80207 5559
rect 84105 5559 84163 5565
rect 84105 5556 84117 5559
rect 80195 5528 84117 5556
rect 80195 5525 80207 5528
rect 80149 5519 80207 5525
rect 84105 5525 84117 5528
rect 84151 5525 84163 5559
rect 84105 5519 84163 5525
rect 93857 5559 93915 5565
rect 93857 5525 93869 5559
rect 93903 5556 93915 5559
rect 103425 5559 103483 5565
rect 103425 5556 103437 5559
rect 93903 5528 103437 5556
rect 93903 5525 93915 5528
rect 93857 5519 93915 5525
rect 103425 5525 103437 5528
rect 103471 5525 103483 5559
rect 103425 5519 103483 5525
rect 113542 5516 113548 5568
rect 113600 5556 113606 5568
rect 160738 5556 160744 5568
rect 113600 5528 160744 5556
rect 113600 5516 113606 5528
rect 160738 5516 160744 5528
rect 160796 5516 160802 5568
rect 168190 5516 168196 5568
rect 168248 5556 168254 5568
rect 236086 5556 236092 5568
rect 168248 5528 236092 5556
rect 168248 5516 168254 5528
rect 236086 5516 236092 5528
rect 236144 5516 236150 5568
rect 384942 5516 384948 5568
rect 385000 5556 385006 5568
rect 454862 5556 454868 5568
rect 385000 5528 454868 5556
rect 385000 5516 385006 5528
rect 454862 5516 454868 5528
rect 454920 5516 454926 5568
rect 51626 5448 51632 5500
rect 51684 5488 51690 5500
rect 175458 5488 175464 5500
rect 51684 5460 175464 5488
rect 51684 5448 51690 5460
rect 175458 5448 175464 5460
rect 175516 5448 175522 5500
rect 183462 5448 183468 5500
rect 183520 5488 183526 5500
rect 183557 5491 183615 5497
rect 183557 5488 183569 5491
rect 183520 5460 183569 5488
rect 183520 5448 183526 5460
rect 183557 5457 183569 5460
rect 183603 5457 183615 5491
rect 183557 5451 183615 5457
rect 187234 5448 187240 5500
rect 187292 5488 187298 5500
rect 245654 5488 245660 5500
rect 187292 5460 245660 5488
rect 187292 5448 187298 5460
rect 245654 5448 245660 5460
rect 245712 5448 245718 5500
rect 362770 5448 362776 5500
rect 362828 5488 362834 5500
rect 412082 5488 412088 5500
rect 362828 5460 412088 5488
rect 362828 5448 362834 5460
rect 412082 5448 412088 5460
rect 412140 5448 412146 5500
rect 416590 5448 416596 5500
rect 416648 5488 416654 5500
rect 416648 5460 419396 5488
rect 416648 5448 416654 5460
rect 48130 5380 48136 5432
rect 48188 5420 48194 5432
rect 173986 5420 173992 5432
rect 48188 5392 173992 5420
rect 48188 5380 48194 5392
rect 173986 5380 173992 5392
rect 174044 5380 174050 5432
rect 174170 5380 174176 5432
rect 174228 5420 174234 5432
rect 181441 5423 181499 5429
rect 181441 5420 181453 5423
rect 174228 5392 181453 5420
rect 174228 5380 174234 5392
rect 181441 5389 181453 5392
rect 181487 5389 181499 5423
rect 181441 5383 181499 5389
rect 181530 5380 181536 5432
rect 181588 5420 181594 5432
rect 191101 5423 191159 5429
rect 181588 5392 181668 5420
rect 181588 5380 181594 5392
rect 33870 5312 33876 5364
rect 33928 5352 33934 5364
rect 55217 5355 55275 5361
rect 55217 5352 55229 5355
rect 33928 5324 55229 5352
rect 33928 5312 33934 5324
rect 55217 5321 55229 5324
rect 55263 5321 55275 5355
rect 55217 5315 55275 5321
rect 64785 5355 64843 5361
rect 64785 5321 64797 5355
rect 64831 5352 64843 5355
rect 74537 5355 74595 5361
rect 74537 5352 74549 5355
rect 64831 5324 74549 5352
rect 64831 5321 64843 5324
rect 64785 5315 64843 5321
rect 74537 5321 74549 5324
rect 74583 5321 74595 5355
rect 74537 5315 74595 5321
rect 84105 5355 84163 5361
rect 84105 5321 84117 5355
rect 84151 5352 84163 5355
rect 93854 5352 93860 5364
rect 84151 5324 93860 5352
rect 84151 5321 84163 5324
rect 84105 5315 84163 5321
rect 93854 5312 93860 5324
rect 93912 5312 93918 5364
rect 103422 5312 103428 5364
rect 103480 5352 103486 5364
rect 113174 5352 113180 5364
rect 103480 5324 113180 5352
rect 103480 5312 103486 5324
rect 113174 5312 113180 5324
rect 113232 5312 113238 5364
rect 122650 5312 122656 5364
rect 122708 5352 122714 5364
rect 132494 5352 132500 5364
rect 122708 5324 132500 5352
rect 122708 5312 122714 5324
rect 132494 5312 132500 5324
rect 132552 5312 132558 5364
rect 141970 5312 141976 5364
rect 142028 5352 142034 5364
rect 152277 5355 152335 5361
rect 142028 5324 152228 5352
rect 142028 5312 142034 5324
rect 30282 5244 30288 5296
rect 30340 5284 30346 5296
rect 152093 5287 152151 5293
rect 152093 5284 152105 5287
rect 30340 5256 152105 5284
rect 30340 5244 30346 5256
rect 152093 5253 152105 5256
rect 152139 5253 152151 5287
rect 152093 5247 152151 5253
rect 26694 5176 26700 5228
rect 26752 5216 26758 5228
rect 55217 5219 55275 5225
rect 55217 5216 55229 5219
rect 26752 5188 55229 5216
rect 26752 5176 26758 5188
rect 55217 5185 55229 5188
rect 55263 5185 55275 5219
rect 55217 5179 55275 5185
rect 64785 5219 64843 5225
rect 64785 5185 64797 5219
rect 64831 5216 64843 5219
rect 74537 5219 74595 5225
rect 74537 5216 74549 5219
rect 64831 5188 74549 5216
rect 64831 5185 64843 5188
rect 64785 5179 64843 5185
rect 74537 5185 74549 5188
rect 74583 5185 74595 5219
rect 74537 5179 74595 5185
rect 84105 5219 84163 5225
rect 84105 5185 84117 5219
rect 84151 5216 84163 5219
rect 93857 5219 93915 5225
rect 93857 5216 93869 5219
rect 84151 5188 93869 5216
rect 84151 5185 84163 5188
rect 84105 5179 84163 5185
rect 93857 5185 93869 5188
rect 93903 5185 93915 5219
rect 93857 5179 93915 5185
rect 103425 5219 103483 5225
rect 103425 5185 103437 5219
rect 103471 5216 103483 5219
rect 113177 5219 113235 5225
rect 113177 5216 113189 5219
rect 103471 5188 113189 5216
rect 103471 5185 103483 5188
rect 103425 5179 103483 5185
rect 113177 5185 113189 5188
rect 113223 5185 113235 5219
rect 113177 5179 113235 5185
rect 122745 5219 122803 5225
rect 122745 5185 122757 5219
rect 122791 5216 122803 5219
rect 132497 5219 132555 5225
rect 132497 5216 132509 5219
rect 122791 5188 132509 5216
rect 122791 5185 122803 5188
rect 122745 5179 122803 5185
rect 132497 5185 132509 5188
rect 132543 5185 132555 5219
rect 132497 5179 132555 5185
rect 142065 5219 142123 5225
rect 142065 5185 142077 5219
rect 142111 5216 142123 5219
rect 152200 5216 152228 5324
rect 152277 5321 152289 5355
rect 152323 5352 152335 5355
rect 152323 5324 152596 5352
rect 152323 5321 152335 5324
rect 152277 5315 152335 5321
rect 152568 5284 152596 5324
rect 152734 5312 152740 5364
rect 152792 5352 152798 5364
rect 162213 5355 162271 5361
rect 152792 5324 162164 5352
rect 152792 5312 152798 5324
rect 160833 5287 160891 5293
rect 160833 5284 160845 5287
rect 152568 5256 160845 5284
rect 160833 5253 160845 5256
rect 160879 5253 160891 5287
rect 162136 5284 162164 5324
rect 162213 5321 162225 5355
rect 162259 5352 162271 5355
rect 167086 5352 167092 5364
rect 162259 5324 167092 5352
rect 162259 5321 162271 5324
rect 162213 5315 162271 5321
rect 167086 5312 167092 5324
rect 167144 5312 167150 5364
rect 181640 5352 181668 5392
rect 191101 5389 191113 5423
rect 191147 5420 191159 5423
rect 244366 5420 244372 5432
rect 191147 5392 244372 5420
rect 191147 5389 191159 5392
rect 191101 5383 191159 5389
rect 244366 5380 244372 5392
rect 244424 5380 244430 5432
rect 360010 5380 360016 5432
rect 360068 5420 360074 5432
rect 408494 5420 408500 5432
rect 360068 5392 408500 5420
rect 360068 5380 360074 5392
rect 408494 5380 408500 5392
rect 408552 5380 408558 5432
rect 419368 5420 419396 5460
rect 419442 5448 419448 5500
rect 419500 5488 419506 5500
rect 422849 5491 422907 5497
rect 422849 5488 422861 5491
rect 419500 5460 422861 5488
rect 419500 5448 419506 5460
rect 422849 5457 422861 5460
rect 422895 5457 422907 5491
rect 422849 5451 422907 5457
rect 422941 5491 422999 5497
rect 422941 5457 422953 5491
rect 422987 5488 422999 5491
rect 422987 5460 432552 5488
rect 422987 5457 422999 5460
rect 422941 5451 422999 5457
rect 424045 5423 424103 5429
rect 424045 5420 424057 5423
rect 419368 5392 424057 5420
rect 424045 5389 424057 5392
rect 424091 5389 424103 5423
rect 424045 5383 424103 5389
rect 424134 5380 424140 5432
rect 424192 5420 424198 5432
rect 429930 5420 429936 5432
rect 424192 5392 429936 5420
rect 424192 5380 424198 5392
rect 429930 5380 429936 5392
rect 429988 5380 429994 5432
rect 431770 5380 431776 5432
rect 431828 5420 431834 5432
rect 432417 5423 432475 5429
rect 432417 5420 432429 5423
rect 431828 5392 432429 5420
rect 431828 5380 431834 5392
rect 432417 5389 432429 5392
rect 432463 5389 432475 5423
rect 432524 5420 432552 5460
rect 432598 5448 432604 5500
rect 432656 5488 432662 5500
rect 540514 5488 540520 5500
rect 432656 5460 540520 5488
rect 432656 5448 432662 5460
rect 540514 5448 540520 5460
rect 540572 5448 540578 5500
rect 432782 5420 432788 5432
rect 432524 5392 432788 5420
rect 432417 5383 432475 5389
rect 432782 5380 432788 5392
rect 432840 5380 432846 5432
rect 544102 5420 544108 5432
rect 432892 5392 544108 5420
rect 242986 5352 242992 5364
rect 181640 5324 242992 5352
rect 242986 5312 242992 5324
rect 243044 5312 243050 5364
rect 364242 5312 364248 5364
rect 364300 5352 364306 5364
rect 415670 5352 415676 5364
rect 364300 5324 415676 5352
rect 364300 5312 364306 5324
rect 415670 5312 415676 5324
rect 415728 5312 415734 5364
rect 430482 5312 430488 5364
rect 430540 5352 430546 5364
rect 432892 5352 432920 5392
rect 544102 5380 544108 5392
rect 544160 5380 544166 5432
rect 430540 5324 432920 5352
rect 430540 5312 430546 5324
rect 433242 5312 433248 5364
rect 433300 5352 433306 5364
rect 441525 5355 441583 5361
rect 433300 5324 433748 5352
rect 433300 5312 433306 5324
rect 178678 5284 178684 5296
rect 162136 5256 178684 5284
rect 160833 5247 160891 5253
rect 178678 5244 178684 5256
rect 178736 5244 178742 5296
rect 181441 5287 181499 5293
rect 181441 5253 181453 5287
rect 181487 5284 181499 5287
rect 238846 5284 238852 5296
rect 181487 5256 238852 5284
rect 181487 5253 181499 5256
rect 181441 5247 181499 5253
rect 238846 5244 238852 5256
rect 238904 5244 238910 5296
rect 365622 5244 365628 5296
rect 365680 5284 365686 5296
rect 419166 5284 419172 5296
rect 365680 5256 419172 5284
rect 365680 5244 365686 5256
rect 419166 5244 419172 5256
rect 419224 5244 419230 5296
rect 433720 5284 433748 5324
rect 441525 5321 441537 5355
rect 441571 5352 441583 5355
rect 547690 5352 547696 5364
rect 441571 5324 547696 5352
rect 441571 5321 441583 5324
rect 441525 5315 441583 5321
rect 547690 5312 547696 5324
rect 547748 5312 547754 5364
rect 551186 5284 551192 5296
rect 423140 5256 432736 5284
rect 433720 5256 551192 5284
rect 162213 5219 162271 5225
rect 162213 5216 162225 5219
rect 142111 5188 149100 5216
rect 152200 5188 162225 5216
rect 142111 5185 142123 5188
rect 142065 5179 142123 5185
rect 21910 5108 21916 5160
rect 21968 5148 21974 5160
rect 148965 5151 149023 5157
rect 148965 5148 148977 5151
rect 21968 5120 148977 5148
rect 21968 5108 21974 5120
rect 148965 5117 148977 5120
rect 149011 5117 149023 5151
rect 149072 5148 149100 5188
rect 162213 5185 162225 5188
rect 162259 5185 162271 5219
rect 162213 5179 162271 5185
rect 170582 5176 170588 5228
rect 170640 5216 170646 5228
rect 237374 5216 237380 5228
rect 170640 5188 237380 5216
rect 170640 5176 170646 5188
rect 237374 5176 237380 5188
rect 237432 5176 237438 5228
rect 368382 5176 368388 5228
rect 368440 5216 368446 5228
rect 422754 5216 422760 5228
rect 368440 5188 422760 5216
rect 368440 5176 368446 5188
rect 422754 5176 422760 5188
rect 422812 5176 422818 5228
rect 162854 5148 162860 5160
rect 149072 5120 162860 5148
rect 148965 5111 149023 5117
rect 162854 5108 162860 5120
rect 162912 5108 162918 5160
rect 164326 5148 164332 5160
rect 162964 5120 164332 5148
rect 17310 5040 17316 5092
rect 17368 5080 17374 5092
rect 158806 5080 158812 5092
rect 17368 5052 158812 5080
rect 17368 5040 17374 5052
rect 158806 5040 158812 5052
rect 158864 5040 158870 5092
rect 160186 5080 160192 5092
rect 158916 5052 160192 5080
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 142154 5012 142160 5024
rect 7708 4984 142160 5012
rect 7708 4972 7714 4984
rect 142154 4972 142160 4984
rect 142212 4972 142218 5024
rect 148965 5015 149023 5021
rect 148965 4981 148977 5015
rect 149011 5012 149023 5015
rect 158916 5012 158944 5052
rect 160186 5040 160192 5052
rect 160244 5040 160250 5092
rect 160833 5083 160891 5089
rect 160833 5049 160845 5083
rect 160879 5080 160891 5083
rect 162964 5080 162992 5120
rect 164326 5108 164332 5120
rect 164384 5108 164390 5160
rect 167178 5108 167184 5160
rect 167236 5148 167242 5160
rect 234798 5148 234804 5160
rect 167236 5120 234804 5148
rect 167236 5108 167242 5120
rect 234798 5108 234804 5120
rect 234856 5108 234862 5160
rect 369762 5108 369768 5160
rect 369820 5148 369826 5160
rect 422205 5151 422263 5157
rect 422205 5148 422217 5151
rect 369820 5120 422217 5148
rect 369820 5108 369826 5120
rect 422205 5117 422217 5120
rect 422251 5117 422263 5151
rect 423140 5148 423168 5256
rect 426342 5176 426348 5228
rect 426400 5216 426406 5228
rect 432509 5219 432567 5225
rect 432509 5216 432521 5219
rect 426400 5188 432521 5216
rect 426400 5176 426406 5188
rect 432509 5185 432521 5188
rect 432555 5185 432567 5219
rect 432509 5179 432567 5185
rect 422205 5111 422263 5117
rect 423048 5120 423168 5148
rect 423309 5151 423367 5157
rect 160879 5052 162992 5080
rect 160879 5049 160891 5052
rect 160833 5043 160891 5049
rect 163498 5040 163504 5092
rect 163556 5080 163562 5092
rect 233234 5080 233240 5092
rect 163556 5052 233240 5080
rect 163556 5040 163562 5052
rect 233234 5040 233240 5052
rect 233292 5040 233298 5092
rect 371050 5040 371056 5092
rect 371108 5080 371114 5092
rect 403529 5083 403587 5089
rect 403529 5080 403541 5083
rect 371108 5052 403541 5080
rect 371108 5040 371114 5052
rect 403529 5049 403541 5052
rect 403575 5049 403587 5083
rect 403529 5043 403587 5049
rect 403618 5040 403624 5092
rect 403676 5080 403682 5092
rect 412545 5083 412603 5089
rect 403676 5052 412496 5080
rect 403676 5040 403682 5052
rect 149011 4984 158944 5012
rect 149011 4981 149023 4984
rect 148965 4975 149023 4981
rect 158990 4972 158996 5024
rect 159048 5012 159054 5024
rect 230474 5012 230480 5024
rect 159048 4984 230480 5012
rect 159048 4972 159054 4984
rect 230474 4972 230480 4984
rect 230532 4972 230538 5024
rect 373810 4972 373816 5024
rect 373868 5012 373874 5024
rect 379330 5012 379336 5024
rect 373868 4984 379336 5012
rect 373868 4972 373874 4984
rect 379330 4972 379336 4984
rect 379388 4972 379394 5024
rect 379514 4972 379520 5024
rect 379572 5012 379578 5024
rect 398742 5012 398748 5024
rect 379572 4984 398748 5012
rect 379572 4972 379578 4984
rect 398742 4972 398748 4984
rect 398800 4972 398806 5024
rect 412468 5012 412496 5052
rect 412545 5049 412557 5083
rect 412591 5080 412603 5083
rect 420086 5080 420092 5092
rect 412591 5052 420092 5080
rect 412591 5049 412603 5052
rect 412545 5043 412603 5049
rect 420086 5040 420092 5052
rect 420144 5040 420150 5092
rect 423048 5012 423076 5120
rect 423309 5117 423321 5151
rect 423355 5148 423367 5151
rect 426437 5151 426495 5157
rect 426437 5148 426449 5151
rect 423355 5120 426449 5148
rect 423355 5117 423367 5120
rect 423309 5111 423367 5117
rect 426437 5117 426449 5120
rect 426483 5117 426495 5151
rect 426437 5111 426495 5117
rect 427630 5108 427636 5160
rect 427688 5148 427694 5160
rect 432598 5148 432604 5160
rect 427688 5120 432604 5148
rect 427688 5108 427694 5120
rect 432598 5108 432604 5120
rect 432656 5108 432662 5160
rect 432708 5148 432736 5256
rect 551186 5244 551192 5256
rect 551244 5244 551250 5296
rect 432877 5219 432935 5225
rect 432877 5185 432889 5219
rect 432923 5216 432935 5219
rect 437109 5219 437167 5225
rect 437109 5216 437121 5219
rect 432923 5188 437121 5216
rect 432923 5185 432935 5188
rect 432877 5179 432935 5185
rect 437109 5185 437121 5188
rect 437155 5185 437167 5219
rect 437109 5179 437167 5185
rect 437382 5176 437388 5228
rect 437440 5216 437446 5228
rect 446493 5219 446551 5225
rect 437440 5188 446444 5216
rect 437440 5176 437446 5188
rect 433518 5148 433524 5160
rect 432708 5120 433524 5148
rect 433518 5108 433524 5120
rect 433576 5108 433582 5160
rect 436002 5108 436008 5160
rect 436060 5148 436066 5160
rect 440697 5151 440755 5157
rect 440697 5148 440709 5151
rect 436060 5120 440709 5148
rect 436060 5108 436066 5120
rect 440697 5117 440709 5120
rect 440743 5117 440755 5151
rect 440697 5111 440755 5117
rect 441522 5108 441528 5160
rect 441580 5148 441586 5160
rect 446416 5148 446444 5188
rect 446493 5185 446505 5219
rect 446539 5216 446551 5219
rect 554774 5216 554780 5228
rect 446539 5188 554780 5216
rect 446539 5185 446551 5188
rect 446493 5179 446551 5185
rect 554774 5176 554780 5188
rect 554832 5176 554838 5228
rect 558362 5148 558368 5160
rect 441580 5120 446352 5148
rect 446416 5120 558368 5148
rect 441580 5108 441586 5120
rect 423140 5052 432644 5080
rect 423140 5021 423168 5052
rect 412468 4984 423076 5012
rect 423125 5015 423183 5021
rect 423125 4981 423137 5015
rect 423171 4981 423183 5015
rect 423125 4975 423183 4981
rect 423217 5015 423275 5021
rect 423217 4981 423229 5015
rect 423263 5012 423275 5015
rect 423263 4984 432552 5012
rect 423263 4981 423275 4984
rect 423217 4975 423275 4981
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 150802 4944 150808 4956
rect 2924 4916 150808 4944
rect 2924 4904 2930 4916
rect 150802 4904 150808 4916
rect 150860 4904 150866 4956
rect 150894 4904 150900 4956
rect 150952 4944 150958 4956
rect 153194 4944 153200 4956
rect 150952 4916 153200 4944
rect 150952 4904 150958 4916
rect 153194 4904 153200 4916
rect 153252 4904 153258 4956
rect 155218 4904 155224 4956
rect 155276 4944 155282 4956
rect 229094 4944 229100 4956
rect 155276 4916 229100 4944
rect 155276 4904 155282 4916
rect 229094 4904 229100 4916
rect 229152 4904 229158 4956
rect 375282 4904 375288 4956
rect 375340 4944 375346 4956
rect 375340 4916 423076 4944
rect 375340 4904 375346 4916
rect 566 4836 572 4888
rect 624 4876 630 4888
rect 149054 4876 149060 4888
rect 624 4848 149060 4876
rect 624 4836 630 4848
rect 149054 4836 149060 4848
rect 149112 4836 149118 4888
rect 149238 4836 149244 4888
rect 149296 4876 149302 4888
rect 226334 4876 226340 4888
rect 149296 4848 226340 4876
rect 149296 4836 149302 4848
rect 226334 4836 226340 4848
rect 226392 4836 226398 4888
rect 237190 4836 237196 4888
rect 237248 4876 237254 4888
rect 270586 4876 270592 4888
rect 237248 4848 270592 4876
rect 237248 4836 237254 4848
rect 270586 4836 270592 4848
rect 270644 4836 270650 4888
rect 379422 4836 379428 4888
rect 379480 4876 379486 4888
rect 398834 4876 398840 4888
rect 379480 4848 398840 4876
rect 379480 4836 379486 4848
rect 398834 4836 398840 4848
rect 398892 4836 398898 4888
rect 422941 4879 422999 4885
rect 422941 4876 422953 4879
rect 412560 4848 422953 4876
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 150526 4808 150532 4820
rect 1728 4780 150532 4808
rect 1728 4768 1734 4780
rect 150526 4768 150532 4780
rect 150584 4768 150590 4820
rect 151538 4768 151544 4820
rect 151596 4808 151602 4820
rect 227898 4808 227904 4820
rect 151596 4780 227904 4808
rect 151596 4768 151602 4780
rect 227898 4768 227904 4780
rect 227956 4768 227962 4820
rect 233694 4768 233700 4820
rect 233752 4808 233758 4820
rect 269206 4808 269212 4820
rect 233752 4780 269212 4808
rect 233752 4768 233758 4780
rect 269206 4768 269212 4780
rect 269264 4768 269270 4820
rect 376662 4768 376668 4820
rect 376720 4808 376726 4820
rect 400217 4811 400275 4817
rect 400217 4808 400229 4811
rect 376720 4780 400229 4808
rect 376720 4768 376726 4780
rect 400217 4777 400229 4780
rect 400263 4777 400275 4811
rect 404906 4808 404912 4820
rect 400217 4771 400275 4777
rect 400324 4780 404912 4808
rect 55214 4700 55220 4752
rect 55272 4740 55278 4752
rect 178034 4740 178040 4752
rect 55272 4712 178040 4740
rect 55272 4700 55278 4712
rect 178034 4700 178040 4712
rect 178092 4700 178098 4752
rect 183557 4743 183615 4749
rect 183557 4709 183569 4743
rect 183603 4740 183615 4743
rect 188341 4743 188399 4749
rect 188341 4740 188353 4743
rect 183603 4712 188353 4740
rect 183603 4709 183615 4712
rect 183557 4703 183615 4709
rect 188341 4709 188353 4712
rect 188387 4709 188399 4743
rect 188341 4703 188399 4709
rect 188430 4700 188436 4752
rect 188488 4740 188494 4752
rect 245930 4740 245936 4752
rect 188488 4712 245936 4740
rect 188488 4700 188494 4712
rect 245930 4700 245936 4712
rect 245988 4700 245994 4752
rect 358722 4700 358728 4752
rect 358780 4740 358786 4752
rect 400324 4740 400352 4780
rect 404906 4768 404912 4780
rect 404964 4768 404970 4820
rect 404998 4768 405004 4820
rect 405056 4808 405062 4820
rect 412560 4808 412588 4848
rect 422941 4845 422953 4848
rect 422987 4845 422999 4879
rect 423048 4876 423076 4916
rect 432414 4876 432420 4888
rect 423048 4848 432420 4876
rect 422941 4839 422999 4845
rect 432414 4836 432420 4848
rect 432472 4836 432478 4888
rect 432524 4876 432552 4984
rect 432616 4944 432644 5052
rect 432782 5040 432788 5092
rect 432840 5080 432846 5092
rect 441617 5083 441675 5089
rect 441617 5080 441629 5083
rect 432840 5052 441629 5080
rect 432840 5040 432846 5052
rect 441617 5049 441629 5052
rect 441663 5049 441675 5083
rect 446324 5080 446352 5120
rect 558362 5108 558368 5120
rect 558420 5108 558426 5160
rect 565538 5080 565544 5092
rect 446324 5052 565544 5080
rect 441617 5043 441675 5049
rect 565538 5040 565544 5052
rect 565596 5040 565602 5092
rect 432690 4972 432696 5024
rect 432748 5012 432754 5024
rect 437014 5012 437020 5024
rect 432748 4984 437020 5012
rect 432748 4972 432754 4984
rect 437014 4972 437020 4984
rect 437072 4972 437078 5024
rect 437109 5015 437167 5021
rect 437109 4981 437121 5015
rect 437155 5012 437167 5015
rect 438305 5015 438363 5021
rect 438305 5012 438317 5015
rect 437155 4984 438317 5012
rect 437155 4981 437167 4984
rect 437109 4975 437167 4981
rect 438305 4981 438317 4984
rect 438351 4981 438363 5015
rect 438305 4975 438363 4981
rect 438670 4972 438676 5024
rect 438728 5012 438734 5024
rect 561950 5012 561956 5024
rect 438728 4984 561956 5012
rect 438728 4972 438734 4984
rect 561950 4972 561956 4984
rect 562008 4972 562014 5024
rect 440602 4944 440608 4956
rect 432616 4916 440608 4944
rect 440602 4904 440608 4916
rect 440660 4904 440666 4956
rect 440697 4947 440755 4953
rect 440697 4913 440709 4947
rect 440743 4944 440755 4947
rect 446493 4947 446551 4953
rect 446493 4944 446505 4947
rect 440743 4916 446505 4944
rect 440743 4913 440755 4916
rect 440697 4907 440755 4913
rect 446493 4913 446505 4916
rect 446539 4913 446551 4947
rect 446493 4907 446551 4913
rect 446585 4947 446643 4953
rect 446585 4913 446597 4947
rect 446631 4944 446643 4947
rect 569034 4944 569040 4956
rect 446631 4916 569040 4944
rect 446631 4913 446643 4916
rect 446585 4907 446643 4913
rect 569034 4904 569040 4916
rect 569092 4904 569098 4956
rect 432785 4879 432843 4885
rect 432524 4848 432736 4876
rect 423125 4811 423183 4817
rect 423125 4808 423137 4811
rect 405056 4780 412588 4808
rect 417436 4780 423137 4808
rect 405056 4768 405062 4780
rect 358780 4712 400352 4740
rect 400401 4743 400459 4749
rect 358780 4700 358786 4712
rect 400401 4709 400413 4743
rect 400447 4740 400459 4743
rect 417436 4740 417464 4780
rect 423125 4777 423137 4780
rect 423171 4777 423183 4811
rect 423125 4771 423183 4777
rect 423309 4811 423367 4817
rect 423309 4777 423321 4811
rect 423355 4808 423367 4811
rect 427630 4808 427636 4820
rect 423355 4780 427636 4808
rect 423355 4777 423367 4780
rect 423309 4771 423367 4777
rect 427630 4768 427636 4780
rect 427688 4768 427694 4820
rect 427817 4811 427875 4817
rect 427817 4777 427829 4811
rect 427863 4808 427875 4811
rect 431126 4808 431132 4820
rect 427863 4780 431132 4808
rect 427863 4777 427875 4780
rect 427817 4771 427875 4777
rect 431126 4768 431132 4780
rect 431184 4768 431190 4820
rect 432601 4811 432659 4817
rect 432601 4777 432613 4811
rect 432647 4777 432659 4811
rect 432708 4808 432736 4848
rect 432785 4845 432797 4879
rect 432831 4876 432843 4879
rect 438210 4876 438216 4888
rect 432831 4848 438216 4876
rect 432831 4845 432843 4848
rect 432785 4839 432843 4845
rect 438210 4836 438216 4848
rect 438268 4836 438274 4888
rect 438305 4879 438363 4885
rect 438305 4845 438317 4879
rect 438351 4876 438363 4879
rect 441525 4879 441583 4885
rect 441525 4876 441537 4879
rect 438351 4848 441537 4876
rect 438351 4845 438363 4848
rect 438305 4839 438363 4845
rect 441525 4845 441537 4848
rect 441571 4845 441583 4879
rect 441525 4839 441583 4845
rect 441893 4879 441951 4885
rect 441893 4845 441905 4879
rect 441939 4876 441951 4879
rect 444190 4876 444196 4888
rect 441939 4848 444196 4876
rect 441939 4845 441951 4848
rect 441893 4839 441951 4845
rect 444190 4836 444196 4848
rect 444248 4836 444254 4888
rect 444282 4836 444288 4888
rect 444340 4876 444346 4888
rect 572622 4876 572628 4888
rect 444340 4848 572628 4876
rect 444340 4836 444346 4848
rect 572622 4836 572628 4848
rect 572680 4836 572686 4888
rect 441798 4808 441804 4820
rect 432708 4780 441804 4808
rect 432601 4771 432659 4777
rect 400447 4712 417464 4740
rect 400447 4709 400459 4712
rect 400401 4703 400459 4709
rect 422202 4700 422208 4752
rect 422260 4740 422266 4752
rect 422849 4743 422907 4749
rect 422849 4740 422861 4743
rect 422260 4712 422861 4740
rect 422260 4700 422266 4712
rect 422849 4709 422861 4712
rect 422895 4709 422907 4743
rect 432616 4740 432644 4771
rect 441798 4768 441804 4780
rect 441856 4768 441862 4820
rect 442810 4768 442816 4820
rect 442868 4808 442874 4820
rect 446585 4811 446643 4817
rect 446585 4808 446597 4811
rect 442868 4780 446597 4808
rect 442868 4768 442874 4780
rect 446585 4777 446597 4780
rect 446631 4777 446643 4811
rect 446585 4771 446643 4777
rect 447042 4768 447048 4820
rect 447100 4808 447106 4820
rect 576210 4808 576216 4820
rect 447100 4780 576216 4808
rect 447100 4768 447106 4780
rect 576210 4768 576216 4780
rect 576268 4768 576274 4820
rect 422849 4703 422907 4709
rect 422956 4712 432644 4740
rect 432693 4743 432751 4749
rect 58802 4632 58808 4684
rect 58860 4672 58866 4684
rect 179506 4672 179512 4684
rect 58860 4644 179512 4672
rect 58860 4632 58866 4644
rect 179506 4632 179512 4644
rect 179564 4632 179570 4684
rect 184842 4632 184848 4684
rect 184900 4672 184906 4684
rect 191101 4675 191159 4681
rect 191101 4672 191113 4675
rect 184900 4644 191113 4672
rect 184900 4632 184906 4644
rect 191101 4641 191113 4644
rect 191147 4641 191159 4675
rect 191101 4635 191159 4641
rect 194410 4632 194416 4684
rect 194468 4672 194474 4684
rect 249978 4672 249984 4684
rect 194468 4644 249984 4672
rect 194468 4632 194474 4644
rect 249978 4632 249984 4644
rect 250036 4632 250042 4684
rect 354582 4632 354588 4684
rect 354640 4672 354646 4684
rect 397822 4672 397828 4684
rect 354640 4644 397828 4672
rect 354640 4632 354646 4644
rect 397822 4632 397828 4644
rect 397880 4632 397886 4684
rect 398098 4632 398104 4684
rect 398156 4672 398162 4684
rect 398834 4672 398840 4684
rect 398156 4644 398840 4672
rect 398156 4632 398162 4644
rect 398834 4632 398840 4644
rect 398892 4632 398898 4684
rect 422757 4675 422815 4681
rect 422757 4672 422769 4675
rect 412376 4644 422769 4672
rect 55217 4607 55275 4613
rect 55217 4573 55229 4607
rect 55263 4604 55275 4607
rect 64785 4607 64843 4613
rect 64785 4604 64797 4607
rect 55263 4576 64797 4604
rect 55263 4573 55275 4576
rect 55217 4567 55275 4573
rect 64785 4573 64797 4576
rect 64831 4573 64843 4607
rect 64785 4567 64843 4573
rect 65978 4564 65984 4616
rect 66036 4604 66042 4616
rect 183554 4604 183560 4616
rect 66036 4576 183560 4604
rect 66036 4564 66042 4576
rect 183554 4564 183560 4576
rect 183612 4564 183618 4616
rect 192018 4564 192024 4616
rect 192076 4604 192082 4616
rect 248506 4604 248512 4616
rect 192076 4576 248512 4604
rect 192076 4564 192082 4576
rect 248506 4564 248512 4576
rect 248564 4564 248570 4616
rect 353202 4564 353208 4616
rect 353260 4604 353266 4616
rect 394234 4604 394240 4616
rect 353260 4576 394240 4604
rect 353260 4564 353266 4576
rect 394234 4564 394240 4576
rect 394292 4564 394298 4616
rect 394418 4564 394424 4616
rect 394476 4604 394482 4616
rect 403621 4607 403679 4613
rect 403621 4604 403633 4607
rect 394476 4576 403633 4604
rect 394476 4564 394482 4576
rect 403621 4573 403633 4576
rect 403667 4573 403679 4607
rect 403621 4567 403679 4573
rect 403710 4564 403716 4616
rect 403768 4604 403774 4616
rect 412376 4604 412404 4644
rect 422757 4641 422769 4644
rect 422803 4641 422815 4675
rect 422757 4635 422815 4641
rect 403768 4576 412404 4604
rect 412453 4607 412511 4613
rect 403768 4564 403774 4576
rect 412453 4573 412465 4607
rect 412499 4604 412511 4607
rect 422956 4604 422984 4712
rect 432693 4709 432705 4743
rect 432739 4740 432751 4743
rect 536926 4740 536932 4752
rect 432739 4712 536932 4740
rect 432739 4709 432751 4712
rect 432693 4703 432751 4709
rect 536926 4700 536932 4712
rect 536984 4700 536990 4752
rect 424778 4632 424784 4684
rect 424836 4672 424842 4684
rect 533430 4672 533436 4684
rect 424836 4644 533436 4672
rect 424836 4632 424842 4644
rect 533430 4632 533436 4644
rect 533488 4632 533494 4684
rect 412499 4576 422984 4604
rect 423033 4607 423091 4613
rect 412499 4573 412511 4576
rect 412453 4567 412511 4573
rect 423033 4573 423045 4607
rect 423079 4604 423091 4607
rect 529842 4604 529848 4616
rect 423079 4576 529848 4604
rect 423079 4573 423091 4576
rect 423033 4567 423091 4573
rect 529842 4564 529848 4576
rect 529900 4564 529906 4616
rect 62390 4496 62396 4548
rect 62448 4536 62454 4548
rect 180978 4536 180984 4548
rect 62448 4508 180984 4536
rect 62448 4496 62454 4508
rect 180978 4496 180984 4508
rect 181036 4496 181042 4548
rect 190822 4496 190828 4548
rect 190880 4536 190886 4548
rect 247310 4536 247316 4548
rect 190880 4508 247316 4536
rect 190880 4496 190886 4508
rect 247310 4496 247316 4508
rect 247368 4496 247374 4548
rect 357158 4496 357164 4548
rect 357216 4536 357222 4548
rect 401318 4536 401324 4548
rect 357216 4508 401324 4536
rect 357216 4496 357222 4508
rect 401318 4496 401324 4508
rect 401376 4496 401382 4548
rect 401410 4496 401416 4548
rect 401468 4536 401474 4548
rect 403434 4536 403440 4548
rect 401468 4508 403440 4536
rect 401468 4496 401474 4508
rect 403434 4496 403440 4508
rect 403492 4496 403498 4548
rect 403529 4539 403587 4545
rect 403529 4505 403541 4539
rect 403575 4536 403587 4539
rect 412545 4539 412603 4545
rect 412545 4536 412557 4539
rect 403575 4508 412557 4536
rect 403575 4505 403587 4508
rect 403529 4499 403587 4505
rect 412545 4505 412557 4508
rect 412591 4505 412603 4539
rect 412545 4499 412603 4505
rect 422205 4539 422263 4545
rect 422205 4505 422217 4539
rect 422251 4536 422263 4539
rect 426342 4536 426348 4548
rect 422251 4508 426348 4536
rect 422251 4505 422263 4508
rect 422205 4499 422263 4505
rect 426342 4496 426348 4508
rect 426400 4496 426406 4548
rect 426437 4539 426495 4545
rect 426437 4505 426449 4539
rect 426483 4536 426495 4539
rect 526254 4536 526260 4548
rect 426483 4508 526260 4536
rect 426483 4505 426495 4508
rect 426437 4499 426495 4505
rect 526254 4496 526260 4508
rect 526312 4496 526318 4548
rect 55309 4471 55367 4477
rect 55309 4437 55321 4471
rect 55355 4468 55367 4471
rect 64693 4471 64751 4477
rect 64693 4468 64705 4471
rect 55355 4440 64705 4468
rect 55355 4437 55367 4440
rect 55309 4431 55367 4437
rect 64693 4437 64705 4440
rect 64739 4437 64751 4471
rect 64693 4431 64751 4437
rect 69474 4428 69480 4480
rect 69532 4468 69538 4480
rect 185210 4468 185216 4480
rect 69532 4440 185216 4468
rect 69532 4428 69538 4440
rect 185210 4428 185216 4440
rect 185268 4428 185274 4480
rect 195606 4428 195612 4480
rect 195664 4468 195670 4480
rect 249886 4468 249892 4480
rect 195664 4440 249892 4468
rect 195664 4428 195670 4440
rect 249886 4428 249892 4440
rect 249944 4428 249950 4480
rect 351822 4428 351828 4480
rect 351880 4468 351886 4480
rect 391842 4468 391848 4480
rect 351880 4440 391848 4468
rect 351880 4428 351886 4440
rect 391842 4428 391848 4440
rect 391900 4428 391906 4480
rect 391952 4440 394648 4468
rect 73062 4360 73068 4412
rect 73120 4400 73126 4412
rect 186406 4400 186412 4412
rect 73120 4372 186412 4400
rect 73120 4360 73126 4372
rect 186406 4360 186412 4372
rect 186464 4360 186470 4412
rect 188341 4403 188399 4409
rect 188341 4369 188353 4403
rect 188387 4400 188399 4403
rect 188387 4372 189212 4400
rect 188387 4369 188399 4372
rect 188341 4363 188399 4369
rect 76650 4292 76656 4344
rect 76708 4332 76714 4344
rect 189074 4332 189080 4344
rect 76708 4304 189080 4332
rect 76708 4292 76714 4304
rect 189074 4292 189080 4304
rect 189132 4292 189138 4344
rect 189184 4332 189212 4372
rect 198090 4360 198096 4412
rect 198148 4400 198154 4412
rect 251266 4400 251272 4412
rect 198148 4372 251272 4400
rect 198148 4360 198154 4372
rect 251266 4360 251272 4372
rect 251324 4360 251330 4412
rect 351730 4360 351736 4412
rect 351788 4400 351794 4412
rect 390646 4400 390652 4412
rect 351788 4372 390652 4400
rect 351788 4360 351794 4372
rect 390646 4360 390652 4372
rect 390704 4360 390710 4412
rect 391382 4360 391388 4412
rect 391440 4400 391446 4412
rect 391952 4400 391980 4440
rect 391440 4372 391980 4400
rect 393869 4403 393927 4409
rect 391440 4360 391446 4372
rect 393869 4369 393881 4403
rect 393915 4400 393927 4403
rect 394620 4400 394648 4440
rect 394694 4428 394700 4480
rect 394752 4468 394758 4480
rect 423950 4468 423956 4480
rect 394752 4440 423956 4468
rect 394752 4428 394758 4440
rect 423950 4428 423956 4440
rect 424008 4428 424014 4480
rect 424045 4471 424103 4477
rect 424045 4437 424057 4471
rect 424091 4468 424103 4471
rect 519078 4468 519084 4480
rect 424091 4440 519084 4468
rect 424091 4437 424103 4440
rect 424045 4431 424103 4437
rect 519078 4428 519084 4440
rect 519136 4428 519142 4480
rect 427817 4403 427875 4409
rect 427817 4400 427829 4403
rect 393915 4372 394096 4400
rect 394620 4372 427829 4400
rect 393915 4369 393927 4372
rect 393869 4363 393927 4369
rect 200758 4332 200764 4344
rect 189184 4304 200764 4332
rect 200758 4292 200764 4304
rect 200816 4292 200822 4344
rect 201494 4292 201500 4344
rect 201552 4332 201558 4344
rect 252830 4332 252836 4344
rect 201552 4304 252836 4332
rect 201552 4292 201558 4304
rect 252830 4292 252836 4304
rect 252888 4292 252894 4344
rect 350442 4292 350448 4344
rect 350500 4332 350506 4344
rect 388254 4332 388260 4344
rect 350500 4304 388260 4332
rect 350500 4292 350506 4304
rect 388254 4292 388260 4304
rect 388312 4292 388318 4344
rect 388349 4335 388407 4341
rect 388349 4301 388361 4335
rect 388395 4332 388407 4335
rect 394068 4332 394096 4372
rect 427817 4369 427829 4372
rect 427863 4369 427875 4403
rect 427817 4363 427875 4369
rect 427906 4360 427912 4412
rect 427964 4400 427970 4412
rect 522666 4400 522672 4412
rect 427964 4372 522672 4400
rect 427964 4360 427970 4372
rect 522666 4360 522672 4372
rect 522724 4360 522730 4412
rect 409690 4332 409696 4344
rect 388395 4304 394004 4332
rect 394068 4304 409696 4332
rect 388395 4301 388407 4304
rect 388349 4295 388407 4301
rect 74629 4267 74687 4273
rect 74629 4233 74641 4267
rect 74675 4264 74687 4267
rect 80149 4267 80207 4273
rect 80149 4264 80161 4267
rect 74675 4236 80161 4264
rect 74675 4233 74687 4236
rect 74629 4227 74687 4233
rect 80149 4233 80161 4236
rect 80195 4233 80207 4267
rect 80149 4227 80207 4233
rect 80238 4224 80244 4276
rect 80296 4264 80302 4276
rect 190454 4264 190460 4276
rect 80296 4236 190460 4264
rect 80296 4224 80302 4236
rect 190454 4224 190460 4236
rect 190512 4224 190518 4276
rect 205082 4224 205088 4276
rect 205140 4264 205146 4276
rect 255406 4264 255412 4276
rect 205140 4236 255412 4264
rect 205140 4224 205146 4236
rect 255406 4224 255412 4236
rect 255464 4224 255470 4276
rect 347682 4224 347688 4276
rect 347740 4264 347746 4276
rect 384666 4264 384672 4276
rect 347740 4236 384672 4264
rect 347740 4224 347746 4236
rect 384666 4224 384672 4236
rect 384724 4224 384730 4276
rect 384776 4236 388484 4264
rect 74537 4199 74595 4205
rect 74537 4165 74549 4199
rect 74583 4196 74595 4199
rect 83737 4199 83795 4205
rect 83737 4196 83749 4199
rect 74583 4168 83749 4196
rect 74583 4165 74595 4168
rect 74537 4159 74595 4165
rect 83737 4165 83749 4168
rect 83783 4165 83795 4199
rect 83737 4159 83795 4165
rect 83826 4156 83832 4208
rect 83884 4196 83890 4208
rect 191834 4196 191840 4208
rect 83884 4168 191840 4196
rect 83884 4156 83890 4168
rect 191834 4156 191840 4168
rect 191892 4156 191898 4208
rect 212258 4156 212264 4208
rect 212316 4196 212322 4208
rect 258074 4196 258080 4208
rect 212316 4168 258080 4196
rect 212316 4156 212322 4168
rect 258074 4156 258080 4168
rect 258132 4156 258138 4208
rect 346210 4156 346216 4208
rect 346268 4196 346274 4208
rect 381170 4196 381176 4208
rect 346268 4168 381176 4196
rect 346268 4156 346274 4168
rect 381170 4156 381176 4168
rect 381228 4156 381234 4208
rect 382182 4156 382188 4208
rect 382240 4196 382246 4208
rect 382240 4168 384436 4196
rect 382240 4156 382246 4168
rect 39758 4088 39764 4140
rect 39816 4128 39822 4140
rect 42058 4128 42064 4140
rect 39816 4100 42064 4128
rect 39816 4088 39822 4100
rect 42058 4088 42064 4100
rect 42116 4088 42122 4140
rect 61194 4088 61200 4140
rect 61252 4128 61258 4140
rect 175918 4128 175924 4140
rect 61252 4100 175924 4128
rect 61252 4088 61258 4100
rect 175918 4088 175924 4100
rect 175976 4088 175982 4140
rect 191193 4131 191251 4137
rect 191193 4097 191205 4131
rect 191239 4128 191251 4131
rect 196713 4131 196771 4137
rect 196713 4128 196725 4131
rect 191239 4100 196725 4128
rect 191239 4097 191251 4100
rect 191193 4091 191251 4097
rect 196713 4097 196725 4100
rect 196759 4097 196771 4131
rect 196713 4091 196771 4097
rect 196802 4088 196808 4140
rect 196860 4128 196866 4140
rect 197262 4128 197268 4140
rect 196860 4100 197268 4128
rect 196860 4088 196866 4100
rect 197262 4088 197268 4100
rect 197320 4088 197326 4140
rect 199194 4088 199200 4140
rect 199252 4128 199258 4140
rect 203518 4128 203524 4140
rect 199252 4100 203524 4128
rect 199252 4088 199258 4100
rect 203518 4088 203524 4100
rect 203576 4088 203582 4140
rect 207474 4088 207480 4140
rect 207532 4128 207538 4140
rect 208302 4128 208308 4140
rect 207532 4100 208308 4128
rect 207532 4088 207538 4100
rect 208302 4088 208308 4100
rect 208360 4088 208366 4140
rect 211062 4088 211068 4140
rect 211120 4128 211126 4140
rect 211798 4128 211804 4140
rect 211120 4100 211804 4128
rect 211120 4088 211126 4100
rect 211798 4088 211804 4100
rect 211856 4088 211862 4140
rect 214650 4088 214656 4140
rect 214708 4128 214714 4140
rect 215202 4128 215208 4140
rect 214708 4100 215208 4128
rect 214708 4088 214714 4100
rect 215202 4088 215208 4100
rect 215260 4088 215266 4140
rect 222930 4088 222936 4140
rect 222988 4128 222994 4140
rect 263686 4128 263692 4140
rect 222988 4100 263692 4128
rect 222988 4088 222994 4100
rect 263686 4088 263692 4100
rect 263744 4088 263750 4140
rect 265802 4088 265808 4140
rect 265860 4128 265866 4140
rect 266262 4128 266268 4140
rect 265860 4100 266268 4128
rect 265860 4088 265866 4100
rect 266262 4088 266268 4100
rect 266320 4088 266326 4140
rect 268102 4088 268108 4140
rect 268160 4128 268166 4140
rect 269022 4128 269028 4140
rect 268160 4100 269028 4128
rect 268160 4088 268166 4100
rect 269022 4088 269028 4100
rect 269080 4088 269086 4140
rect 269298 4088 269304 4140
rect 269356 4128 269362 4140
rect 270402 4128 270408 4140
rect 269356 4100 270408 4128
rect 269356 4088 269362 4100
rect 270402 4088 270408 4100
rect 270460 4088 270466 4140
rect 274082 4088 274088 4140
rect 274140 4128 274146 4140
rect 274542 4128 274548 4140
rect 274140 4100 274548 4128
rect 274140 4088 274146 4100
rect 274542 4088 274548 4100
rect 274600 4088 274606 4140
rect 291930 4088 291936 4140
rect 291988 4128 291994 4140
rect 292482 4128 292488 4140
rect 291988 4100 292488 4128
rect 291988 4088 291994 4100
rect 292482 4088 292488 4100
rect 292540 4088 292546 4140
rect 295518 4088 295524 4140
rect 295576 4128 295582 4140
rect 298738 4128 298744 4140
rect 295576 4100 298744 4128
rect 295576 4088 295582 4100
rect 298738 4088 298744 4100
rect 298796 4088 298802 4140
rect 303798 4088 303804 4140
rect 303856 4128 303862 4140
rect 304902 4128 304908 4140
rect 303856 4100 304908 4128
rect 303856 4088 303862 4100
rect 304902 4088 304908 4100
rect 304960 4088 304966 4140
rect 304994 4088 305000 4140
rect 305052 4128 305058 4140
rect 306190 4128 306196 4140
rect 305052 4100 306196 4128
rect 305052 4088 305058 4100
rect 306190 4088 306196 4100
rect 306248 4088 306254 4140
rect 308030 4088 308036 4140
rect 308088 4128 308094 4140
rect 308582 4128 308588 4140
rect 308088 4100 308588 4128
rect 308088 4088 308094 4100
rect 308582 4088 308588 4100
rect 308640 4088 308646 4140
rect 310422 4088 310428 4140
rect 310480 4128 310486 4140
rect 310974 4128 310980 4140
rect 310480 4100 310980 4128
rect 310480 4088 310486 4100
rect 310974 4088 310980 4100
rect 311032 4088 311038 4140
rect 324130 4088 324136 4140
rect 324188 4128 324194 4140
rect 337102 4128 337108 4140
rect 324188 4100 337108 4128
rect 324188 4088 324194 4100
rect 337102 4088 337108 4100
rect 337160 4088 337166 4140
rect 338850 4088 338856 4140
rect 338908 4128 338914 4140
rect 338908 4100 342852 4128
rect 338908 4088 338914 4100
rect 54018 4020 54024 4072
rect 54076 4060 54082 4072
rect 174538 4060 174544 4072
rect 54076 4032 174544 4060
rect 54076 4020 54082 4032
rect 174538 4020 174544 4032
rect 174596 4020 174602 4072
rect 189626 4020 189632 4072
rect 189684 4060 189690 4072
rect 198182 4060 198188 4072
rect 189684 4032 198188 4060
rect 189684 4020 189690 4032
rect 198182 4020 198188 4032
rect 198240 4020 198246 4072
rect 220538 4020 220544 4072
rect 220596 4060 220602 4072
rect 261478 4060 261484 4072
rect 220596 4032 261484 4060
rect 220596 4020 220602 4032
rect 261478 4020 261484 4032
rect 261536 4020 261542 4072
rect 268286 4060 268292 4072
rect 262508 4032 268292 4060
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 17218 3992 17224 4004
rect 14884 3964 17224 3992
rect 14884 3952 14890 3964
rect 17218 3952 17224 3964
rect 17276 3952 17282 4004
rect 43346 3952 43352 4004
rect 43404 3992 43410 4004
rect 171134 3992 171140 4004
rect 43404 3964 171140 3992
rect 43404 3952 43410 3964
rect 171134 3952 171140 3964
rect 171192 3952 171198 4004
rect 186038 3952 186044 4004
rect 186096 3992 186102 4004
rect 199378 3992 199384 4004
rect 186096 3964 199384 3992
rect 186096 3952 186102 3964
rect 199378 3952 199384 3964
rect 199436 3952 199442 4004
rect 202690 3952 202696 4004
rect 202748 3992 202754 4004
rect 209317 3995 209375 4001
rect 202748 3964 208808 3992
rect 202748 3952 202754 3964
rect 24302 3884 24308 3936
rect 24360 3924 24366 3936
rect 28258 3924 28264 3936
rect 24360 3896 28264 3924
rect 24360 3884 24366 3896
rect 28258 3884 28264 3896
rect 28316 3884 28322 3936
rect 42150 3884 42156 3936
rect 42208 3924 42214 3936
rect 171226 3924 171232 3936
rect 42208 3896 171232 3924
rect 42208 3884 42214 3896
rect 171226 3884 171232 3896
rect 171284 3884 171290 3936
rect 177758 3884 177764 3936
rect 177816 3924 177822 3936
rect 177816 3896 181668 3924
rect 177816 3884 177822 3896
rect 36170 3816 36176 3868
rect 36228 3856 36234 3868
rect 168374 3856 168380 3868
rect 36228 3828 168380 3856
rect 36228 3816 36234 3828
rect 168374 3816 168380 3828
rect 168432 3816 168438 3868
rect 180150 3816 180156 3868
rect 180208 3856 180214 3868
rect 181640 3856 181668 3896
rect 182542 3884 182548 3936
rect 182600 3924 182606 3936
rect 202138 3924 202144 3936
rect 182600 3896 202144 3924
rect 182600 3884 182606 3896
rect 202138 3884 202144 3896
rect 202196 3884 202202 3936
rect 208780 3924 208808 3964
rect 209317 3961 209329 3995
rect 209363 3992 209375 3995
rect 216493 3995 216551 4001
rect 216493 3992 216505 3995
rect 209363 3964 216505 3992
rect 209363 3961 209375 3964
rect 209317 3955 209375 3961
rect 216493 3961 216505 3964
rect 216539 3961 216551 3995
rect 216493 3955 216551 3961
rect 219342 3952 219348 4004
rect 219400 3992 219406 4004
rect 262398 3992 262404 4004
rect 219400 3964 262404 3992
rect 219400 3952 219406 3964
rect 262398 3952 262404 3964
rect 262456 3952 262462 4004
rect 211890 3924 211896 3936
rect 208780 3896 211896 3924
rect 211890 3884 211896 3896
rect 211948 3884 211954 3936
rect 215846 3884 215852 3936
rect 215904 3924 215910 3936
rect 261018 3924 261024 3936
rect 215904 3896 261024 3924
rect 215904 3884 215910 3896
rect 261018 3884 261024 3896
rect 261076 3884 261082 3936
rect 262508 3924 262536 4032
rect 268286 4020 268292 4032
rect 268344 4020 268350 4072
rect 268381 4063 268439 4069
rect 268381 4029 268393 4063
rect 268427 4060 268439 4063
rect 276014 4060 276020 4072
rect 268427 4032 276020 4060
rect 268427 4029 268439 4032
rect 268381 4023 268439 4029
rect 276014 4020 276020 4032
rect 276072 4020 276078 4072
rect 302602 4020 302608 4072
rect 302660 4060 302666 4072
rect 304258 4060 304264 4072
rect 302660 4032 304264 4060
rect 302660 4020 302666 4032
rect 304258 4020 304264 4032
rect 304316 4020 304322 4072
rect 321462 4020 321468 4072
rect 321520 4060 321526 4072
rect 332410 4060 332416 4072
rect 321520 4032 332416 4060
rect 321520 4020 321526 4032
rect 332410 4020 332416 4032
rect 332468 4020 332474 4072
rect 333238 4020 333244 4072
rect 333296 4060 333302 4072
rect 342717 4063 342775 4069
rect 342717 4060 342729 4063
rect 333296 4032 342729 4060
rect 333296 4020 333302 4032
rect 342717 4029 342729 4032
rect 342763 4029 342775 4063
rect 342824 4060 342852 4100
rect 342898 4088 342904 4140
rect 342956 4128 342962 4140
rect 344278 4128 344284 4140
rect 342956 4100 344284 4128
rect 342956 4088 342962 4100
rect 344278 4088 344284 4100
rect 344336 4088 344342 4140
rect 345658 4088 345664 4140
rect 345716 4128 345722 4140
rect 360930 4128 360936 4140
rect 345716 4100 360936 4128
rect 345716 4088 345722 4100
rect 360930 4088 360936 4100
rect 360988 4088 360994 4140
rect 376018 4088 376024 4140
rect 376076 4128 376082 4140
rect 377582 4128 377588 4140
rect 376076 4100 377588 4128
rect 376076 4088 376082 4100
rect 377582 4088 377588 4100
rect 377640 4088 377646 4140
rect 384408 4128 384436 4168
rect 384776 4128 384804 4236
rect 384850 4156 384856 4208
rect 384908 4196 384914 4208
rect 388349 4199 388407 4205
rect 388349 4196 388361 4199
rect 384908 4168 388361 4196
rect 384908 4156 384914 4168
rect 388349 4165 388361 4168
rect 388395 4165 388407 4199
rect 388456 4196 388484 4236
rect 388622 4224 388628 4276
rect 388680 4264 388686 4276
rect 393869 4267 393927 4273
rect 393869 4264 393881 4267
rect 388680 4236 393881 4264
rect 388680 4224 388686 4236
rect 393869 4233 393881 4236
rect 393915 4233 393927 4267
rect 393976 4264 394004 4304
rect 409690 4292 409696 4304
rect 409748 4292 409754 4344
rect 415302 4292 415308 4344
rect 415360 4332 415366 4344
rect 515582 4332 515588 4344
rect 415360 4304 515588 4332
rect 415360 4292 415366 4304
rect 515582 4292 515588 4304
rect 515640 4292 515646 4344
rect 402514 4264 402520 4276
rect 393976 4236 402520 4264
rect 393869 4227 393927 4233
rect 402514 4224 402520 4236
rect 402572 4224 402578 4276
rect 403621 4267 403679 4273
rect 403621 4233 403633 4267
rect 403667 4264 403679 4267
rect 412453 4267 412511 4273
rect 412453 4264 412465 4267
rect 403667 4236 412465 4264
rect 403667 4233 403679 4236
rect 403621 4227 403679 4233
rect 412453 4233 412465 4236
rect 412499 4233 412511 4267
rect 412453 4227 412511 4233
rect 413922 4224 413928 4276
rect 413980 4264 413986 4276
rect 511994 4264 512000 4276
rect 413980 4236 512000 4264
rect 413980 4224 413986 4236
rect 511994 4224 512000 4236
rect 512052 4224 512058 4276
rect 451274 4196 451280 4208
rect 388456 4168 451280 4196
rect 388349 4159 388407 4165
rect 451274 4156 451280 4168
rect 451332 4156 451338 4208
rect 384408 4100 384804 4128
rect 385678 4088 385684 4140
rect 385736 4128 385742 4140
rect 387058 4128 387064 4140
rect 385736 4100 387064 4128
rect 385736 4088 385742 4100
rect 387058 4088 387064 4100
rect 387116 4088 387122 4140
rect 395430 4088 395436 4140
rect 395488 4128 395494 4140
rect 475102 4128 475108 4140
rect 395488 4100 475108 4128
rect 395488 4088 395494 4100
rect 475102 4088 475108 4100
rect 475160 4088 475166 4140
rect 507118 4088 507124 4140
rect 507176 4128 507182 4140
rect 514386 4128 514392 4140
rect 507176 4100 514392 4128
rect 507176 4088 507182 4100
rect 514386 4088 514392 4100
rect 514444 4088 514450 4140
rect 525058 4088 525064 4140
rect 525116 4128 525122 4140
rect 557166 4128 557172 4140
rect 525116 4100 557172 4128
rect 525116 4088 525122 4100
rect 557166 4088 557172 4100
rect 557224 4088 557230 4140
rect 345753 4063 345811 4069
rect 345753 4060 345765 4063
rect 342824 4032 345765 4060
rect 342717 4023 342775 4029
rect 345753 4029 345765 4032
rect 345799 4029 345811 4063
rect 345753 4023 345811 4029
rect 349062 4020 349068 4072
rect 349120 4060 349126 4072
rect 385862 4060 385868 4072
rect 349120 4032 385868 4060
rect 349120 4020 349126 4032
rect 385862 4020 385868 4032
rect 385920 4020 385926 4072
rect 395246 4020 395252 4072
rect 395304 4060 395310 4072
rect 410886 4060 410892 4072
rect 395304 4032 410892 4060
rect 395304 4020 395310 4032
rect 410886 4020 410892 4032
rect 410944 4020 410950 4072
rect 423214 4020 423220 4072
rect 423272 4060 423278 4072
rect 510798 4060 510804 4072
rect 423272 4032 510804 4060
rect 423272 4020 423278 4032
rect 510798 4020 510804 4032
rect 510856 4020 510862 4072
rect 511258 4020 511264 4072
rect 511316 4060 511322 4072
rect 521470 4060 521476 4072
rect 511316 4032 521476 4060
rect 511316 4020 511322 4032
rect 521470 4020 521476 4032
rect 521528 4020 521534 4072
rect 527818 4020 527824 4072
rect 527876 4060 527882 4072
rect 564342 4060 564348 4072
rect 527876 4032 564348 4060
rect 527876 4020 527882 4032
rect 564342 4020 564348 4032
rect 564400 4020 564406 4072
rect 264606 3952 264612 4004
rect 264664 3992 264670 4004
rect 285766 3992 285772 4004
rect 264664 3964 285772 3992
rect 264664 3952 264670 3964
rect 285766 3952 285772 3964
rect 285824 3952 285830 4004
rect 328362 3952 328368 4004
rect 328420 3992 328426 4004
rect 345474 3992 345480 4004
rect 328420 3964 345480 3992
rect 328420 3952 328426 3964
rect 345474 3952 345480 3964
rect 345532 3952 345538 4004
rect 355962 3952 355968 4004
rect 356020 3992 356026 4004
rect 400214 3992 400220 4004
rect 356020 3964 400220 3992
rect 356020 3952 356026 3964
rect 400214 3952 400220 3964
rect 400272 3952 400278 4004
rect 416682 3952 416688 4004
rect 416740 3992 416746 4004
rect 517882 3992 517888 4004
rect 416740 3964 517888 3992
rect 416740 3952 416746 3964
rect 517882 3952 517888 3964
rect 517940 3952 517946 4004
rect 529198 3952 529204 4004
rect 529256 3992 529262 4004
rect 571426 3992 571432 4004
rect 529256 3964 571432 3992
rect 529256 3952 529262 3964
rect 571426 3952 571432 3964
rect 571484 3952 571490 4004
rect 261128 3896 262536 3924
rect 204898 3856 204904 3868
rect 180208 3828 181576 3856
rect 181640 3828 204904 3856
rect 180208 3816 180214 3828
rect 25498 3748 25504 3800
rect 25556 3788 25562 3800
rect 31018 3788 31024 3800
rect 25556 3760 31024 3788
rect 25556 3748 25562 3760
rect 31018 3748 31024 3760
rect 31076 3748 31082 3800
rect 34974 3748 34980 3800
rect 35032 3788 35038 3800
rect 166994 3788 167000 3800
rect 35032 3760 167000 3788
rect 35032 3748 35038 3760
rect 166994 3748 167000 3760
rect 167052 3748 167058 3800
rect 176562 3748 176568 3800
rect 176620 3788 176626 3800
rect 176620 3760 181484 3788
rect 176620 3748 176626 3760
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 24118 3720 24124 3732
rect 16080 3692 24124 3720
rect 16080 3680 16086 3692
rect 24118 3680 24124 3692
rect 24176 3680 24182 3732
rect 29086 3680 29092 3732
rect 29144 3720 29150 3732
rect 164234 3720 164240 3732
rect 29144 3692 164240 3720
rect 29144 3680 29150 3692
rect 164234 3680 164240 3692
rect 164292 3680 164298 3732
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 160094 3652 160100 3664
rect 20772 3624 160100 3652
rect 20772 3612 20778 3624
rect 160094 3612 160100 3624
rect 160152 3612 160158 3664
rect 172974 3612 172980 3664
rect 173032 3652 173038 3664
rect 181349 3655 181407 3661
rect 181349 3652 181361 3655
rect 173032 3624 181361 3652
rect 173032 3612 173038 3624
rect 181349 3621 181361 3624
rect 181395 3621 181407 3655
rect 181456 3652 181484 3760
rect 181548 3720 181576 3828
rect 204898 3816 204904 3828
rect 204956 3816 204962 3868
rect 208670 3816 208676 3868
rect 208728 3856 208734 3868
rect 256786 3856 256792 3868
rect 208728 3828 256792 3856
rect 208728 3816 208734 3828
rect 256786 3816 256792 3828
rect 256844 3816 256850 3868
rect 256881 3859 256939 3865
rect 256881 3825 256893 3859
rect 256927 3856 256939 3859
rect 261128 3856 261156 3896
rect 263410 3884 263416 3936
rect 263468 3924 263474 3936
rect 284478 3924 284484 3936
rect 263468 3896 284484 3924
rect 263468 3884 263474 3896
rect 284478 3884 284484 3896
rect 284536 3884 284542 3936
rect 328270 3884 328276 3936
rect 328328 3924 328334 3936
rect 346670 3924 346676 3936
rect 328328 3896 346676 3924
rect 328328 3884 328334 3896
rect 346670 3884 346676 3896
rect 346728 3884 346734 3936
rect 360102 3884 360108 3936
rect 360160 3924 360166 3936
rect 407298 3924 407304 3936
rect 360160 3896 407304 3924
rect 360160 3884 360166 3896
rect 407298 3884 407304 3896
rect 407356 3884 407362 3936
rect 409138 3884 409144 3936
rect 409196 3924 409202 3936
rect 417970 3924 417976 3936
rect 409196 3896 417976 3924
rect 409196 3884 409202 3896
rect 417970 3884 417976 3896
rect 418028 3884 418034 3936
rect 421650 3884 421656 3936
rect 421708 3924 421714 3936
rect 525058 3924 525064 3936
rect 421708 3896 525064 3924
rect 421708 3884 421714 3896
rect 525058 3884 525064 3896
rect 525116 3884 525122 3936
rect 530578 3884 530584 3936
rect 530636 3924 530642 3936
rect 578602 3924 578608 3936
rect 530636 3896 578608 3924
rect 530636 3884 530642 3896
rect 578602 3884 578608 3896
rect 578660 3884 578666 3936
rect 283006 3856 283012 3868
rect 256927 3828 261156 3856
rect 261220 3828 283012 3856
rect 256927 3825 256939 3828
rect 256881 3819 256939 3825
rect 191009 3791 191067 3797
rect 191009 3757 191021 3791
rect 191055 3788 191067 3791
rect 239493 3791 239551 3797
rect 191055 3760 239444 3788
rect 191055 3757 191067 3760
rect 191009 3751 191067 3757
rect 235813 3723 235871 3729
rect 235813 3720 235825 3723
rect 181548 3692 235825 3720
rect 235813 3689 235825 3692
rect 235859 3689 235871 3723
rect 238754 3720 238760 3732
rect 235813 3683 235871 3689
rect 235920 3692 238760 3720
rect 191193 3655 191251 3661
rect 191193 3652 191205 3655
rect 181456 3624 191205 3652
rect 181349 3615 181407 3621
rect 191193 3621 191205 3624
rect 191239 3621 191251 3655
rect 191193 3615 191251 3621
rect 196713 3655 196771 3661
rect 196713 3621 196725 3655
rect 196759 3652 196771 3655
rect 209317 3655 209375 3661
rect 209317 3652 209329 3655
rect 196759 3624 209329 3652
rect 196759 3621 196771 3624
rect 196713 3615 196771 3621
rect 209317 3621 209329 3624
rect 209363 3621 209375 3655
rect 209317 3615 209375 3621
rect 216493 3655 216551 3661
rect 216493 3621 216505 3655
rect 216539 3652 216551 3655
rect 225233 3655 225291 3661
rect 225233 3652 225245 3655
rect 216539 3624 225245 3652
rect 216539 3621 216551 3624
rect 216493 3615 216551 3621
rect 225233 3621 225245 3624
rect 225279 3621 225291 3655
rect 225233 3615 225291 3621
rect 225322 3612 225328 3664
rect 225380 3652 225386 3664
rect 226242 3652 226248 3664
rect 225380 3624 226248 3652
rect 225380 3612 225386 3624
rect 226242 3612 226248 3624
rect 226300 3612 226306 3664
rect 226337 3655 226395 3661
rect 226337 3621 226349 3655
rect 226383 3652 226395 3655
rect 226383 3624 226564 3652
rect 226383 3621 226395 3624
rect 226337 3615 226395 3621
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 13078 3584 13084 3596
rect 6512 3556 13084 3584
rect 6512 3544 6518 3556
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 158714 3584 158720 3596
rect 19576 3556 158720 3584
rect 19576 3544 19582 3556
rect 158714 3544 158720 3556
rect 158772 3544 158778 3596
rect 186225 3587 186283 3593
rect 186225 3553 186237 3587
rect 186271 3584 186283 3587
rect 191101 3587 191159 3593
rect 191101 3584 191113 3587
rect 186271 3556 191113 3584
rect 186271 3553 186283 3556
rect 186225 3547 186283 3553
rect 191101 3553 191113 3556
rect 191147 3553 191159 3587
rect 191101 3547 191159 3553
rect 200761 3587 200819 3593
rect 200761 3553 200773 3587
rect 200807 3584 200819 3587
rect 208765 3587 208823 3593
rect 208765 3584 208777 3587
rect 200807 3556 208777 3584
rect 200807 3553 200819 3556
rect 200761 3547 200819 3553
rect 208765 3553 208777 3556
rect 208811 3553 208823 3587
rect 208765 3547 208823 3553
rect 220081 3587 220139 3593
rect 220081 3553 220093 3587
rect 220127 3584 220139 3587
rect 226536 3584 226564 3624
rect 228910 3612 228916 3664
rect 228968 3652 228974 3664
rect 231210 3652 231216 3664
rect 228968 3624 231216 3652
rect 228968 3612 228974 3624
rect 231210 3612 231216 3624
rect 231268 3612 231274 3664
rect 231302 3612 231308 3664
rect 231360 3652 231366 3664
rect 231762 3652 231768 3664
rect 231360 3624 231768 3652
rect 231360 3612 231366 3624
rect 231762 3612 231768 3624
rect 231820 3612 231826 3664
rect 231857 3655 231915 3661
rect 231857 3621 231869 3655
rect 231903 3652 231915 3655
rect 235920 3652 235948 3692
rect 238754 3680 238760 3692
rect 238812 3680 238818 3732
rect 239416 3720 239444 3760
rect 239493 3757 239505 3791
rect 239539 3788 239551 3791
rect 240226 3788 240232 3800
rect 239539 3760 240232 3788
rect 239539 3757 239551 3760
rect 239493 3751 239551 3757
rect 240226 3748 240232 3760
rect 240284 3748 240290 3800
rect 240778 3748 240784 3800
rect 240836 3788 240842 3800
rect 241422 3788 241428 3800
rect 240836 3760 241428 3788
rect 240836 3748 240842 3760
rect 241422 3748 241428 3760
rect 241480 3748 241486 3800
rect 243170 3748 243176 3800
rect 243228 3788 243234 3800
rect 244182 3788 244188 3800
rect 243228 3760 244188 3788
rect 243228 3748 243234 3760
rect 244182 3748 244188 3760
rect 244240 3748 244246 3800
rect 249150 3748 249156 3800
rect 249208 3788 249214 3800
rect 249702 3788 249708 3800
rect 249208 3760 249708 3788
rect 249208 3748 249214 3760
rect 249702 3748 249708 3760
rect 249760 3748 249766 3800
rect 250346 3748 250352 3800
rect 250404 3788 250410 3800
rect 251082 3788 251088 3800
rect 250404 3760 251088 3788
rect 250404 3748 250410 3760
rect 251082 3748 251088 3760
rect 251140 3748 251146 3800
rect 251450 3748 251456 3800
rect 251508 3788 251514 3800
rect 252462 3788 252468 3800
rect 251508 3760 252468 3788
rect 251508 3748 251514 3760
rect 252462 3748 252468 3760
rect 252520 3748 252526 3800
rect 261018 3748 261024 3800
rect 261076 3788 261082 3800
rect 261220 3788 261248 3828
rect 283006 3816 283012 3828
rect 283064 3816 283070 3868
rect 319990 3816 319996 3868
rect 320048 3856 320054 3868
rect 330018 3856 330024 3868
rect 320048 3828 330024 3856
rect 320048 3816 320054 3828
rect 330018 3816 330024 3828
rect 330076 3816 330082 3868
rect 331122 3816 331128 3868
rect 331180 3856 331186 3868
rect 352558 3856 352564 3868
rect 331180 3828 352564 3856
rect 331180 3816 331186 3828
rect 352558 3816 352564 3828
rect 352616 3816 352622 3868
rect 362862 3816 362868 3868
rect 362920 3856 362926 3868
rect 414474 3856 414480 3868
rect 362920 3828 414480 3856
rect 362920 3816 362926 3828
rect 414474 3816 414480 3828
rect 414532 3816 414538 3868
rect 423582 3816 423588 3868
rect 423640 3856 423646 3868
rect 532234 3856 532240 3868
rect 423640 3828 532240 3856
rect 423640 3816 423646 3828
rect 532234 3816 532240 3828
rect 532292 3816 532298 3868
rect 261076 3760 261248 3788
rect 263597 3791 263655 3797
rect 261076 3748 261082 3760
rect 263597 3757 263609 3791
rect 263643 3788 263655 3791
rect 268473 3791 268531 3797
rect 268473 3788 268485 3791
rect 263643 3760 268485 3788
rect 263643 3757 263655 3760
rect 263597 3751 263655 3757
rect 268473 3757 268485 3760
rect 268519 3757 268531 3791
rect 268473 3751 268531 3757
rect 320082 3748 320088 3800
rect 320140 3788 320146 3800
rect 331214 3788 331220 3800
rect 320140 3760 331220 3788
rect 320140 3748 320146 3760
rect 331214 3748 331220 3760
rect 331272 3748 331278 3800
rect 333882 3748 333888 3800
rect 333940 3788 333946 3800
rect 356146 3788 356152 3800
rect 333940 3760 356152 3788
rect 333940 3748 333946 3760
rect 356146 3748 356152 3760
rect 356204 3748 356210 3800
rect 356698 3748 356704 3800
rect 356756 3788 356762 3800
rect 364518 3788 364524 3800
rect 356756 3760 364524 3788
rect 356756 3748 356762 3760
rect 364518 3748 364524 3760
rect 364576 3748 364582 3800
rect 367002 3748 367008 3800
rect 367060 3788 367066 3800
rect 420362 3788 420368 3800
rect 367060 3760 420368 3788
rect 367060 3748 367066 3760
rect 420362 3748 420368 3760
rect 420420 3748 420426 3800
rect 427722 3748 427728 3800
rect 427780 3788 427786 3800
rect 539318 3788 539324 3800
rect 427780 3760 539324 3788
rect 427780 3748 427786 3760
rect 539318 3748 539324 3760
rect 539376 3748 539382 3800
rect 244458 3720 244464 3732
rect 239416 3692 244464 3720
rect 244458 3680 244464 3692
rect 244516 3680 244522 3732
rect 250438 3720 250444 3732
rect 244568 3692 250444 3720
rect 231903 3624 235948 3652
rect 231903 3621 231915 3624
rect 231857 3615 231915 3621
rect 235994 3612 236000 3664
rect 236052 3652 236058 3664
rect 243538 3652 243544 3664
rect 236052 3624 243544 3652
rect 236052 3612 236058 3624
rect 243538 3612 243544 3624
rect 243596 3612 243602 3664
rect 244277 3655 244335 3661
rect 244277 3621 244289 3655
rect 244323 3652 244335 3655
rect 244568 3652 244596 3692
rect 250438 3680 250444 3692
rect 250496 3680 250502 3732
rect 252646 3680 252652 3732
rect 252704 3720 252710 3732
rect 278866 3720 278872 3732
rect 252704 3692 278872 3720
rect 252704 3680 252710 3692
rect 278866 3680 278872 3692
rect 278924 3680 278930 3732
rect 285950 3680 285956 3732
rect 286008 3720 286014 3732
rect 294598 3720 294604 3732
rect 286008 3692 294604 3720
rect 286008 3680 286014 3692
rect 294598 3680 294604 3692
rect 294656 3680 294662 3732
rect 321370 3680 321376 3732
rect 321428 3720 321434 3732
rect 333606 3720 333612 3732
rect 321428 3692 333612 3720
rect 321428 3680 321434 3692
rect 333606 3680 333612 3692
rect 333664 3680 333670 3732
rect 335262 3680 335268 3732
rect 335320 3720 335326 3732
rect 359734 3720 359740 3732
rect 335320 3692 359740 3720
rect 335320 3680 335326 3692
rect 359734 3680 359740 3692
rect 359792 3680 359798 3732
rect 366910 3680 366916 3732
rect 366968 3720 366974 3732
rect 421558 3720 421564 3732
rect 366968 3692 421564 3720
rect 366968 3680 366974 3692
rect 421558 3680 421564 3692
rect 421616 3680 421622 3732
rect 431862 3680 431868 3732
rect 431920 3720 431926 3732
rect 546494 3720 546500 3732
rect 431920 3692 546500 3720
rect 431920 3680 431926 3692
rect 546494 3680 546500 3692
rect 546552 3680 546558 3732
rect 244323 3624 244596 3652
rect 244323 3621 244335 3624
rect 244277 3615 244335 3621
rect 246758 3612 246764 3664
rect 246816 3652 246822 3664
rect 268381 3655 268439 3661
rect 268381 3652 268393 3655
rect 246816 3624 268393 3652
rect 246816 3612 246822 3624
rect 268381 3621 268393 3624
rect 268427 3621 268439 3655
rect 268381 3615 268439 3621
rect 268473 3655 268531 3661
rect 268473 3621 268485 3655
rect 268519 3652 268531 3655
rect 273254 3652 273260 3664
rect 268519 3624 273260 3652
rect 268519 3621 268531 3624
rect 268473 3615 268531 3621
rect 273254 3612 273260 3624
rect 273312 3612 273318 3664
rect 282454 3612 282460 3664
rect 282512 3652 282518 3664
rect 294138 3652 294144 3664
rect 282512 3624 294144 3652
rect 282512 3612 282518 3624
rect 294138 3612 294144 3624
rect 294196 3612 294202 3664
rect 300302 3612 300308 3664
rect 300360 3652 300366 3664
rect 303614 3652 303620 3664
rect 300360 3624 303620 3652
rect 300360 3612 300366 3624
rect 303614 3612 303620 3624
rect 303672 3612 303678 3664
rect 316770 3612 316776 3664
rect 316828 3652 316834 3664
rect 320450 3652 320456 3664
rect 316828 3624 320456 3652
rect 316828 3612 316834 3624
rect 320450 3612 320456 3624
rect 320508 3612 320514 3664
rect 322750 3612 322756 3664
rect 322808 3652 322814 3664
rect 335906 3652 335912 3664
rect 322808 3624 335912 3652
rect 322808 3612 322814 3624
rect 335906 3612 335912 3624
rect 335964 3612 335970 3664
rect 339402 3612 339408 3664
rect 339460 3652 339466 3664
rect 345753 3655 345811 3661
rect 339460 3624 345704 3652
rect 339460 3612 339466 3624
rect 236270 3584 236276 3596
rect 220127 3556 226472 3584
rect 226536 3556 236276 3584
rect 220127 3553 220139 3556
rect 220081 3547 220139 3553
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 154850 3516 154856 3528
rect 11296 3488 154856 3516
rect 11296 3476 11302 3488
rect 154850 3476 154856 3488
rect 154908 3476 154914 3528
rect 169386 3476 169392 3528
rect 169444 3516 169450 3528
rect 226337 3519 226395 3525
rect 226337 3516 226349 3519
rect 169444 3488 226349 3516
rect 169444 3476 169450 3488
rect 226337 3485 226349 3488
rect 226383 3485 226395 3519
rect 226444 3516 226472 3556
rect 236270 3544 236276 3556
rect 236328 3544 236334 3596
rect 241514 3584 241520 3596
rect 236380 3556 241520 3584
rect 231857 3519 231915 3525
rect 231857 3516 231869 3519
rect 226444 3488 231869 3516
rect 226337 3479 226395 3485
rect 231857 3485 231869 3488
rect 231903 3485 231915 3519
rect 231857 3479 231915 3485
rect 231949 3519 232007 3525
rect 231949 3485 231961 3519
rect 231995 3516 232007 3519
rect 235721 3519 235779 3525
rect 235721 3516 235733 3519
rect 231995 3488 235733 3516
rect 231995 3485 232007 3488
rect 231949 3479 232007 3485
rect 235721 3485 235733 3488
rect 235767 3485 235779 3519
rect 235721 3479 235779 3485
rect 235813 3519 235871 3525
rect 235813 3485 235825 3519
rect 235859 3516 235871 3519
rect 236380 3516 236408 3556
rect 241514 3544 241520 3556
rect 241572 3544 241578 3596
rect 241974 3544 241980 3596
rect 242032 3584 242038 3596
rect 263597 3587 263655 3593
rect 263597 3584 263609 3587
rect 242032 3556 263609 3584
rect 242032 3544 242038 3556
rect 263597 3553 263609 3556
rect 263643 3553 263655 3587
rect 263597 3547 263655 3553
rect 277670 3544 277676 3596
rect 277728 3584 277734 3596
rect 286318 3584 286324 3596
rect 277728 3556 286324 3584
rect 277728 3544 277734 3556
rect 286318 3544 286324 3556
rect 286376 3544 286382 3596
rect 316678 3544 316684 3596
rect 316736 3584 316742 3596
rect 318058 3584 318064 3596
rect 316736 3556 318064 3584
rect 316736 3544 316742 3556
rect 318058 3544 318064 3556
rect 318116 3544 318122 3596
rect 324222 3544 324228 3596
rect 324280 3584 324286 3596
rect 338298 3584 338304 3596
rect 324280 3556 338304 3584
rect 324280 3544 324286 3556
rect 338298 3544 338304 3556
rect 338356 3544 338362 3596
rect 340782 3544 340788 3596
rect 340840 3584 340846 3596
rect 345569 3587 345627 3593
rect 345569 3584 345581 3587
rect 340840 3556 345581 3584
rect 340840 3544 340846 3556
rect 345569 3553 345581 3556
rect 345615 3553 345627 3587
rect 345676 3584 345704 3624
rect 345753 3621 345765 3655
rect 345799 3652 345811 3655
rect 363322 3652 363328 3664
rect 345799 3624 363328 3652
rect 345799 3621 345811 3624
rect 345753 3615 345811 3621
rect 363322 3612 363328 3624
rect 363380 3612 363386 3664
rect 371142 3612 371148 3664
rect 371200 3652 371206 3664
rect 428734 3652 428740 3664
rect 371200 3624 428740 3652
rect 371200 3612 371206 3624
rect 428734 3612 428740 3624
rect 428792 3612 428798 3664
rect 434622 3612 434628 3664
rect 434680 3652 434686 3664
rect 553578 3652 553584 3664
rect 434680 3624 553584 3652
rect 434680 3612 434686 3624
rect 553578 3612 553584 3624
rect 553636 3612 553642 3664
rect 366910 3584 366916 3596
rect 345676 3556 366916 3584
rect 345569 3547 345627 3553
rect 366910 3544 366916 3556
rect 366968 3544 366974 3596
rect 372522 3544 372528 3596
rect 372580 3584 372586 3596
rect 432322 3584 432328 3596
rect 372580 3556 432328 3584
rect 372580 3544 372586 3556
rect 432322 3544 432328 3556
rect 432380 3544 432386 3596
rect 438762 3544 438768 3596
rect 438820 3584 438826 3596
rect 560754 3584 560760 3596
rect 438820 3556 560760 3584
rect 438820 3544 438826 3556
rect 560754 3544 560760 3556
rect 560812 3544 560818 3596
rect 235859 3488 236408 3516
rect 236457 3519 236515 3525
rect 235859 3485 235871 3488
rect 235813 3479 235871 3485
rect 236457 3485 236469 3519
rect 236503 3516 236515 3519
rect 239493 3519 239551 3525
rect 239493 3516 239505 3519
rect 236503 3488 239505 3516
rect 236503 3485 236515 3488
rect 236457 3479 236515 3485
rect 239493 3485 239505 3488
rect 239539 3485 239551 3519
rect 239493 3479 239551 3485
rect 239582 3476 239588 3528
rect 239640 3516 239646 3528
rect 271966 3516 271972 3528
rect 239640 3488 271972 3516
rect 239640 3476 239646 3488
rect 271966 3476 271972 3488
rect 272024 3476 272030 3528
rect 301406 3476 301412 3528
rect 301464 3516 301470 3528
rect 302878 3516 302884 3528
rect 301464 3488 302884 3516
rect 301464 3476 301470 3488
rect 302878 3476 302884 3488
rect 302936 3476 302942 3528
rect 312538 3476 312544 3528
rect 312596 3516 312602 3528
rect 313366 3516 313372 3528
rect 312596 3488 313372 3516
rect 312596 3476 312602 3488
rect 313366 3476 313372 3488
rect 313424 3476 313430 3528
rect 322198 3476 322204 3528
rect 322256 3516 322262 3528
rect 325234 3516 325240 3528
rect 322256 3488 325240 3516
rect 322256 3476 322262 3488
rect 325234 3476 325240 3488
rect 325292 3476 325298 3528
rect 325602 3476 325608 3528
rect 325660 3516 325666 3528
rect 339494 3516 339500 3528
rect 325660 3488 339500 3516
rect 325660 3476 325666 3488
rect 339494 3476 339500 3488
rect 339552 3476 339558 3528
rect 350445 3519 350503 3525
rect 350445 3485 350457 3519
rect 350491 3516 350503 3519
rect 370406 3516 370412 3528
rect 350491 3488 370412 3516
rect 350491 3485 350503 3488
rect 350445 3479 350503 3485
rect 370406 3476 370412 3488
rect 370464 3476 370470 3528
rect 373902 3476 373908 3528
rect 373960 3516 373966 3528
rect 435818 3516 435824 3528
rect 373960 3488 435824 3516
rect 373960 3476 373966 3488
rect 435818 3476 435824 3488
rect 435876 3476 435882 3528
rect 442902 3476 442908 3528
rect 442960 3516 442966 3528
rect 567838 3516 567844 3528
rect 442960 3488 567844 3516
rect 442960 3476 442966 3488
rect 567838 3476 567844 3488
rect 567896 3476 567902 3528
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 154666 3448 154672 3460
rect 10100 3420 154672 3448
rect 10100 3408 10106 3420
rect 154666 3408 154672 3420
rect 154724 3408 154730 3460
rect 165890 3408 165896 3460
rect 165948 3448 165954 3460
rect 234614 3448 234620 3460
rect 165948 3420 234620 3448
rect 165948 3408 165954 3420
rect 234614 3408 234620 3420
rect 234672 3408 234678 3460
rect 234798 3408 234804 3460
rect 234856 3448 234862 3460
rect 268470 3448 268476 3460
rect 234856 3420 268476 3448
rect 234856 3408 234862 3420
rect 268470 3408 268476 3420
rect 268528 3408 268534 3460
rect 270494 3408 270500 3460
rect 270552 3448 270558 3460
rect 270552 3420 276428 3448
rect 270552 3408 270558 3420
rect 32674 3340 32680 3392
rect 32732 3380 32738 3392
rect 35158 3380 35164 3392
rect 32732 3352 35164 3380
rect 32732 3340 32738 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 68278 3340 68284 3392
rect 68336 3380 68342 3392
rect 177298 3380 177304 3392
rect 68336 3352 177304 3380
rect 68336 3340 68342 3352
rect 177298 3340 177304 3352
rect 177356 3340 177362 3392
rect 183738 3340 183744 3392
rect 183796 3380 183802 3392
rect 191009 3383 191067 3389
rect 191009 3380 191021 3383
rect 183796 3352 191021 3380
rect 183796 3340 183802 3352
rect 191009 3349 191021 3352
rect 191055 3349 191067 3383
rect 191009 3343 191067 3349
rect 200390 3340 200396 3392
rect 200448 3380 200454 3392
rect 201402 3380 201408 3392
rect 200448 3352 201408 3380
rect 200448 3340 200454 3352
rect 201402 3340 201408 3352
rect 201460 3340 201466 3392
rect 225233 3383 225291 3389
rect 225233 3349 225245 3383
rect 225279 3380 225291 3383
rect 231949 3383 232007 3389
rect 231949 3380 231961 3383
rect 225279 3352 231961 3380
rect 225279 3349 225291 3352
rect 225233 3343 225291 3349
rect 231949 3349 231961 3352
rect 231995 3349 232007 3383
rect 231949 3343 232007 3349
rect 232041 3383 232099 3389
rect 232041 3349 232053 3383
rect 232087 3380 232099 3383
rect 232087 3352 258580 3380
rect 232087 3349 232099 3352
rect 232041 3343 232099 3349
rect 38562 3272 38568 3324
rect 38620 3312 38626 3324
rect 71038 3312 71044 3324
rect 38620 3284 71044 3312
rect 38620 3272 38626 3284
rect 71038 3272 71044 3284
rect 71096 3272 71102 3324
rect 75454 3272 75460 3324
rect 75512 3312 75518 3324
rect 180058 3312 180064 3324
rect 75512 3284 180064 3312
rect 75512 3272 75518 3284
rect 180058 3272 180064 3284
rect 180116 3272 180122 3324
rect 181349 3315 181407 3321
rect 181349 3281 181361 3315
rect 181395 3312 181407 3315
rect 186225 3315 186283 3321
rect 186225 3312 186237 3315
rect 181395 3284 186237 3312
rect 181395 3281 181407 3284
rect 181349 3275 181407 3281
rect 186225 3281 186237 3284
rect 186271 3281 186283 3315
rect 186225 3275 186283 3281
rect 208765 3315 208823 3321
rect 208765 3281 208777 3315
rect 208811 3312 208823 3315
rect 220081 3315 220139 3321
rect 220081 3312 220093 3315
rect 208811 3284 220093 3312
rect 208811 3281 208823 3284
rect 208765 3275 208823 3281
rect 220081 3281 220093 3284
rect 220127 3281 220139 3315
rect 220081 3275 220139 3281
rect 220173 3315 220231 3321
rect 220173 3281 220185 3315
rect 220219 3312 220231 3315
rect 249061 3315 249119 3321
rect 249061 3312 249073 3315
rect 220219 3284 249073 3312
rect 220219 3281 220231 3284
rect 220173 3275 220231 3281
rect 249061 3281 249073 3284
rect 249107 3281 249119 3315
rect 253753 3315 253811 3321
rect 253753 3312 253765 3315
rect 249061 3275 249119 3281
rect 249168 3284 253765 3312
rect 45738 3204 45744 3256
rect 45796 3244 45802 3256
rect 75178 3244 75184 3256
rect 45796 3216 75184 3244
rect 45796 3204 45802 3216
rect 75178 3204 75184 3216
rect 75236 3204 75242 3256
rect 82630 3204 82636 3256
rect 82688 3244 82694 3256
rect 181438 3244 181444 3256
rect 82688 3216 181444 3244
rect 82688 3204 82694 3216
rect 181438 3204 181444 3216
rect 181496 3204 181502 3256
rect 191101 3247 191159 3253
rect 191101 3213 191113 3247
rect 191147 3244 191159 3247
rect 200761 3247 200819 3253
rect 200761 3244 200773 3247
rect 191147 3216 200773 3244
rect 191147 3213 191159 3216
rect 191101 3207 191159 3213
rect 200761 3213 200773 3216
rect 200807 3213 200819 3247
rect 200761 3207 200819 3213
rect 209866 3204 209872 3256
rect 209924 3244 209930 3256
rect 244277 3247 244335 3253
rect 244277 3244 244289 3247
rect 209924 3216 244289 3244
rect 209924 3204 209930 3216
rect 244277 3213 244289 3216
rect 244323 3213 244335 3247
rect 244277 3207 244335 3213
rect 244366 3204 244372 3256
rect 244424 3244 244430 3256
rect 249168 3244 249196 3284
rect 253753 3281 253765 3284
rect 253799 3281 253811 3315
rect 253753 3275 253811 3281
rect 253842 3272 253848 3324
rect 253900 3312 253906 3324
rect 254670 3312 254676 3324
rect 253900 3284 254676 3312
rect 253900 3272 253906 3284
rect 254670 3272 254676 3284
rect 254728 3272 254734 3324
rect 254765 3315 254823 3321
rect 254765 3281 254777 3315
rect 254811 3312 254823 3315
rect 256881 3315 256939 3321
rect 256881 3312 256893 3315
rect 254811 3284 256893 3312
rect 254811 3281 254823 3284
rect 254765 3275 254823 3281
rect 256881 3281 256893 3284
rect 256927 3281 256939 3315
rect 256881 3275 256939 3281
rect 257430 3272 257436 3324
rect 257488 3312 257494 3324
rect 257982 3312 257988 3324
rect 257488 3284 257988 3312
rect 257488 3272 257494 3284
rect 257982 3272 257988 3284
rect 258040 3272 258046 3324
rect 258552 3312 258580 3352
rect 258626 3340 258632 3392
rect 258684 3380 258690 3392
rect 259362 3380 259368 3392
rect 258684 3352 259368 3380
rect 258684 3340 258690 3352
rect 259362 3340 259368 3352
rect 259420 3340 259426 3392
rect 261570 3380 261576 3392
rect 259472 3352 261576 3380
rect 259472 3312 259500 3352
rect 261570 3340 261576 3352
rect 261628 3340 261634 3392
rect 262214 3340 262220 3392
rect 262272 3380 262278 3392
rect 263502 3380 263508 3392
rect 262272 3352 263508 3380
rect 262272 3340 262278 3352
rect 263502 3340 263508 3352
rect 263560 3340 263566 3392
rect 276400 3380 276428 3420
rect 276474 3408 276480 3460
rect 276532 3448 276538 3460
rect 277302 3448 277308 3460
rect 276532 3420 277308 3448
rect 276532 3408 276538 3420
rect 277302 3408 277308 3420
rect 277360 3408 277366 3460
rect 278866 3408 278872 3460
rect 278924 3448 278930 3460
rect 278924 3420 287376 3448
rect 278924 3408 278930 3420
rect 284938 3380 284944 3392
rect 276400 3352 284944 3380
rect 284938 3340 284944 3352
rect 284996 3340 285002 3392
rect 287348 3380 287376 3420
rect 289538 3408 289544 3460
rect 289596 3448 289602 3460
rect 297358 3448 297364 3460
rect 289596 3420 297364 3448
rect 289596 3408 289602 3420
rect 297358 3408 297364 3420
rect 297416 3408 297422 3460
rect 297910 3408 297916 3460
rect 297968 3448 297974 3460
rect 301590 3448 301596 3460
rect 297968 3420 301596 3448
rect 297968 3408 297974 3420
rect 301590 3408 301596 3420
rect 301648 3408 301654 3460
rect 311802 3408 311808 3460
rect 311860 3448 311866 3460
rect 314562 3448 314568 3460
rect 311860 3420 314568 3448
rect 311860 3408 311866 3420
rect 314562 3408 314568 3420
rect 314620 3408 314626 3460
rect 315942 3408 315948 3460
rect 316000 3448 316006 3460
rect 322842 3448 322848 3460
rect 316000 3420 322848 3448
rect 316000 3408 316006 3420
rect 322842 3408 322848 3420
rect 322900 3408 322906 3460
rect 326982 3408 326988 3460
rect 327040 3448 327046 3460
rect 343082 3448 343088 3460
rect 327040 3420 343088 3448
rect 327040 3408 327046 3420
rect 343082 3408 343088 3420
rect 343140 3408 343146 3460
rect 344922 3408 344928 3460
rect 344980 3448 344986 3460
rect 378778 3448 378784 3460
rect 344980 3420 378784 3448
rect 344980 3408 344986 3420
rect 378778 3408 378784 3420
rect 378836 3408 378842 3460
rect 442994 3448 443000 3460
rect 390756 3420 443000 3448
rect 291838 3380 291844 3392
rect 287348 3352 291844 3380
rect 291838 3340 291844 3352
rect 291896 3340 291902 3392
rect 294322 3340 294328 3392
rect 294380 3380 294386 3392
rect 297450 3380 297456 3392
rect 294380 3352 297456 3380
rect 294380 3340 294386 3352
rect 297450 3340 297456 3352
rect 297508 3340 297514 3392
rect 322934 3340 322940 3392
rect 322992 3380 322998 3392
rect 334710 3380 334716 3392
rect 322992 3352 334716 3380
rect 322992 3340 322998 3352
rect 334710 3340 334716 3352
rect 334768 3340 334774 3392
rect 340138 3340 340144 3392
rect 340196 3380 340202 3392
rect 342717 3383 342775 3389
rect 340196 3352 340828 3380
rect 340196 3340 340202 3352
rect 258552 3284 259500 3312
rect 259822 3272 259828 3324
rect 259880 3312 259886 3324
rect 280798 3312 280804 3324
rect 259880 3284 280804 3312
rect 259880 3272 259886 3284
rect 280798 3272 280804 3284
rect 280856 3272 280862 3324
rect 284754 3272 284760 3324
rect 284812 3312 284818 3324
rect 290458 3312 290464 3324
rect 284812 3284 290464 3312
rect 284812 3272 284818 3284
rect 290458 3272 290464 3284
rect 290516 3272 290522 3324
rect 323578 3272 323584 3324
rect 323636 3312 323642 3324
rect 328822 3312 328828 3324
rect 323636 3284 328828 3312
rect 323636 3272 323642 3284
rect 328822 3272 328828 3284
rect 328880 3272 328886 3324
rect 330478 3272 330484 3324
rect 330536 3312 330542 3324
rect 340690 3312 340696 3324
rect 330536 3284 340696 3312
rect 330536 3272 330542 3284
rect 340690 3272 340696 3284
rect 340748 3272 340754 3324
rect 340800 3312 340828 3352
rect 342717 3349 342729 3383
rect 342763 3380 342775 3383
rect 349062 3380 349068 3392
rect 342763 3352 349068 3380
rect 342763 3349 342775 3352
rect 342717 3343 342775 3349
rect 349062 3340 349068 3352
rect 349120 3340 349126 3392
rect 353754 3380 353760 3392
rect 350368 3352 353760 3380
rect 350258 3312 350264 3324
rect 340800 3284 350264 3312
rect 350258 3272 350264 3284
rect 350316 3272 350322 3324
rect 244424 3216 249196 3244
rect 250533 3247 250591 3253
rect 244424 3204 244430 3216
rect 250533 3213 250545 3247
rect 250579 3244 250591 3247
rect 254578 3244 254584 3256
rect 250579 3216 254584 3244
rect 250579 3213 250591 3216
rect 250533 3207 250591 3213
rect 254578 3204 254584 3216
rect 254636 3204 254642 3256
rect 320818 3204 320824 3256
rect 320876 3244 320882 3256
rect 324038 3244 324044 3256
rect 320876 3216 324044 3244
rect 320876 3204 320882 3216
rect 324038 3204 324044 3216
rect 324096 3204 324102 3256
rect 50522 3136 50528 3188
rect 50580 3176 50586 3188
rect 77938 3176 77944 3188
rect 50580 3148 77944 3176
rect 50580 3136 50586 3148
rect 77938 3136 77944 3148
rect 77996 3136 78002 3188
rect 89714 3136 89720 3188
rect 89772 3176 89778 3188
rect 93118 3176 93124 3188
rect 89772 3148 93124 3176
rect 89772 3136 89778 3148
rect 93118 3136 93124 3148
rect 93176 3136 93182 3188
rect 184198 3176 184204 3188
rect 93228 3148 184204 3176
rect 57606 3068 57612 3120
rect 57664 3108 57670 3120
rect 84838 3108 84844 3120
rect 57664 3080 84844 3108
rect 57664 3068 57670 3080
rect 84838 3068 84844 3080
rect 84896 3068 84902 3120
rect 86126 3068 86132 3120
rect 86184 3108 86190 3120
rect 93228 3108 93256 3148
rect 184198 3136 184204 3148
rect 184256 3136 184262 3188
rect 217042 3136 217048 3188
rect 217100 3176 217106 3188
rect 220173 3179 220231 3185
rect 220173 3176 220185 3179
rect 217100 3148 220185 3176
rect 217100 3136 217106 3148
rect 220173 3145 220185 3148
rect 220219 3145 220231 3179
rect 220173 3139 220231 3145
rect 224126 3136 224132 3188
rect 224184 3176 224190 3188
rect 262858 3176 262864 3188
rect 224184 3148 262864 3176
rect 224184 3136 224190 3148
rect 262858 3136 262864 3148
rect 262916 3136 262922 3188
rect 299106 3136 299112 3188
rect 299164 3176 299170 3188
rect 301498 3176 301504 3188
rect 299164 3148 301504 3176
rect 299164 3136 299170 3148
rect 301498 3136 301504 3148
rect 301556 3136 301562 3188
rect 341518 3136 341524 3188
rect 341576 3176 341582 3188
rect 350368 3176 350396 3352
rect 353754 3340 353760 3352
rect 353812 3340 353818 3392
rect 359458 3340 359464 3392
rect 359516 3380 359522 3392
rect 371602 3380 371608 3392
rect 359516 3352 371608 3380
rect 359516 3340 359522 3352
rect 371602 3340 371608 3352
rect 371660 3340 371666 3392
rect 358078 3272 358084 3324
rect 358136 3312 358142 3324
rect 368014 3312 368020 3324
rect 358136 3284 368020 3312
rect 358136 3272 358142 3284
rect 368014 3272 368020 3284
rect 368072 3272 368078 3324
rect 380158 3272 380164 3324
rect 380216 3312 380222 3324
rect 389450 3312 389456 3324
rect 380216 3284 389456 3312
rect 380216 3272 380222 3284
rect 389450 3272 389456 3284
rect 389508 3272 389514 3324
rect 380250 3204 380256 3256
rect 380308 3244 380314 3256
rect 390756 3244 390784 3420
rect 442994 3408 443000 3420
rect 443052 3408 443058 3460
rect 445662 3408 445668 3460
rect 445720 3448 445726 3460
rect 575014 3448 575020 3460
rect 445720 3420 575020 3448
rect 445720 3408 445726 3420
rect 575014 3408 575020 3420
rect 575072 3408 575078 3460
rect 391198 3340 391204 3392
rect 391256 3380 391262 3392
rect 403710 3380 403716 3392
rect 391256 3352 403716 3380
rect 391256 3340 391262 3352
rect 403710 3340 403716 3352
rect 403768 3340 403774 3392
rect 403802 3340 403808 3392
rect 403860 3380 403866 3392
rect 482278 3380 482284 3392
rect 403860 3352 482284 3380
rect 403860 3340 403866 3352
rect 482278 3340 482284 3352
rect 482336 3340 482342 3392
rect 523678 3340 523684 3392
rect 523736 3380 523742 3392
rect 550082 3380 550088 3392
rect 523736 3352 550088 3380
rect 523736 3340 523742 3352
rect 550082 3340 550088 3352
rect 550140 3340 550146 3392
rect 392578 3272 392584 3324
rect 392636 3312 392642 3324
rect 392636 3284 394096 3312
rect 392636 3272 392642 3284
rect 380308 3216 390784 3244
rect 394068 3244 394096 3284
rect 424318 3272 424324 3324
rect 424376 3312 424382 3324
rect 503622 3312 503628 3324
rect 424376 3284 503628 3312
rect 424376 3272 424382 3284
rect 503622 3272 503628 3284
rect 503680 3272 503686 3324
rect 520918 3272 520924 3324
rect 520976 3312 520982 3324
rect 542906 3312 542912 3324
rect 520976 3284 542912 3312
rect 520976 3272 520982 3284
rect 542906 3272 542912 3284
rect 542964 3272 542970 3324
rect 467926 3244 467932 3256
rect 394068 3216 467932 3244
rect 380308 3204 380314 3216
rect 467926 3204 467932 3216
rect 467984 3204 467990 3256
rect 518158 3204 518164 3256
rect 518216 3244 518222 3256
rect 535730 3244 535736 3256
rect 518216 3216 535736 3244
rect 518216 3204 518222 3216
rect 535730 3204 535736 3216
rect 535788 3204 535794 3256
rect 341576 3148 350396 3176
rect 341576 3136 341582 3148
rect 384298 3136 384304 3188
rect 384356 3176 384362 3188
rect 393038 3176 393044 3188
rect 384356 3148 393044 3176
rect 384356 3136 384362 3148
rect 393038 3136 393044 3148
rect 393096 3136 393102 3188
rect 460842 3176 460848 3188
rect 393976 3148 460848 3176
rect 86184 3080 93256 3108
rect 86184 3068 86190 3080
rect 93302 3068 93308 3120
rect 93360 3108 93366 3120
rect 185578 3108 185584 3120
rect 93360 3080 185584 3108
rect 93360 3068 93366 3080
rect 185578 3068 185584 3080
rect 185636 3068 185642 3120
rect 221734 3068 221740 3120
rect 221792 3108 221798 3120
rect 232041 3111 232099 3117
rect 232041 3108 232053 3111
rect 221792 3080 232053 3108
rect 221792 3068 221798 3080
rect 232041 3077 232053 3080
rect 232087 3077 232099 3111
rect 232041 3071 232099 3077
rect 232133 3111 232191 3117
rect 232133 3077 232145 3111
rect 232179 3108 232191 3111
rect 266446 3108 266452 3120
rect 232179 3080 266452 3108
rect 232179 3077 232191 3080
rect 232133 3071 232191 3077
rect 266446 3068 266452 3080
rect 266504 3068 266510 3120
rect 266998 3068 267004 3120
rect 267056 3108 267062 3120
rect 267642 3108 267648 3120
rect 267056 3080 267648 3108
rect 267056 3068 267062 3080
rect 267642 3068 267648 3080
rect 267700 3068 267706 3120
rect 345569 3111 345627 3117
rect 345569 3077 345581 3111
rect 345615 3108 345627 3111
rect 350445 3111 350503 3117
rect 350445 3108 350457 3111
rect 345615 3080 350457 3108
rect 345615 3077 345627 3080
rect 345569 3071 345627 3077
rect 350445 3077 350457 3080
rect 350491 3077 350503 3111
rect 350445 3071 350503 3077
rect 377398 3068 377404 3120
rect 377456 3108 377462 3120
rect 382366 3108 382372 3120
rect 377456 3080 382372 3108
rect 377456 3068 377462 3080
rect 382366 3068 382372 3080
rect 382424 3068 382430 3120
rect 388530 3068 388536 3120
rect 388588 3108 388594 3120
rect 393976 3108 394004 3148
rect 460842 3136 460848 3148
rect 460900 3136 460906 3188
rect 514018 3136 514024 3188
rect 514076 3176 514082 3188
rect 528646 3176 528652 3188
rect 514076 3148 528652 3176
rect 514076 3136 514082 3148
rect 528646 3136 528652 3148
rect 528704 3136 528710 3188
rect 450170 3108 450176 3120
rect 388588 3080 394004 3108
rect 396736 3080 450176 3108
rect 388588 3068 388594 3080
rect 46934 3000 46940 3052
rect 46992 3040 46998 3052
rect 95878 3040 95884 3052
rect 46992 3012 95884 3040
rect 46992 3000 46998 3012
rect 95878 3000 95884 3012
rect 95936 3000 95942 3052
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 98638 3040 98644 3052
rect 96948 3012 98644 3040
rect 96948 3000 96954 3012
rect 98638 3000 98644 3012
rect 98696 3000 98702 3052
rect 103974 3000 103980 3052
rect 104032 3040 104038 3052
rect 104802 3040 104808 3052
rect 104032 3012 104808 3040
rect 104032 3000 104038 3012
rect 104802 3000 104808 3012
rect 104860 3000 104866 3052
rect 111150 3000 111156 3052
rect 111208 3040 111214 3052
rect 111702 3040 111708 3052
rect 111208 3012 111708 3040
rect 111208 3000 111214 3012
rect 111702 3000 111708 3012
rect 111760 3000 111766 3052
rect 186958 3040 186964 3052
rect 111812 3012 186964 3040
rect 71866 2932 71872 2984
rect 71924 2972 71930 2984
rect 86218 2972 86224 2984
rect 71924 2944 86224 2972
rect 71924 2932 71930 2944
rect 86218 2932 86224 2944
rect 86276 2932 86282 2984
rect 100478 2932 100484 2984
rect 100536 2972 100542 2984
rect 111812 2972 111840 3012
rect 186958 3000 186964 3012
rect 187016 3000 187022 3052
rect 193214 3000 193220 3052
rect 193272 3040 193278 3052
rect 197998 3040 198004 3052
rect 193272 3012 198004 3040
rect 193272 3000 193278 3012
rect 197998 3000 198004 3012
rect 198056 3000 198062 3052
rect 206278 3000 206284 3052
rect 206336 3040 206342 3052
rect 226978 3040 226984 3052
rect 206336 3012 226984 3040
rect 206336 3000 206342 3012
rect 226978 3000 226984 3012
rect 227036 3000 227042 3052
rect 230106 3000 230112 3052
rect 230164 3040 230170 3052
rect 267826 3040 267832 3052
rect 230164 3012 267832 3040
rect 230164 3000 230170 3012
rect 267826 3000 267832 3012
rect 267884 3000 267890 3052
rect 275278 3000 275284 3052
rect 275336 3040 275342 3052
rect 275922 3040 275928 3052
rect 275336 3012 275928 3040
rect 275336 3000 275342 3012
rect 275922 3000 275928 3012
rect 275980 3000 275986 3052
rect 287146 3000 287152 3052
rect 287204 3040 287210 3052
rect 288250 3040 288256 3052
rect 287204 3012 288256 3040
rect 287204 3000 287210 3012
rect 288250 3000 288256 3012
rect 288308 3000 288314 3052
rect 293126 3000 293132 3052
rect 293184 3040 293190 3052
rect 298830 3040 298836 3052
rect 293184 3012 298836 3040
rect 293184 3000 293190 3012
rect 298830 3000 298836 3012
rect 298888 3000 298894 3052
rect 338758 3000 338764 3052
rect 338816 3040 338822 3052
rect 341886 3040 341892 3052
rect 338816 3012 341892 3040
rect 338816 3000 338822 3012
rect 341886 3000 341892 3012
rect 341944 3000 341950 3052
rect 388438 3000 388444 3052
rect 388496 3040 388502 3052
rect 396626 3040 396632 3052
rect 388496 3012 396632 3040
rect 388496 3000 388502 3012
rect 396626 3000 396632 3012
rect 396684 3000 396690 3052
rect 188614 2972 188620 2984
rect 100536 2944 111840 2972
rect 111904 2944 188620 2972
rect 100536 2932 100542 2944
rect 64782 2864 64788 2916
rect 64840 2904 64846 2916
rect 106918 2904 106924 2916
rect 64840 2876 106924 2904
rect 64840 2864 64846 2876
rect 106918 2864 106924 2876
rect 106976 2864 106982 2916
rect 79042 2796 79048 2848
rect 79100 2836 79106 2848
rect 88978 2836 88984 2848
rect 79100 2808 88984 2836
rect 79100 2796 79106 2808
rect 88978 2796 88984 2808
rect 89036 2796 89042 2848
rect 107562 2796 107568 2848
rect 107620 2836 107626 2848
rect 111904 2836 111932 2944
rect 188614 2932 188620 2944
rect 188672 2932 188678 2984
rect 226518 2932 226524 2984
rect 226576 2972 226582 2984
rect 264974 2972 264980 2984
rect 226576 2944 264980 2972
rect 226576 2932 226582 2944
rect 264974 2932 264980 2944
rect 265032 2932 265038 2984
rect 283650 2932 283656 2984
rect 283708 2972 283714 2984
rect 284202 2972 284208 2984
rect 283708 2944 284208 2972
rect 283708 2932 283714 2944
rect 284202 2932 284208 2944
rect 284260 2932 284266 2984
rect 384390 2932 384396 2984
rect 384448 2972 384454 2984
rect 386417 2975 386475 2981
rect 386417 2972 386429 2975
rect 384448 2944 386429 2972
rect 384448 2932 384454 2944
rect 386417 2941 386429 2944
rect 386463 2941 386475 2975
rect 386417 2935 386475 2941
rect 114738 2864 114744 2916
rect 114796 2904 114802 2916
rect 115842 2904 115848 2916
rect 114796 2876 115848 2904
rect 114796 2864 114802 2876
rect 115842 2864 115848 2876
rect 115900 2864 115906 2916
rect 121822 2864 121828 2916
rect 121880 2904 121886 2916
rect 122742 2904 122748 2916
rect 121880 2876 122748 2904
rect 121880 2864 121886 2876
rect 122742 2864 122748 2876
rect 122800 2864 122806 2916
rect 125410 2864 125416 2916
rect 125468 2904 125474 2916
rect 127621 2907 127679 2913
rect 125468 2876 127572 2904
rect 125468 2864 125474 2876
rect 107620 2808 111932 2836
rect 107620 2796 107626 2808
rect 118234 2796 118240 2848
rect 118292 2836 118298 2848
rect 127437 2839 127495 2845
rect 127437 2836 127449 2839
rect 118292 2808 127449 2836
rect 118292 2796 118298 2808
rect 127437 2805 127449 2808
rect 127483 2805 127495 2839
rect 127437 2799 127495 2805
rect 127544 2768 127572 2876
rect 127621 2873 127633 2907
rect 127667 2904 127679 2907
rect 188338 2904 188344 2916
rect 127667 2876 188344 2904
rect 127667 2873 127679 2876
rect 127621 2867 127679 2873
rect 188338 2864 188344 2876
rect 188396 2864 188402 2916
rect 227714 2864 227720 2916
rect 227772 2904 227778 2916
rect 232133 2907 232191 2913
rect 232133 2904 232145 2907
rect 227772 2876 232145 2904
rect 227772 2864 227778 2876
rect 232133 2873 232145 2876
rect 232179 2873 232191 2907
rect 232133 2867 232191 2873
rect 232498 2864 232504 2916
rect 232556 2904 232562 2916
rect 269206 2904 269212 2916
rect 232556 2876 269212 2904
rect 232556 2864 232562 2876
rect 269206 2864 269212 2876
rect 269264 2864 269270 2916
rect 296714 2864 296720 2916
rect 296772 2904 296778 2916
rect 302418 2904 302424 2916
rect 296772 2876 302424 2904
rect 296772 2864 296778 2876
rect 302418 2864 302424 2876
rect 302476 2864 302482 2916
rect 395985 2907 396043 2913
rect 395985 2873 395997 2907
rect 396031 2904 396043 2907
rect 396736 2904 396764 3080
rect 450170 3068 450176 3080
rect 450228 3068 450234 3120
rect 411898 3000 411904 3052
rect 411956 3040 411962 3052
rect 425146 3040 425152 3052
rect 411956 3012 425152 3040
rect 411956 3000 411962 3012
rect 425146 3000 425152 3012
rect 425204 3000 425210 3052
rect 435358 3000 435364 3052
rect 435416 3040 435422 3052
rect 496538 3040 496544 3052
rect 435416 3012 496544 3040
rect 435416 3000 435422 3012
rect 496538 3000 496544 3012
rect 496596 3000 496602 3052
rect 502978 3000 502984 3052
rect 503036 3040 503042 3052
rect 507210 3040 507216 3052
rect 503036 3012 507216 3040
rect 503036 3000 503042 3012
rect 507210 3000 507216 3012
rect 507268 3000 507274 3052
rect 421466 2932 421472 2984
rect 421524 2972 421530 2984
rect 481082 2972 481088 2984
rect 421524 2944 481088 2972
rect 421524 2932 421530 2944
rect 481082 2932 481088 2944
rect 481140 2932 481146 2984
rect 396031 2876 396764 2904
rect 396031 2873 396043 2876
rect 395985 2867 396043 2873
rect 420178 2864 420184 2916
rect 420236 2904 420242 2916
rect 477494 2904 477500 2916
rect 420236 2876 477500 2904
rect 420236 2864 420242 2876
rect 477494 2864 477500 2876
rect 477552 2864 477558 2916
rect 191098 2836 191104 2848
rect 127728 2808 191104 2836
rect 127728 2768 127756 2808
rect 191098 2796 191104 2808
rect 191156 2796 191162 2848
rect 218146 2796 218152 2848
rect 218204 2836 218210 2848
rect 249061 2839 249119 2845
rect 218204 2808 249012 2836
rect 218204 2796 218210 2808
rect 127544 2740 127756 2768
rect 248984 2768 249012 2808
rect 249061 2805 249073 2839
rect 249107 2836 249119 2839
rect 257338 2836 257344 2848
rect 249107 2808 257344 2836
rect 249107 2805 249119 2808
rect 249061 2799 249119 2805
rect 257338 2796 257344 2808
rect 257396 2796 257402 2848
rect 290737 2839 290795 2845
rect 290737 2805 290749 2839
rect 290783 2836 290795 2839
rect 291102 2836 291108 2848
rect 290783 2808 291108 2836
rect 290783 2805 290795 2808
rect 290737 2799 290795 2805
rect 291102 2796 291108 2808
rect 291160 2796 291166 2848
rect 431218 2796 431224 2848
rect 431276 2836 431282 2848
rect 489362 2836 489368 2848
rect 431276 2808 489368 2836
rect 431276 2796 431282 2808
rect 489362 2796 489368 2808
rect 489420 2796 489426 2848
rect 250533 2771 250591 2777
rect 250533 2768 250545 2771
rect 248984 2740 250545 2768
rect 250533 2737 250545 2740
rect 250579 2737 250591 2771
rect 250533 2731 250591 2737
rect 386417 2771 386475 2777
rect 386417 2737 386429 2771
rect 386463 2768 386475 2771
rect 395985 2771 396043 2777
rect 395985 2768 395997 2771
rect 386463 2740 395997 2768
rect 386463 2737 386475 2740
rect 386417 2731 386475 2737
rect 395985 2737 395997 2740
rect 396031 2737 396043 2771
rect 395985 2731 396043 2737
rect 373997 2703 374055 2709
rect 373997 2669 374009 2703
rect 374043 2700 374055 2703
rect 374270 2700 374276 2712
rect 374043 2672 374276 2700
rect 374043 2669 374055 2672
rect 373997 2663 374055 2669
rect 374270 2660 374276 2672
rect 374328 2660 374334 2712
rect 374086 1504 374092 1556
rect 374144 1544 374150 1556
rect 375190 1544 375196 1556
rect 374144 1516 375196 1544
rect 374144 1504 374150 1516
rect 375190 1504 375196 1516
rect 375248 1504 375254 1556
rect 238386 552 238392 604
rect 238444 592 238450 604
rect 238570 592 238576 604
rect 238444 564 238576 592
rect 238444 552 238450 564
rect 238570 552 238576 564
rect 238628 552 238634 604
rect 256234 552 256240 604
rect 256292 592 256298 604
rect 256602 592 256608 604
rect 256292 564 256608 592
rect 256292 552 256298 564
rect 256602 552 256608 564
rect 256660 552 256666 604
rect 281258 552 281264 604
rect 281316 592 281322 604
rect 281442 592 281448 604
rect 281316 564 281448 592
rect 281316 552 281322 564
rect 281442 552 281448 564
rect 281500 552 281506 604
rect 290734 592 290740 604
rect 290695 564 290740 592
rect 290734 552 290740 564
rect 290792 552 290798 604
rect 325786 552 325792 604
rect 325844 592 325850 604
rect 326430 592 326436 604
rect 325844 564 326436 592
rect 325844 552 325850 564
rect 326430 552 326436 564
rect 326488 552 326494 604
rect 350810 552 350816 604
rect 350868 592 350874 604
rect 351362 592 351368 604
rect 350868 564 351368 592
rect 350868 552 350874 564
rect 351362 552 351368 564
rect 351420 552 351426 604
rect 361850 552 361856 604
rect 361908 592 361914 604
rect 362126 592 362132 604
rect 361908 564 362132 592
rect 361908 552 361914 564
rect 362126 552 362132 564
rect 362184 552 362190 604
rect 368474 552 368480 604
rect 368532 592 368538 604
rect 369210 592 369216 604
rect 368532 564 369216 592
rect 368532 552 368538 564
rect 369210 552 369216 564
rect 369268 552 369274 604
rect 372614 552 372620 604
rect 372672 592 372678 604
rect 372798 592 372804 604
rect 372672 564 372804 592
rect 372672 552 372678 564
rect 372798 552 372804 564
rect 372856 552 372862 604
rect 373994 592 374000 604
rect 373955 564 374000 592
rect 373994 552 374000 564
rect 374052 552 374058 604
rect 379698 552 379704 604
rect 379756 592 379762 604
rect 379974 592 379980 604
rect 379756 564 379980 592
rect 379756 552 379762 564
rect 379974 552 379980 564
rect 380032 552 380038 604
rect 382458 552 382464 604
rect 382516 592 382522 604
rect 383562 592 383568 604
rect 382516 564 383568 592
rect 382516 552 382522 564
rect 383562 552 383568 564
rect 383620 552 383626 604
rect 439038 552 439044 604
rect 439096 592 439102 604
rect 439406 592 439412 604
rect 439096 564 439412 592
rect 439096 552 439102 564
rect 439406 552 439412 564
rect 439464 552 439470 604
rect 445754 552 445760 604
rect 445812 592 445818 604
rect 446582 592 446588 604
rect 445812 564 446588 592
rect 445812 552 445818 564
rect 446582 552 446588 564
rect 446640 552 446646 604
rect 470594 552 470600 604
rect 470652 592 470658 604
rect 471514 592 471520 604
rect 470652 564 471520 592
rect 470652 552 470658 564
rect 471514 552 471520 564
rect 471572 552 471578 604
rect 473354 552 473360 604
rect 473412 592 473418 604
rect 473906 592 473912 604
rect 473412 564 473912 592
rect 473412 552 473418 564
rect 473906 552 473912 564
rect 473964 552 473970 604
rect 477586 552 477592 604
rect 477644 592 477650 604
rect 478690 592 478696 604
rect 477644 564 478696 592
rect 477644 552 477650 564
rect 478690 552 478696 564
rect 478748 552 478754 604
rect 499574 552 499580 604
rect 499632 592 499638 604
rect 500126 592 500132 604
rect 499632 564 500132 592
rect 499632 552 499638 564
rect 500126 552 500132 564
rect 500184 552 500190 604
<< via1 >>
rect 154120 700952 154172 701004
rect 318800 700952 318852 701004
rect 137836 700884 137888 700936
rect 316040 700884 316092 700936
rect 278688 700816 278740 700868
rect 462320 700816 462372 700868
rect 281448 700748 281500 700800
rect 478512 700748 478564 700800
rect 105452 700680 105504 700732
rect 321560 700680 321612 700732
rect 89168 700612 89220 700664
rect 327080 700612 327132 700664
rect 72976 700544 73028 700596
rect 324320 700544 324372 700596
rect 270408 700476 270460 700528
rect 527180 700476 527232 700528
rect 273168 700408 273220 700460
rect 543464 700408 543516 700460
rect 40500 700340 40552 700392
rect 328460 700340 328512 700392
rect 24308 700272 24360 700324
rect 333980 700272 334032 700324
rect 170312 700204 170364 700256
rect 313280 700204 313332 700256
rect 288348 700136 288400 700188
rect 413652 700136 413704 700188
rect 286968 700068 287020 700120
rect 397460 700068 397512 700120
rect 202788 700000 202840 700052
rect 307760 700000 307812 700052
rect 218980 699932 219032 699984
rect 310520 699932 310572 699984
rect 296628 699864 296680 699916
rect 348792 699864 348844 699916
rect 293868 699796 293920 699848
rect 332508 699796 332560 699848
rect 267648 699728 267700 699780
rect 300860 699728 300912 699780
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 283840 699660 283892 699712
rect 303620 699660 303672 699712
rect 263508 696940 263560 696992
rect 580172 696940 580224 696992
rect 299664 688576 299716 688628
rect 300124 688576 300176 688628
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 266268 685856 266320 685908
rect 580172 685856 580224 685908
rect 299572 684428 299624 684480
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 336740 681708 336792 681760
rect 364340 676175 364392 676184
rect 364340 676141 364349 676175
rect 364349 676141 364383 676175
rect 364383 676141 364392 676175
rect 364340 676132 364392 676141
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 260748 673480 260800 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 342260 667904 342312 667956
rect 299940 666544 299992 666596
rect 364432 666544 364484 666596
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 339500 652740 339552 652792
rect 255228 650020 255280 650072
rect 580172 650020 580224 650072
rect 299664 647232 299716 647284
rect 299756 647232 299808 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 299664 640364 299716 640416
rect 299756 640364 299808 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 257988 638936 258040 638988
rect 580172 638936 580224 638988
rect 364340 634788 364392 634840
rect 364524 634788 364576 634840
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 299572 630640 299624 630692
rect 299756 630640 299808 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 252468 626560 252520 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 345020 623772 345072 623824
rect 364340 615476 364392 615528
rect 364524 615476 364576 615528
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 3424 609968 3476 610020
rect 349160 609968 349212 610020
rect 299664 608583 299716 608592
rect 299664 608549 299673 608583
rect 299673 608549 299707 608583
rect 299707 608549 299716 608583
rect 299664 608540 299716 608549
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 246948 603100 247000 603152
rect 580172 603100 580224 603152
rect 299848 601672 299900 601724
rect 429568 601672 429620 601724
rect 559288 601672 559340 601724
rect 299848 598927 299900 598936
rect 299848 598893 299857 598927
rect 299857 598893 299891 598927
rect 299891 598893 299900 598927
rect 299848 598884 299900 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 364340 596164 364392 596216
rect 364524 596164 364576 596216
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 347780 594804 347832 594856
rect 249708 592016 249760 592068
rect 580172 592016 580224 592068
rect 299940 589296 299992 589348
rect 429660 589296 429712 589348
rect 559380 589296 559432 589348
rect 364156 589228 364208 589280
rect 364432 589228 364484 589280
rect 493876 589228 493928 589280
rect 494152 589228 494204 589280
rect 299940 582428 299992 582480
rect 429660 582428 429712 582480
rect 559380 582428 559432 582480
rect 299848 582292 299900 582344
rect 429568 582292 429620 582344
rect 559288 582292 559340 582344
rect 245568 579640 245620 579692
rect 580172 579640 580224 579692
rect 3424 567196 3476 567248
rect 351920 567196 351972 567248
rect 299572 563116 299624 563168
rect 429292 563116 429344 563168
rect 559012 563116 559064 563168
rect 299572 562980 299624 563032
rect 429292 562980 429344 563032
rect 559012 562980 559064 563032
rect 299572 560235 299624 560244
rect 299572 560201 299581 560235
rect 299581 560201 299615 560235
rect 299615 560201 299624 560235
rect 299572 560192 299624 560201
rect 559012 560235 559064 560244
rect 559012 560201 559021 560235
rect 559021 560201 559055 560235
rect 559055 560201 559064 560235
rect 559012 560192 559064 560201
rect 240048 556180 240100 556232
rect 580172 556180 580224 556232
rect 429200 553435 429252 553444
rect 429200 553401 429209 553435
rect 429209 553401 429243 553435
rect 429243 553401 429252 553435
rect 429200 553392 429252 553401
rect 3424 552100 3476 552152
rect 357440 552100 357492 552152
rect 156420 552032 156472 552084
rect 577504 552032 577556 552084
rect 299664 550604 299716 550656
rect 429200 550647 429252 550656
rect 429200 550613 429209 550647
rect 429209 550613 429243 550647
rect 429243 550613 429252 550647
rect 429200 550604 429252 550613
rect 559104 550604 559156 550656
rect 235908 550128 235960 550180
rect 306380 550128 306432 550180
rect 290924 550060 290976 550112
rect 364340 550060 364392 550112
rect 283104 549992 283156 550044
rect 429200 549992 429252 550044
rect 275376 549924 275428 549976
rect 494060 549924 494112 549976
rect 267648 549856 267700 549908
rect 559104 549856 559156 549908
rect 298652 549244 298704 549296
rect 299572 549244 299624 549296
rect 226248 549176 226300 549228
rect 449532 549176 449584 549228
rect 223672 549108 223724 549160
rect 449624 549108 449676 549160
rect 218428 549040 218480 549092
rect 449348 549040 449400 549092
rect 2964 548972 3016 549024
rect 355508 548972 355560 549024
rect 4712 548904 4764 548956
rect 365904 548904 365956 548956
rect 5264 548836 5316 548888
rect 371056 548836 371108 548888
rect 3056 548768 3108 548820
rect 368480 548768 368532 548820
rect 5356 548700 5408 548752
rect 373632 548700 373684 548752
rect 3148 548632 3200 548684
rect 376208 548632 376260 548684
rect 5172 548564 5224 548616
rect 378784 548564 378836 548616
rect 6368 548496 6420 548548
rect 381360 548496 381412 548548
rect 3240 548428 3292 548480
rect 384028 548428 384080 548480
rect 6276 548360 6328 548412
rect 389180 548360 389232 548412
rect 4068 548292 4120 548344
rect 391756 548292 391808 548344
rect 5080 548224 5132 548276
rect 394332 548224 394384 548276
rect 6184 548156 6236 548208
rect 396908 548156 396960 548208
rect 10324 548088 10376 548140
rect 404636 548088 404688 548140
rect 3976 548020 4028 548072
rect 399484 548020 399536 548072
rect 19984 547952 20036 548004
rect 420184 547952 420236 548004
rect 4896 547884 4948 547936
rect 409880 547884 409932 547936
rect 149704 545504 149756 545556
rect 401692 545504 401744 545556
rect 184756 545436 184808 545488
rect 449256 545436 449308 545488
rect 177488 545368 177540 545420
rect 449164 545368 449216 545420
rect 242072 545300 242124 545352
rect 580172 545300 580224 545352
rect 5448 545232 5500 545284
rect 363052 545232 363104 545284
rect 192852 545164 192904 545216
rect 580724 545164 580776 545216
rect 187608 545096 187660 545148
rect 580540 545096 580592 545148
rect 236920 544892 236972 544944
rect 449072 544892 449124 544944
rect 229008 544824 229060 544876
rect 449716 544824 449768 544876
rect 216128 544756 216180 544808
rect 449440 544756 449492 544808
rect 161848 544731 161900 544740
rect 161848 544697 161857 544731
rect 161857 544697 161891 544731
rect 161891 544697 161900 544731
rect 161848 544688 161900 544697
rect 164056 544731 164108 544740
rect 164056 544697 164065 544731
rect 164065 544697 164099 544731
rect 164099 544697 164108 544731
rect 164056 544688 164108 544697
rect 169576 544731 169628 544740
rect 169576 544697 169585 544731
rect 169585 544697 169619 544731
rect 169619 544697 169628 544731
rect 169576 544688 169628 544697
rect 172152 544731 172204 544740
rect 172152 544697 172161 544731
rect 172161 544697 172195 544731
rect 172195 544697 172204 544731
rect 172152 544688 172204 544697
rect 174912 544731 174964 544740
rect 174912 544697 174921 544731
rect 174921 544697 174955 544731
rect 174955 544697 174964 544731
rect 174912 544688 174964 544697
rect 180064 544731 180116 544740
rect 180064 544697 180073 544731
rect 180073 544697 180107 544731
rect 180107 544697 180116 544731
rect 180064 544688 180116 544697
rect 182640 544731 182692 544740
rect 182640 544697 182649 544731
rect 182649 544697 182683 544731
rect 182683 544697 182692 544731
rect 182640 544688 182692 544697
rect 195520 544731 195572 544740
rect 195520 544697 195529 544731
rect 195529 544697 195563 544731
rect 195563 544697 195572 544731
rect 195520 544688 195572 544697
rect 200672 544731 200724 544740
rect 200672 544697 200681 544731
rect 200681 544697 200715 544731
rect 200715 544697 200724 544731
rect 200672 544688 200724 544697
rect 234344 544688 234396 544740
rect 580080 544688 580132 544740
rect 6460 544620 6512 544672
rect 360476 544620 360528 544672
rect 412180 544663 412232 544672
rect 412180 544629 412189 544663
rect 412189 544629 412223 544663
rect 412223 544629 412232 544663
rect 412180 544620 412232 544629
rect 417332 544663 417384 544672
rect 417332 544629 417341 544663
rect 417341 544629 417375 544663
rect 417375 544629 417384 544663
rect 417332 544620 417384 544629
rect 427820 544663 427872 544672
rect 427820 544629 427829 544663
rect 427829 544629 427863 544663
rect 427863 544629 427872 544663
rect 432788 544663 432840 544672
rect 427820 544620 427872 544629
rect 432788 544629 432797 544663
rect 432797 544629 432831 544663
rect 432831 544629 432840 544663
rect 432788 544620 432840 544629
rect 438216 544663 438268 544672
rect 438216 544629 438225 544663
rect 438225 544629 438259 544663
rect 438259 544629 438268 544663
rect 438216 544620 438268 544629
rect 443092 544663 443144 544672
rect 443092 544629 443101 544663
rect 443101 544629 443135 544663
rect 443135 544629 443144 544663
rect 443092 544620 443144 544629
rect 580908 544552 580960 544604
rect 580632 544484 580684 544536
rect 578056 544416 578108 544468
rect 580448 544348 580500 544400
rect 577964 544280 578016 544332
rect 4988 544212 5040 544264
rect 580356 544144 580408 544196
rect 577872 544076 577924 544128
rect 3884 544008 3936 544060
rect 577688 543940 577740 543992
rect 3792 543872 3844 543924
rect 3608 543804 3660 543856
rect 3424 543736 3476 543788
rect 3516 542784 3568 542836
rect 580264 542852 580316 542904
rect 449072 534012 449124 534064
rect 579896 534012 579948 534064
rect 449808 510552 449860 510604
rect 579896 510552 579948 510604
rect 2964 509940 3016 509992
rect 6460 509940 6512 509992
rect 2780 495524 2832 495576
rect 4712 495524 4764 495576
rect 449716 487092 449768 487144
rect 580080 487092 580132 487144
rect 2780 481108 2832 481160
rect 5448 481108 5500 481160
rect 449624 463632 449676 463684
rect 580080 463632 580132 463684
rect 449532 452548 449584 452600
rect 580080 452548 580132 452600
rect 2780 438540 2832 438592
rect 5356 438540 5408 438592
rect 2780 424804 2832 424856
rect 5264 424804 5316 424856
rect 449440 416712 449492 416764
rect 580080 416712 580132 416764
rect 449348 405628 449400 405680
rect 580080 405628 580132 405680
rect 2964 380604 3016 380656
rect 6368 380604 6420 380656
rect 2780 366936 2832 366988
rect 5172 366936 5224 366988
rect 3148 324096 3200 324148
rect 6276 324096 6328 324148
rect 3148 280100 3200 280152
rect 6184 280100 6236 280152
rect 2780 266160 2832 266212
rect 5080 266160 5132 266212
rect 346952 243176 347004 243228
rect 368940 243040 368992 243092
rect 369768 243040 369820 243092
rect 186872 242972 186924 243024
rect 71044 242836 71096 242888
rect 169760 242836 169812 242888
rect 42064 242768 42116 242820
rect 103428 242768 103480 242820
rect 190552 242836 190604 242888
rect 199660 242836 199712 242888
rect 210700 242836 210752 242888
rect 211896 242836 211948 242888
rect 254124 242836 254176 242888
rect 257988 242836 258040 242888
rect 183376 242768 183428 242820
rect 86224 242700 86276 242752
rect 260196 242768 260248 242820
rect 267556 242768 267608 242820
rect 286508 242836 286560 242888
rect 312728 242836 312780 242888
rect 316040 242836 316092 242888
rect 341432 242836 341484 242888
rect 346308 242836 346360 242888
rect 282184 242768 282236 242820
rect 284944 242768 284996 242820
rect 288900 242768 288952 242820
rect 331680 242768 331732 242820
rect 341524 242768 341576 242820
rect 345112 242768 345164 242820
rect 367744 242904 367796 242956
rect 414480 242904 414532 242956
rect 377404 242836 377456 242888
rect 398104 242836 398156 242888
rect 399484 242836 399536 242888
rect 485780 242836 485832 242888
rect 364708 242768 364760 242820
rect 370136 242768 370188 242820
rect 371148 242768 371200 242820
rect 375656 242768 375708 242820
rect 439044 242768 439096 242820
rect 443460 242768 443512 242820
rect 199384 242700 199436 242752
rect 245568 242700 245620 242752
rect 245660 242700 245712 242752
rect 280344 242700 280396 242752
rect 294788 242700 294840 242752
rect 296812 242700 296864 242752
rect 314568 242700 314620 242752
rect 316776 242700 316828 242752
rect 329840 242700 329892 242752
rect 340144 242700 340196 242752
rect 343272 242700 343324 242752
rect 88984 242632 89036 242684
rect 183468 242632 183520 242684
rect 188344 242632 188396 242684
rect 211804 242632 211856 242684
rect 258356 242632 258408 242684
rect 259368 242632 259420 242684
rect 282828 242632 282880 242684
rect 286324 242632 286376 242684
rect 292580 242632 292632 242684
rect 313924 242632 313976 242684
rect 319076 242632 319128 242684
rect 328644 242632 328696 242684
rect 342076 242632 342128 242684
rect 378140 242700 378192 242752
rect 379428 242700 379480 242752
rect 93124 242564 93176 242616
rect 196072 242564 196124 242616
rect 208308 242564 208360 242616
rect 256516 242564 256568 242616
rect 113180 242496 113232 242548
rect 122748 242496 122800 242548
rect 170404 242496 170456 242548
rect 180064 242496 180116 242548
rect 188712 242496 188764 242548
rect 203616 242496 203668 242548
rect 252284 242496 252336 242548
rect 254584 242496 254636 242548
rect 262036 242564 262088 242616
rect 266268 242564 266320 242616
rect 284668 242564 284720 242616
rect 313372 242564 313424 242616
rect 316684 242564 316736 242616
rect 325608 242564 325660 242616
rect 338764 242564 338816 242616
rect 351828 242632 351880 242684
rect 367100 242632 367152 242684
rect 367652 242632 367704 242684
rect 376944 242632 376996 242684
rect 405004 242700 405056 242752
rect 435364 242700 435416 242752
rect 436192 242700 436244 242752
rect 525064 242700 525116 242752
rect 385684 242632 385736 242684
rect 403164 242632 403216 242684
rect 492680 242632 492732 242684
rect 379704 242564 379756 242616
rect 401324 242564 401376 242616
rect 425152 242564 425204 242616
rect 432512 242564 432564 242616
rect 523684 242564 523736 242616
rect 256700 242496 256752 242548
rect 281540 242496 281592 242548
rect 288256 242496 288308 242548
rect 297456 242496 297508 242548
rect 333520 242496 333572 242548
rect 35164 242428 35216 242480
rect 166724 242428 166776 242480
rect 176108 242428 176160 242480
rect 181352 242428 181404 242480
rect 184204 242428 184256 242480
rect 194232 242428 194284 242480
rect 198280 242428 198332 242480
rect 247408 242428 247460 242480
rect 248328 242428 248380 242480
rect 277308 242428 277360 242480
rect 277400 242428 277452 242480
rect 291936 242428 291988 242480
rect 292488 242428 292540 242480
rect 299940 242428 299992 242480
rect 347964 242428 348016 242480
rect 349988 242428 350040 242480
rect 357348 242496 357400 242548
rect 367100 242496 367152 242548
rect 367468 242496 367520 242548
rect 391204 242496 391256 242548
rect 397644 242496 397696 242548
rect 403624 242496 403676 242548
rect 502984 242496 503036 242548
rect 359464 242428 359516 242480
rect 31024 242360 31076 242412
rect 163044 242360 163096 242412
rect 187148 242360 187200 242412
rect 201500 242360 201552 242412
rect 204168 242360 204220 242412
rect 254676 242360 254728 242412
rect 255228 242360 255280 242412
rect 280988 242360 281040 242412
rect 288348 242360 288400 242412
rect 298100 242360 298152 242412
rect 326804 242360 326856 242412
rect 342904 242360 342956 242412
rect 24124 242292 24176 242344
rect 158168 242292 158220 242344
rect 185584 242292 185636 242344
rect 197912 242292 197964 242344
rect 198188 242292 198240 242344
rect 249708 242292 249760 242344
rect 277952 242292 278004 242344
rect 284208 242292 284260 242344
rect 295616 242292 295668 242344
rect 315212 242292 315264 242344
rect 321652 242292 321704 242344
rect 324964 242292 325016 242344
rect 330484 242292 330536 242344
rect 336004 242292 336056 242344
rect 355232 242292 355284 242344
rect 355508 242292 355560 242344
rect 361856 242428 361908 242480
rect 395344 242428 395396 242480
rect 397092 242428 397144 242480
rect 421564 242428 421616 242480
rect 431224 242428 431276 242480
rect 518164 242428 518216 242480
rect 369584 242360 369636 242412
rect 382464 242360 382516 242412
rect 389732 242360 389784 242412
rect 395252 242360 395304 242412
rect 420184 242360 420236 242412
rect 421472 242360 421524 242412
rect 514024 242360 514076 242412
rect 361028 242292 361080 242344
rect 409144 242292 409196 242344
rect 410524 242292 410576 242344
rect 416044 242292 416096 242344
rect 416688 242292 416740 242344
rect 507124 242292 507176 242344
rect 28264 242224 28316 242276
rect 162400 242224 162452 242276
rect 163504 242224 163556 242276
rect 200948 242224 201000 242276
rect 201408 242224 201460 242276
rect 252836 242224 252888 242276
rect 254676 242224 254728 242276
rect 281448 242224 281500 242276
rect 294420 242224 294472 242276
rect 317604 242224 317656 242276
rect 325792 242224 325844 242276
rect 337752 242224 337804 242276
rect 357440 242224 357492 242276
rect 368388 242224 368440 242276
rect 411260 242224 411312 242276
rect 411720 242224 411772 242276
rect 412548 242224 412600 242276
rect 422944 242224 422996 242276
rect 428832 242224 428884 242276
rect 520924 242224 520976 242276
rect 17224 242156 17276 242208
rect 157524 242156 157576 242208
rect 181628 242156 181680 242208
rect 192392 242156 192444 242208
rect 197268 242156 197320 242208
rect 249156 242156 249208 242208
rect 252468 242156 252520 242208
rect 279148 242156 279200 242208
rect 280068 242156 280120 242208
rect 293776 242156 293828 242208
rect 318248 242156 318300 242208
rect 327264 242156 327316 242208
rect 332324 242156 332376 242208
rect 348792 242156 348844 242208
rect 388628 242156 388680 242208
rect 392216 242156 392268 242208
rect 406844 242156 406896 242208
rect 499580 242156 499632 242208
rect 98644 242088 98696 242140
rect 103428 242088 103480 242140
rect 104808 242088 104860 242140
rect 203340 242088 203392 242140
rect 215208 242088 215260 242140
rect 226248 242088 226300 242140
rect 265716 242088 265768 242140
rect 267648 242088 267700 242140
rect 287060 242088 287112 242140
rect 343916 242088 343968 242140
rect 77944 242020 77996 242072
rect 175832 242020 175884 242072
rect 202144 242020 202196 242072
rect 243728 242020 243780 242072
rect 244188 242020 244240 242072
rect 268476 242020 268528 242072
rect 275468 242020 275520 242072
rect 275928 242020 275980 242072
rect 291384 242020 291436 242072
rect 342720 242020 342772 242072
rect 374092 242020 374144 242072
rect 374276 242088 374328 242140
rect 384304 242088 384356 242140
rect 384856 242088 384908 242140
rect 408684 242088 408736 242140
rect 412916 242088 412968 242140
rect 413928 242088 413980 242140
rect 415400 242088 415452 242140
rect 416504 242088 416556 242140
rect 417240 242088 417292 242140
rect 418068 242088 418120 242140
rect 419632 242088 419684 242140
rect 421656 242088 421708 242140
rect 440424 242088 440476 242140
rect 441528 242088 441580 242140
rect 441712 242088 441764 242140
rect 443000 242088 443052 242140
rect 445760 242088 445812 242140
rect 447140 242088 447192 242140
rect 376024 242020 376076 242072
rect 379336 242020 379388 242072
rect 442724 242020 442776 242072
rect 442908 242020 442960 242072
rect 444748 242020 444800 242072
rect 445576 242020 445628 242072
rect 445944 242020 445996 242072
rect 447048 242020 447100 242072
rect 447784 242020 447836 242072
rect 448428 242020 448480 242072
rect 448980 242020 449032 242072
rect 449808 242020 449860 242072
rect 529204 242088 529256 242140
rect 530584 242020 530636 242072
rect 75184 241952 75236 242004
rect 173440 241952 173492 242004
rect 177304 241952 177356 242004
rect 185032 241952 185084 242004
rect 200764 241952 200816 242004
rect 228456 241952 228508 242004
rect 231768 241952 231820 242004
rect 268752 241952 268804 242004
rect 269028 241952 269080 242004
rect 287704 241952 287756 242004
rect 372804 241952 372856 242004
rect 375104 241952 375156 242004
rect 394056 241952 394108 242004
rect 395804 241952 395856 242004
rect 477592 241952 477644 242004
rect 111708 241884 111760 241936
rect 207020 241884 207072 241936
rect 232504 241884 232556 241936
rect 261576 241884 261628 241936
rect 263876 241884 263928 241936
rect 271788 241884 271840 241936
rect 289544 241884 289596 241936
rect 335360 241884 335412 241936
rect 350816 241884 350868 241936
rect 380164 241884 380216 241936
rect 84844 241816 84896 241868
rect 179512 241816 179564 241868
rect 188436 241816 188488 241868
rect 204812 241816 204864 241868
rect 204904 241816 204956 241868
rect 241244 241816 241296 241868
rect 241428 241816 241480 241868
rect 273628 241816 273680 241868
rect 278504 241816 278556 241868
rect 339592 241816 339644 241868
rect 368480 241816 368532 241868
rect 371424 241816 371476 241868
rect 391388 241884 391440 241936
rect 393412 241884 393464 241936
rect 473360 241884 473412 241936
rect 388536 241816 388588 241868
rect 115848 241748 115900 241800
rect 208860 241748 208912 241800
rect 272432 241748 272484 241800
rect 273168 241748 273220 241800
rect 290096 241748 290148 241800
rect 291108 241748 291160 241800
rect 299296 241748 299348 241800
rect 334164 241748 334216 241800
rect 122748 241680 122800 241732
rect 212540 241680 212592 241732
rect 226984 241680 227036 241732
rect 255872 241680 255924 241732
rect 257344 241680 257396 241732
rect 261392 241680 261444 241732
rect 262864 241680 262916 241732
rect 265072 241680 265124 241732
rect 270408 241680 270460 241732
rect 287980 241680 288032 241732
rect 318892 241680 318944 241732
rect 323584 241680 323636 241732
rect 330760 241680 330812 241732
rect 345664 241680 345716 241732
rect 349436 241680 349488 241732
rect 350448 241680 350500 241732
rect 365812 241748 365864 241800
rect 367376 241748 367428 241800
rect 368388 241748 368440 241800
rect 369124 241748 369176 241800
rect 357440 241680 357492 241732
rect 384488 241748 384540 241800
rect 95884 241612 95936 241664
rect 174084 241612 174136 241664
rect 174544 241612 174596 241664
rect 177672 241612 177724 241664
rect 191104 241612 191156 241664
rect 214380 241612 214432 241664
rect 243544 241612 243596 241664
rect 271236 241612 271288 241664
rect 106924 241544 106976 241596
rect 183192 241544 183244 241596
rect 250996 241544 251048 241596
rect 251088 241544 251140 241596
rect 274548 241612 274600 241664
rect 290740 241612 290792 241664
rect 298744 241612 298796 241664
rect 301780 241612 301832 241664
rect 302884 241612 302936 241664
rect 304816 241612 304868 241664
rect 317052 241612 317104 241664
rect 322204 241612 322256 241664
rect 337200 241612 337252 241664
rect 276112 241544 276164 241596
rect 290464 241544 290516 241596
rect 296260 241544 296312 241596
rect 297456 241544 297508 241596
rect 301136 241544 301188 241596
rect 301504 241544 301556 241596
rect 303620 241544 303672 241596
rect 304264 241544 304316 241596
rect 305368 241544 305420 241596
rect 310336 241544 310388 241596
rect 311900 241544 311952 241596
rect 312176 241544 312228 241596
rect 314844 241544 314896 241596
rect 316408 241544 316460 241596
rect 320824 241544 320876 241596
rect 329196 241544 329248 241596
rect 333244 241544 333296 241596
rect 336556 241544 336608 241596
rect 338856 241544 338908 241596
rect 339040 241612 339092 241664
rect 358084 241612 358136 241664
rect 356704 241544 356756 241596
rect 357072 241544 357124 241596
rect 360384 241612 360436 241664
rect 369124 241612 369176 241664
rect 377496 241612 377548 241664
rect 380256 241612 380308 241664
rect 375564 241544 375616 241596
rect 391296 241680 391348 241732
rect 470600 241816 470652 241868
rect 466460 241748 466512 241800
rect 463700 241680 463752 241732
rect 383016 241612 383068 241664
rect 113180 241476 113232 241528
rect 122656 241476 122708 241528
rect 160836 241476 160888 241528
rect 208216 241476 208268 241528
rect 238668 241519 238720 241528
rect 238668 241485 238677 241519
rect 238677 241485 238711 241519
rect 238711 241485 238720 241519
rect 238668 241476 238720 241485
rect 250444 241476 250496 241528
rect 257712 241476 257764 241528
rect 261484 241476 261536 241528
rect 263232 241476 263284 241528
rect 263508 241476 263560 241528
rect 274824 241476 274876 241528
rect 280804 241476 280856 241528
rect 283380 241476 283432 241528
rect 291844 241476 291896 241528
rect 293224 241476 293276 241528
rect 297364 241476 297416 241528
rect 298652 241476 298704 241528
rect 298836 241476 298888 241528
rect 300492 241476 300544 241528
rect 301596 241476 301648 241528
rect 302976 241476 303028 241528
rect 304908 241476 304960 241528
rect 306012 241476 306064 241528
rect 307208 241476 307260 241528
rect 309692 241476 309744 241528
rect 310428 241476 310480 241528
rect 310888 241476 310940 241528
rect 312544 241476 312596 241528
rect 320640 241476 320692 241528
rect 321468 241476 321520 241528
rect 321928 241476 321980 241528
rect 322848 241476 322900 241528
rect 323124 241476 323176 241528
rect 324136 241476 324188 241528
rect 324320 241476 324372 241528
rect 325608 241476 325660 241528
rect 326160 241476 326212 241528
rect 326988 241476 327040 241528
rect 327448 241476 327500 241528
rect 328368 241476 328420 241528
rect 332876 241476 332928 241528
rect 333888 241476 333940 241528
rect 338396 241476 338448 241528
rect 339408 241476 339460 241528
rect 340880 241476 340932 241528
rect 198280 241451 198332 241460
rect 198280 241417 198289 241451
rect 198289 241417 198323 241451
rect 198323 241417 198332 241451
rect 198280 241408 198332 241417
rect 303804 241451 303856 241460
rect 303804 241417 303813 241451
rect 303813 241417 303847 241451
rect 303847 241417 303856 241451
rect 303804 241408 303856 241417
rect 306288 241408 306340 241460
rect 348148 241476 348200 241528
rect 349068 241476 349120 241528
rect 352472 241476 352524 241528
rect 353208 241476 353260 241528
rect 354772 241476 354824 241528
rect 354864 241476 354916 241528
rect 355876 241476 355928 241528
rect 356152 241476 356204 241528
rect 357348 241476 357400 241528
rect 357992 241476 358044 241528
rect 358728 241476 358780 241528
rect 359188 241476 359240 241528
rect 360108 241476 360160 241528
rect 361580 241476 361632 241528
rect 362776 241476 362828 241528
rect 363420 241476 363472 241528
rect 364248 241476 364300 241528
rect 365904 241476 365956 241528
rect 367008 241476 367060 241528
rect 356336 241408 356388 241460
rect 372620 241476 372672 241528
rect 373816 241476 373868 241528
rect 374460 241476 374512 241528
rect 375288 241476 375340 241528
rect 381176 241544 381228 241596
rect 384396 241544 384448 241596
rect 386696 241544 386748 241596
rect 388536 241544 388588 241596
rect 390376 241612 390428 241664
rect 392584 241612 392636 241664
rect 456800 241612 456852 241664
rect 452660 241544 452712 241596
rect 379980 241476 380032 241528
rect 380808 241476 380860 241528
rect 382372 241476 382424 241528
rect 383568 241476 383620 241528
rect 383660 241476 383712 241528
rect 384948 241476 385000 241528
rect 385408 241476 385460 241528
rect 386328 241476 386380 241528
rect 387892 241476 387944 241528
rect 388996 241476 389048 241528
rect 390928 241476 390980 241528
rect 391848 241476 391900 241528
rect 393964 241476 394016 241528
rect 395436 241476 395488 241528
rect 396448 241476 396500 241528
rect 397368 241476 397420 241528
rect 398932 241476 398984 241528
rect 400128 241476 400180 241528
rect 400772 241476 400824 241528
rect 401508 241476 401560 241528
rect 401968 241476 402020 241528
rect 402796 241476 402848 241528
rect 404360 241476 404412 241528
rect 405648 241476 405700 241528
rect 406200 241476 406252 241528
rect 407028 241476 407080 241528
rect 407488 241476 407540 241528
rect 408316 241476 408368 241528
rect 409880 241476 409932 241528
rect 411168 241476 411220 241528
rect 411260 241476 411312 241528
rect 411904 241476 411956 241528
rect 412364 241476 412416 241528
rect 418436 241476 418488 241528
rect 419448 241476 419500 241528
rect 420920 241476 420972 241528
rect 422116 241476 422168 241528
rect 423864 241476 423916 241528
rect 423956 241476 424008 241528
rect 424784 241476 424836 241528
rect 425796 241476 425848 241528
rect 426348 241476 426400 241528
rect 426992 241476 427044 241528
rect 427728 241476 427780 241528
rect 428188 241476 428240 241528
rect 429108 241476 429160 241528
rect 429476 241476 429528 241528
rect 430488 241476 430540 241528
rect 430672 241476 430724 241528
rect 423220 241451 423272 241460
rect 423220 241417 423229 241451
rect 423229 241417 423263 241451
rect 423263 241417 423272 241451
rect 423220 241408 423272 241417
rect 431684 241476 431736 241528
rect 431868 241476 431920 241528
rect 433708 241476 433760 241528
rect 434536 241476 434588 241528
rect 434904 241476 434956 241528
rect 436008 241476 436060 241528
rect 436744 241476 436796 241528
rect 437388 241476 437440 241528
rect 438032 241476 438084 241528
rect 438768 241476 438820 241528
rect 439228 241476 439280 241528
rect 440148 241476 440200 241528
rect 440240 241476 440292 241528
rect 527824 241476 527876 241528
rect 431868 241340 431920 241392
rect 237748 239368 237800 239420
rect 149060 239300 149112 239352
rect 149980 239300 150032 239352
rect 150716 239300 150768 239352
rect 151176 239300 151228 239352
rect 158720 239300 158772 239352
rect 159732 239300 159784 239352
rect 164332 239300 164384 239352
rect 165252 239300 165304 239352
rect 167000 239300 167052 239352
rect 167644 239300 167696 239352
rect 171140 239300 171192 239352
rect 171876 239300 171928 239352
rect 190552 239300 190604 239352
rect 191380 239300 191432 239352
rect 196072 239300 196124 239352
rect 196900 239300 196952 239352
rect 201592 239300 201644 239352
rect 202420 239300 202472 239352
rect 212632 239300 212684 239352
rect 213460 239300 213512 239352
rect 215300 239300 215352 239352
rect 215852 239300 215904 239352
rect 220820 239300 220872 239352
rect 221372 239300 221424 239352
rect 222200 239300 222252 239352
rect 223212 239300 223264 239352
rect 227812 239300 227864 239352
rect 228732 239300 228784 239352
rect 230480 239300 230532 239352
rect 231124 239300 231176 239352
rect 231860 239300 231912 239352
rect 232412 239300 232464 239352
rect 233332 239300 233384 239352
rect 234252 239300 234304 239352
rect 241520 239300 241572 239352
rect 242164 239300 242216 239352
rect 244372 239300 244424 239352
rect 244556 239300 244608 239352
rect 247224 239300 247276 239352
rect 247776 239300 247828 239352
rect 249892 239300 249944 239352
rect 250076 239300 250128 239352
rect 270500 239300 270552 239352
rect 271512 239300 271564 239352
rect 272064 239300 272116 239352
rect 272800 239300 272852 239352
rect 276020 239300 276072 239352
rect 276480 239300 276532 239352
rect 423312 239232 423364 239284
rect 269212 238688 269264 238740
rect 269580 238688 269632 238740
rect 3056 237328 3108 237380
rect 10324 237328 10376 237380
rect 222476 236648 222528 236700
rect 222660 236648 222712 236700
rect 223764 236648 223816 236700
rect 224408 236648 224460 236700
rect 233240 236648 233292 236700
rect 233516 236648 233568 236700
rect 194968 235943 195020 235952
rect 194968 235909 194977 235943
rect 194977 235909 195011 235943
rect 195011 235909 195020 235943
rect 194968 235900 195020 235909
rect 265164 234812 265216 234864
rect 265992 234812 266044 234864
rect 164240 234744 164292 234796
rect 164516 234744 164568 234796
rect 245936 234608 245988 234660
rect 246488 234608 246540 234660
rect 351000 234608 351052 234660
rect 351736 234608 351788 234660
rect 403624 234676 403676 234728
rect 270500 234540 270552 234592
rect 270684 234540 270736 234592
rect 403532 234540 403584 234592
rect 185032 231888 185084 231940
rect 185860 231888 185912 231940
rect 163044 231820 163096 231872
rect 163228 231820 163280 231872
rect 174084 231820 174136 231872
rect 174360 231820 174412 231872
rect 179604 231820 179656 231872
rect 179880 231820 179932 231872
rect 185124 231820 185176 231872
rect 185400 231820 185452 231872
rect 190644 231820 190696 231872
rect 190736 231820 190788 231872
rect 196164 231820 196216 231872
rect 196256 231820 196308 231872
rect 198280 231863 198332 231872
rect 198280 231829 198289 231863
rect 198289 231829 198323 231863
rect 198323 231829 198332 231863
rect 198280 231820 198332 231829
rect 208492 231820 208544 231872
rect 209136 231820 209188 231872
rect 211252 231820 211304 231872
rect 211528 231820 211580 231872
rect 225052 231820 225104 231872
rect 225696 231820 225748 231872
rect 226616 231820 226668 231872
rect 226800 231820 226852 231872
rect 229376 231820 229428 231872
rect 229836 231820 229888 231872
rect 234896 231820 234948 231872
rect 235448 231820 235500 231872
rect 236368 231820 236420 231872
rect 236552 231820 236604 231872
rect 237656 231863 237708 231872
rect 237656 231829 237665 231863
rect 237665 231829 237699 231863
rect 237699 231829 237708 231863
rect 237656 231820 237708 231829
rect 239128 231820 239180 231872
rect 239680 231820 239732 231872
rect 303896 231820 303948 231872
rect 393780 231820 393832 231872
rect 393964 231820 394016 231872
rect 403532 231795 403584 231804
rect 403532 231761 403541 231795
rect 403541 231761 403575 231795
rect 403575 231761 403584 231795
rect 403532 231752 403584 231761
rect 207112 230460 207164 230512
rect 207204 230460 207256 230512
rect 238484 230460 238536 230512
rect 238668 230460 238720 230512
rect 248144 230460 248196 230512
rect 248236 230460 248288 230512
rect 374276 230460 374328 230512
rect 374460 230460 374512 230512
rect 449256 229032 449308 229084
rect 580172 229032 580224 229084
rect 169944 227035 169996 227044
rect 169944 227001 169953 227035
rect 169953 227001 169987 227035
rect 169987 227001 169996 227035
rect 169944 226992 169996 227001
rect 194968 226355 195020 226364
rect 194968 226321 194977 226355
rect 194977 226321 195011 226355
rect 195011 226321 195020 226355
rect 194968 226312 195020 226321
rect 154856 224995 154908 225004
rect 154856 224961 154865 224995
rect 154865 224961 154899 224995
rect 154899 224961 154908 224995
rect 154856 224952 154908 224961
rect 156144 224995 156196 225004
rect 156144 224961 156153 224995
rect 156153 224961 156187 224995
rect 156187 224961 156196 224995
rect 156144 224952 156196 224961
rect 168656 225020 168708 225072
rect 191932 224995 191984 225004
rect 191932 224961 191941 224995
rect 191941 224961 191975 224995
rect 191975 224961 191984 224995
rect 191932 224952 191984 224961
rect 198280 224952 198332 225004
rect 168564 224884 168616 224936
rect 218428 224952 218480 225004
rect 245936 225020 245988 225072
rect 278964 225020 279016 225072
rect 247224 224952 247276 225004
rect 252652 224952 252704 225004
rect 252836 224952 252888 225004
rect 307852 224952 307904 225004
rect 308036 224952 308088 225004
rect 346124 224952 346176 225004
rect 346308 224952 346360 225004
rect 357164 224952 357216 225004
rect 357348 224952 357400 225004
rect 423220 224995 423272 225004
rect 423220 224961 423229 224995
rect 423229 224961 423263 224995
rect 423263 224961 423272 224995
rect 423220 224952 423272 224961
rect 218244 224884 218296 224936
rect 245844 224884 245896 224936
rect 198372 224816 198424 224868
rect 247316 224816 247368 224868
rect 3332 223524 3384 223576
rect 149704 223524 149756 223576
rect 424692 222232 424744 222284
rect 424784 222232 424836 222284
rect 154856 222207 154908 222216
rect 154856 222173 154865 222207
rect 154865 222173 154899 222207
rect 154899 222173 154908 222207
rect 154856 222164 154908 222173
rect 156144 222207 156196 222216
rect 156144 222173 156153 222207
rect 156153 222173 156187 222207
rect 156187 222173 156196 222207
rect 156144 222164 156196 222173
rect 170036 222164 170088 222216
rect 179604 222164 179656 222216
rect 179788 222164 179840 222216
rect 185124 222164 185176 222216
rect 185308 222164 185360 222216
rect 191932 222207 191984 222216
rect 191932 222173 191941 222207
rect 191941 222173 191975 222207
rect 191975 222173 191984 222207
rect 191932 222164 191984 222173
rect 196164 222164 196216 222216
rect 196348 222164 196400 222216
rect 205824 222164 205876 222216
rect 205916 222164 205968 222216
rect 223856 222207 223908 222216
rect 223856 222173 223865 222207
rect 223865 222173 223899 222207
rect 223899 222173 223908 222207
rect 223856 222164 223908 222173
rect 225144 222207 225196 222216
rect 225144 222173 225153 222207
rect 225153 222173 225187 222207
rect 225187 222173 225196 222207
rect 225144 222164 225196 222173
rect 265164 222164 265216 222216
rect 265348 222164 265400 222216
rect 278872 222207 278924 222216
rect 278872 222173 278881 222207
rect 278881 222173 278915 222207
rect 278915 222173 278924 222207
rect 278872 222164 278924 222173
rect 403716 222164 403768 222216
rect 423220 222207 423272 222216
rect 423220 222173 423229 222207
rect 423229 222173 423263 222207
rect 423263 222173 423272 222207
rect 423220 222164 423272 222173
rect 168564 222096 168616 222148
rect 245844 222096 245896 222148
rect 424692 222139 424744 222148
rect 424692 222105 424701 222139
rect 424701 222105 424735 222139
rect 424735 222105 424744 222139
rect 424692 222096 424744 222105
rect 168656 221960 168708 222012
rect 245936 221960 245988 222012
rect 216772 220872 216824 220924
rect 216864 220872 216916 220924
rect 223856 220847 223908 220856
rect 223856 220813 223865 220847
rect 223865 220813 223899 220847
rect 223899 220813 223908 220847
rect 223856 220804 223908 220813
rect 225144 220847 225196 220856
rect 225144 220813 225153 220847
rect 225153 220813 225187 220847
rect 225187 220813 225196 220847
rect 225144 220804 225196 220813
rect 247960 220804 248012 220856
rect 248328 220804 248380 220856
rect 379060 220804 379112 220856
rect 379244 220804 379296 220856
rect 384580 220804 384632 220856
rect 384856 220804 384908 220856
rect 216772 220736 216824 220788
rect 216956 220736 217008 220788
rect 218244 220736 218296 220788
rect 218336 220736 218388 220788
rect 379152 220736 379204 220788
rect 379336 220736 379388 220788
rect 216956 219419 217008 219428
rect 216956 219385 216965 219419
rect 216965 219385 216999 219419
rect 216999 219385 217008 219419
rect 216956 219376 217008 219385
rect 218336 219376 218388 219428
rect 194508 216588 194560 216640
rect 194968 216588 195020 216640
rect 179604 215364 179656 215416
rect 222568 215364 222620 215416
rect 265164 215364 265216 215416
rect 270684 215364 270736 215416
rect 423220 215364 423272 215416
rect 278872 215296 278924 215348
rect 178224 215271 178276 215280
rect 178224 215237 178233 215271
rect 178233 215237 178267 215271
rect 178267 215237 178276 215271
rect 178224 215228 178276 215237
rect 222476 215228 222528 215280
rect 258172 215228 258224 215280
rect 258356 215228 258408 215280
rect 263784 215271 263836 215280
rect 263784 215237 263793 215271
rect 263793 215237 263827 215271
rect 263827 215237 263836 215271
rect 263784 215228 263836 215237
rect 272064 215271 272116 215280
rect 272064 215237 272073 215271
rect 272073 215237 272107 215271
rect 272107 215237 272116 215271
rect 272064 215228 272116 215237
rect 423220 215228 423272 215280
rect 278872 215160 278924 215212
rect 403532 215160 403584 215212
rect 403716 215160 403768 215212
rect 154764 212508 154816 212560
rect 154856 212508 154908 212560
rect 170036 212508 170088 212560
rect 170128 212508 170180 212560
rect 178224 212551 178276 212560
rect 178224 212517 178233 212551
rect 178233 212517 178267 212551
rect 178267 212517 178276 212551
rect 178224 212508 178276 212517
rect 179512 212551 179564 212560
rect 179512 212517 179521 212551
rect 179521 212517 179555 212551
rect 179555 212517 179564 212551
rect 179512 212508 179564 212517
rect 185124 212508 185176 212560
rect 185216 212508 185268 212560
rect 190736 212508 190788 212560
rect 190920 212508 190972 212560
rect 191748 212508 191800 212560
rect 192024 212508 192076 212560
rect 247316 212508 247368 212560
rect 247408 212508 247460 212560
rect 263784 212551 263836 212560
rect 263784 212517 263793 212551
rect 263793 212517 263827 212551
rect 263827 212517 263836 212551
rect 263784 212508 263836 212517
rect 265072 212551 265124 212560
rect 265072 212517 265081 212551
rect 265081 212517 265115 212551
rect 265115 212517 265124 212551
rect 265072 212508 265124 212517
rect 270592 212551 270644 212560
rect 270592 212517 270601 212551
rect 270601 212517 270635 212551
rect 270635 212517 270644 212551
rect 270592 212508 270644 212517
rect 272064 212551 272116 212560
rect 272064 212517 272073 212551
rect 272073 212517 272107 212551
rect 272107 212517 272116 212551
rect 272064 212508 272116 212517
rect 424784 212508 424836 212560
rect 196256 211216 196308 211268
rect 196348 211216 196400 211268
rect 248144 211148 248196 211200
rect 248236 211148 248288 211200
rect 198188 211080 198240 211132
rect 198372 211080 198424 211132
rect 216956 211123 217008 211132
rect 216956 211089 216965 211123
rect 216965 211089 216999 211123
rect 216999 211089 217008 211123
rect 216956 211080 217008 211089
rect 219532 211080 219584 211132
rect 379152 211080 379204 211132
rect 379244 211080 379296 211132
rect 384672 211123 384724 211132
rect 384672 211089 384681 211123
rect 384681 211089 384715 211123
rect 384715 211089 384724 211123
rect 384672 211080 384724 211089
rect 219624 211012 219676 211064
rect 150808 209788 150860 209840
rect 150900 209788 150952 209840
rect 214012 209831 214064 209840
rect 214012 209797 214021 209831
rect 214021 209797 214055 209831
rect 214055 209797 214064 209831
rect 214012 209788 214064 209797
rect 205916 206252 205968 206304
rect 206100 206252 206152 206304
rect 238484 206252 238536 206304
rect 238668 206252 238720 206304
rect 192024 205708 192076 205760
rect 150808 205640 150860 205692
rect 162860 205640 162912 205692
rect 163044 205640 163096 205692
rect 173900 205640 173952 205692
rect 174084 205640 174136 205692
rect 252652 205640 252704 205692
rect 252836 205640 252888 205692
rect 284300 205640 284352 205692
rect 284484 205640 284536 205692
rect 307852 205640 307904 205692
rect 308036 205640 308088 205692
rect 346124 205640 346176 205692
rect 346308 205640 346360 205692
rect 357164 205640 357216 205692
rect 357348 205640 357400 205692
rect 423220 205683 423272 205692
rect 423220 205649 423229 205683
rect 423229 205649 423263 205683
rect 423263 205649 423272 205683
rect 423220 205640 423272 205649
rect 192024 205572 192076 205624
rect 218244 205615 218296 205624
rect 218244 205581 218253 205615
rect 218253 205581 218287 205615
rect 218287 205581 218296 205615
rect 218244 205572 218296 205581
rect 384672 205615 384724 205624
rect 384672 205581 384681 205615
rect 384681 205581 384715 205615
rect 384715 205581 384724 205615
rect 384672 205572 384724 205581
rect 403532 205572 403584 205624
rect 403716 205572 403768 205624
rect 578056 205572 578108 205624
rect 580816 205572 580868 205624
rect 150808 205504 150860 205556
rect 190460 202852 190512 202904
rect 190644 202852 190696 202904
rect 208492 202852 208544 202904
rect 208584 202852 208636 202904
rect 211252 202852 211304 202904
rect 211344 202852 211396 202904
rect 214012 202895 214064 202904
rect 214012 202861 214021 202895
rect 214021 202861 214055 202895
rect 214055 202861 214064 202895
rect 214012 202852 214064 202861
rect 222476 202852 222528 202904
rect 222568 202852 222620 202904
rect 223856 202852 223908 202904
rect 223948 202852 224000 202904
rect 226524 202852 226576 202904
rect 226616 202852 226668 202904
rect 229284 202852 229336 202904
rect 229376 202852 229428 202904
rect 248144 202852 248196 202904
rect 248328 202852 248380 202904
rect 423220 202895 423272 202904
rect 423220 202861 423229 202895
rect 423229 202861 423263 202895
rect 423263 202861 423272 202895
rect 423220 202852 423272 202861
rect 424600 202852 424652 202904
rect 424692 202852 424744 202904
rect 423220 202759 423272 202768
rect 423220 202725 423229 202759
rect 423229 202725 423263 202759
rect 423263 202725 423272 202759
rect 423220 202716 423272 202725
rect 195980 201560 196032 201612
rect 196256 201560 196308 201612
rect 198372 201560 198424 201612
rect 150808 201424 150860 201476
rect 198372 201424 198424 201476
rect 205916 201424 205968 201476
rect 208400 201424 208452 201476
rect 208584 201424 208636 201476
rect 218244 201467 218296 201476
rect 218244 201433 218253 201467
rect 218253 201433 218287 201467
rect 218287 201433 218296 201467
rect 218244 201424 218296 201433
rect 222568 201424 222620 201476
rect 222660 201424 222712 201476
rect 226616 201424 226668 201476
rect 226800 201424 226852 201476
rect 229376 201424 229428 201476
rect 229468 201424 229520 201476
rect 238484 201424 238536 201476
rect 238668 201424 238720 201476
rect 248328 201424 248380 201476
rect 374276 201424 374328 201476
rect 374460 201424 374512 201476
rect 206008 201356 206060 201408
rect 226708 200064 226760 200116
rect 226800 200064 226852 200116
rect 223856 196052 223908 196104
rect 223764 195916 223816 195968
rect 2780 193876 2832 193928
rect 4988 193876 5040 193928
rect 234896 193264 234948 193316
rect 423312 193264 423364 193316
rect 168656 193196 168708 193248
rect 168840 193196 168892 193248
rect 169760 193196 169812 193248
rect 170036 193196 170088 193248
rect 178224 193196 178276 193248
rect 178408 193196 178460 193248
rect 190460 193196 190512 193248
rect 190736 193196 190788 193248
rect 191840 193196 191892 193248
rect 192024 193196 192076 193248
rect 207020 193196 207072 193248
rect 207204 193196 207256 193248
rect 214012 193196 214064 193248
rect 214104 193196 214156 193248
rect 234804 193196 234856 193248
rect 236276 193196 236328 193248
rect 236460 193196 236512 193248
rect 237564 193196 237616 193248
rect 237748 193196 237800 193248
rect 239036 193196 239088 193248
rect 239220 193196 239272 193248
rect 245936 193196 245988 193248
rect 246120 193196 246172 193248
rect 247040 193196 247092 193248
rect 247316 193196 247368 193248
rect 258080 193196 258132 193248
rect 258356 193196 258408 193248
rect 263600 193196 263652 193248
rect 263784 193196 263836 193248
rect 271880 193196 271932 193248
rect 272064 193196 272116 193248
rect 403808 193196 403860 193248
rect 403992 193196 404044 193248
rect 424508 193196 424560 193248
rect 424784 193196 424836 193248
rect 218336 193128 218388 193180
rect 248144 191879 248196 191888
rect 248144 191845 248153 191879
rect 248153 191845 248187 191879
rect 248187 191845 248196 191879
rect 248144 191836 248196 191845
rect 223764 191768 223816 191820
rect 224040 191768 224092 191820
rect 226432 190408 226484 190460
rect 226800 190408 226852 190460
rect 198280 189048 198332 189100
rect 198372 189048 198424 189100
rect 196348 188980 196400 189032
rect 162860 186328 162912 186380
rect 163044 186328 163096 186380
rect 173900 186328 173952 186380
rect 174084 186328 174136 186380
rect 252652 186328 252704 186380
rect 252836 186328 252888 186380
rect 284300 186328 284352 186380
rect 284484 186328 284536 186380
rect 307852 186328 307904 186380
rect 308036 186328 308088 186380
rect 346124 186328 346176 186380
rect 346308 186328 346360 186380
rect 357164 186328 357216 186380
rect 357348 186328 357400 186380
rect 423220 186328 423272 186380
rect 378876 183608 378928 183660
rect 379060 183608 379112 183660
rect 384580 183608 384632 183660
rect 384672 183608 384724 183660
rect 150808 183540 150860 183592
rect 151820 183540 151872 183592
rect 152004 183540 152056 183592
rect 218244 183540 218296 183592
rect 218428 183540 218480 183592
rect 238484 183540 238536 183592
rect 238668 183540 238720 183592
rect 248144 183540 248196 183592
rect 248328 183540 248380 183592
rect 423128 183583 423180 183592
rect 423128 183549 423137 183583
rect 423137 183549 423171 183583
rect 423171 183549 423180 183583
rect 423128 183540 423180 183549
rect 424600 183540 424652 183592
rect 424692 183540 424744 183592
rect 190736 183515 190788 183524
rect 190736 183481 190745 183515
rect 190745 183481 190779 183515
rect 190779 183481 190788 183515
rect 190736 183472 190788 183481
rect 219532 183515 219584 183524
rect 219532 183481 219541 183515
rect 219541 183481 219575 183515
rect 219575 183481 219584 183515
rect 219532 183472 219584 183481
rect 192024 183447 192076 183456
rect 192024 183413 192033 183447
rect 192033 183413 192067 183447
rect 192067 183413 192076 183447
rect 192024 183404 192076 183413
rect 218244 183447 218296 183456
rect 218244 183413 218253 183447
rect 218253 183413 218287 183447
rect 218287 183413 218296 183447
rect 218244 183404 218296 183413
rect 150808 182112 150860 182164
rect 152004 182112 152056 182164
rect 152188 182112 152240 182164
rect 238668 182112 238720 182164
rect 248144 182112 248196 182164
rect 248328 182112 248380 182164
rect 374276 182112 374328 182164
rect 374460 182112 374512 182164
rect 379060 182112 379112 182164
rect 379336 182112 379388 182164
rect 384580 182155 384632 182164
rect 384580 182121 384589 182155
rect 384589 182121 384623 182155
rect 384623 182121 384632 182155
rect 384580 182112 384632 182121
rect 423128 182112 423180 182164
rect 423220 182112 423272 182164
rect 424508 182155 424560 182164
rect 424508 182121 424517 182155
rect 424517 182121 424551 182155
rect 424551 182121 424560 182155
rect 424508 182112 424560 182121
rect 449164 182112 449216 182164
rect 580172 182112 580224 182164
rect 218336 180004 218388 180056
rect 219624 180004 219676 180056
rect 2780 179460 2832 179512
rect 4896 179460 4948 179512
rect 196256 179435 196308 179444
rect 196256 179401 196265 179435
rect 196265 179401 196299 179435
rect 196299 179401 196308 179435
rect 196256 179392 196308 179401
rect 194784 179367 194836 179376
rect 194784 179333 194793 179367
rect 194793 179333 194827 179367
rect 194827 179333 194836 179367
rect 194784 179324 194836 179333
rect 216588 178984 216640 179036
rect 216864 178984 216916 179036
rect 162952 176672 163004 176724
rect 156144 176604 156196 176656
rect 384580 176647 384632 176656
rect 384580 176613 384589 176647
rect 384589 176613 384623 176647
rect 384623 176613 384632 176647
rect 384580 176604 384632 176613
rect 163044 176536 163096 176588
rect 156144 176468 156196 176520
rect 154856 173952 154908 174004
rect 154948 173952 155000 174004
rect 168656 173884 168708 173936
rect 168840 173884 168892 173936
rect 169760 173884 169812 173936
rect 170036 173884 170088 173936
rect 174084 173884 174136 173936
rect 174268 173884 174320 173936
rect 178224 173884 178276 173936
rect 178408 173884 178460 173936
rect 190736 173927 190788 173936
rect 190736 173893 190745 173927
rect 190745 173893 190779 173927
rect 190779 173893 190788 173927
rect 190736 173884 190788 173893
rect 192024 173927 192076 173936
rect 192024 173893 192033 173927
rect 192033 173893 192067 173927
rect 192067 173893 192076 173927
rect 192024 173884 192076 173893
rect 205916 173884 205968 173936
rect 206100 173884 206152 173936
rect 207020 173884 207072 173936
rect 207204 173884 207256 173936
rect 208492 173884 208544 173936
rect 208584 173884 208636 173936
rect 211252 173884 211304 173936
rect 211344 173884 211396 173936
rect 222476 173884 222528 173936
rect 222660 173884 222712 173936
rect 226616 173952 226668 174004
rect 229284 173884 229336 173936
rect 229468 173884 229520 173936
rect 236276 173884 236328 173936
rect 236460 173884 236512 173936
rect 237564 173884 237616 173936
rect 237748 173884 237800 173936
rect 239036 173884 239088 173936
rect 239220 173884 239272 173936
rect 245936 173884 245988 173936
rect 246120 173884 246172 173936
rect 247040 173884 247092 173936
rect 247316 173884 247368 173936
rect 252560 173884 252612 173936
rect 252836 173884 252888 173936
rect 258080 173884 258132 173936
rect 258356 173884 258408 173936
rect 263600 173884 263652 173936
rect 263784 173884 263836 173936
rect 271880 173884 271932 173936
rect 272064 173884 272116 173936
rect 284484 173884 284536 173936
rect 284668 173884 284720 173936
rect 308036 173884 308088 173936
rect 308220 173884 308272 173936
rect 346032 173884 346084 173936
rect 346308 173884 346360 173936
rect 357072 173884 357124 173936
rect 357348 173884 357400 173936
rect 403808 173884 403860 173936
rect 403992 173884 404044 173936
rect 226524 173816 226576 173868
rect 424692 173816 424744 173868
rect 150716 173723 150768 173732
rect 150716 173689 150725 173723
rect 150725 173689 150759 173723
rect 150759 173689 150768 173723
rect 150716 173680 150768 173689
rect 238484 172567 238536 172576
rect 238484 172533 238493 172567
rect 238493 172533 238527 172567
rect 238527 172533 238536 172567
rect 238484 172524 238536 172533
rect 423312 172456 423364 172508
rect 424692 172456 424744 172508
rect 424968 172456 425020 172508
rect 219624 171028 219676 171080
rect 194784 169779 194836 169788
rect 194784 169745 194793 169779
rect 194793 169745 194827 169779
rect 194827 169745 194836 169779
rect 194784 169736 194836 169745
rect 194784 168351 194836 168360
rect 194784 168317 194793 168351
rect 194793 168317 194827 168351
rect 194827 168317 194836 168351
rect 194784 168308 194836 168317
rect 162860 167016 162912 167068
rect 163044 167016 163096 167068
rect 173900 167016 173952 167068
rect 174084 167016 174136 167068
rect 252652 167016 252704 167068
rect 252836 167016 252888 167068
rect 284300 167016 284352 167068
rect 284484 167016 284536 167068
rect 307852 167016 307904 167068
rect 308036 167016 308088 167068
rect 346124 167016 346176 167068
rect 346308 167016 346360 167068
rect 357164 167016 357216 167068
rect 357348 167016 357400 167068
rect 265072 166948 265124 167000
rect 270592 166948 270644 167000
rect 265072 166812 265124 166864
rect 270592 166812 270644 166864
rect 152004 164228 152056 164280
rect 152188 164228 152240 164280
rect 238484 164228 238536 164280
rect 238668 164228 238720 164280
rect 379152 164228 379204 164280
rect 379336 164228 379388 164280
rect 156144 164203 156196 164212
rect 156144 164169 156153 164203
rect 156153 164169 156187 164203
rect 156187 164169 156196 164203
rect 156144 164160 156196 164169
rect 169944 164160 169996 164212
rect 170036 164160 170088 164212
rect 173992 164203 174044 164212
rect 173992 164169 174001 164203
rect 174001 164169 174035 164203
rect 174035 164169 174044 164203
rect 173992 164160 174044 164169
rect 178224 164160 178276 164212
rect 178408 164160 178460 164212
rect 236276 164203 236328 164212
rect 236276 164169 236285 164203
rect 236285 164169 236319 164203
rect 236319 164169 236328 164203
rect 236276 164160 236328 164169
rect 237564 164203 237616 164212
rect 237564 164169 237573 164203
rect 237573 164169 237607 164203
rect 237607 164169 237616 164203
rect 237564 164160 237616 164169
rect 239036 164160 239088 164212
rect 239128 164160 239180 164212
rect 247040 164160 247092 164212
rect 247224 164160 247276 164212
rect 252744 164203 252796 164212
rect 252744 164169 252753 164203
rect 252753 164169 252787 164203
rect 252787 164169 252796 164203
rect 252744 164160 252796 164169
rect 258080 164160 258132 164212
rect 258264 164160 258316 164212
rect 284392 164203 284444 164212
rect 284392 164169 284401 164203
rect 284401 164169 284435 164203
rect 284435 164169 284444 164203
rect 284392 164160 284444 164169
rect 307944 164203 307996 164212
rect 307944 164169 307953 164203
rect 307953 164169 307987 164203
rect 307987 164169 307996 164203
rect 307944 164160 307996 164169
rect 346216 164203 346268 164212
rect 346216 164169 346225 164203
rect 346225 164169 346259 164203
rect 346259 164169 346268 164203
rect 346216 164160 346268 164169
rect 357256 164203 357308 164212
rect 357256 164169 357265 164203
rect 357265 164169 357299 164203
rect 357299 164169 357308 164203
rect 357256 164160 357308 164169
rect 403532 164160 403584 164212
rect 403716 164160 403768 164212
rect 196256 162868 196308 162920
rect 423220 162911 423272 162920
rect 423220 162877 423229 162911
rect 423229 162877 423263 162911
rect 423263 162877 423272 162911
rect 423220 162868 423272 162877
rect 190460 162800 190512 162852
rect 190644 162800 190696 162852
rect 198280 162800 198332 162852
rect 198372 162800 198424 162852
rect 206008 162843 206060 162852
rect 206008 162809 206017 162843
rect 206017 162809 206051 162843
rect 206051 162809 206060 162843
rect 206008 162800 206060 162809
rect 238392 162800 238444 162852
rect 238668 162800 238720 162852
rect 248328 162843 248380 162852
rect 248328 162809 248337 162843
rect 248337 162809 248371 162843
rect 248371 162809 248380 162843
rect 248328 162800 248380 162809
rect 265072 162800 265124 162852
rect 265256 162800 265308 162852
rect 270592 162800 270644 162852
rect 270776 162800 270828 162852
rect 374276 162843 374328 162852
rect 374276 162809 374285 162843
rect 374285 162809 374319 162843
rect 374319 162809 374328 162843
rect 374276 162800 374328 162809
rect 379060 162843 379112 162852
rect 379060 162809 379069 162843
rect 379069 162809 379103 162843
rect 379103 162809 379112 162843
rect 379060 162800 379112 162809
rect 384580 162843 384632 162852
rect 384580 162809 384589 162843
rect 384589 162809 384623 162843
rect 384623 162809 384632 162843
rect 384580 162800 384632 162809
rect 424692 162843 424744 162852
rect 424692 162809 424701 162843
rect 424701 162809 424735 162843
rect 424735 162809 424744 162843
rect 424692 162800 424744 162809
rect 196256 162732 196308 162784
rect 219532 162435 219584 162444
rect 219532 162401 219541 162435
rect 219541 162401 219575 162435
rect 219575 162401 219584 162435
rect 219532 162392 219584 162401
rect 216772 161415 216824 161424
rect 216772 161381 216781 161415
rect 216781 161381 216815 161415
rect 216815 161381 216824 161415
rect 216772 161372 216824 161381
rect 217968 161372 218020 161424
rect 218244 161372 218296 161424
rect 219532 160055 219584 160064
rect 219532 160021 219541 160055
rect 219541 160021 219575 160055
rect 219575 160021 219584 160055
rect 219532 160012 219584 160021
rect 194876 158720 194928 158772
rect 198372 158652 198424 158704
rect 577964 158652 578016 158704
rect 580080 158652 580132 158704
rect 207112 157428 207164 157480
rect 208492 157428 208544 157480
rect 162952 157360 163004 157412
rect 211252 157360 211304 157412
rect 423220 157360 423272 157412
rect 173992 157335 174044 157344
rect 173992 157301 174001 157335
rect 174001 157301 174035 157335
rect 174035 157301 174044 157335
rect 173992 157292 174044 157301
rect 206008 157335 206060 157344
rect 206008 157301 206017 157335
rect 206017 157301 206051 157335
rect 206051 157301 206060 157335
rect 206008 157292 206060 157301
rect 207112 157292 207164 157344
rect 208492 157292 208544 157344
rect 252744 157335 252796 157344
rect 252744 157301 252753 157335
rect 252753 157301 252787 157335
rect 252787 157301 252796 157335
rect 252744 157292 252796 157301
rect 284392 157335 284444 157344
rect 284392 157301 284401 157335
rect 284401 157301 284435 157335
rect 284435 157301 284444 157335
rect 284392 157292 284444 157301
rect 307944 157335 307996 157344
rect 307944 157301 307953 157335
rect 307953 157301 307987 157335
rect 307987 157301 307996 157335
rect 307944 157292 307996 157301
rect 346216 157335 346268 157344
rect 346216 157301 346225 157335
rect 346225 157301 346259 157335
rect 346259 157301 346268 157335
rect 346216 157292 346268 157301
rect 357256 157335 357308 157344
rect 357256 157301 357265 157335
rect 357265 157301 357299 157335
rect 357299 157301 357308 157335
rect 357256 157292 357308 157301
rect 379060 157335 379112 157344
rect 379060 157301 379069 157335
rect 379069 157301 379103 157335
rect 379103 157301 379112 157335
rect 379060 157292 379112 157301
rect 163044 157224 163096 157276
rect 211252 157224 211304 157276
rect 236276 157267 236328 157276
rect 236276 157233 236285 157267
rect 236285 157233 236319 157267
rect 236319 157233 236328 157267
rect 236276 157224 236328 157233
rect 237564 157267 237616 157276
rect 237564 157233 237573 157267
rect 237573 157233 237607 157267
rect 237607 157233 237616 157267
rect 237564 157224 237616 157233
rect 424692 157335 424744 157344
rect 424692 157301 424701 157335
rect 424701 157301 424735 157335
rect 424735 157301 424744 157335
rect 424692 157292 424744 157301
rect 423312 157224 423364 157276
rect 156144 154615 156196 154624
rect 156144 154581 156153 154615
rect 156153 154581 156187 154615
rect 156187 154581 156196 154615
rect 156144 154572 156196 154581
rect 229192 154572 229244 154624
rect 229284 154572 229336 154624
rect 222476 154504 222528 154556
rect 222660 154504 222712 154556
rect 223764 154504 223816 154556
rect 223948 154504 224000 154556
rect 226524 154504 226576 154556
rect 226616 154504 226668 154556
rect 239036 154504 239088 154556
rect 263784 154547 263836 154556
rect 263784 154513 263793 154547
rect 263793 154513 263827 154547
rect 263827 154513 263836 154547
rect 263784 154504 263836 154513
rect 271880 154504 271932 154556
rect 272064 154504 272116 154556
rect 239128 154436 239180 154488
rect 248328 153255 248380 153264
rect 248328 153221 248337 153255
rect 248337 153221 248371 153255
rect 248371 153221 248380 153255
rect 248328 153212 248380 153221
rect 374276 153255 374328 153264
rect 374276 153221 374285 153255
rect 374285 153221 374319 153255
rect 374319 153221 374328 153255
rect 374276 153212 374328 153221
rect 384580 153255 384632 153264
rect 384580 153221 384589 153255
rect 384589 153221 384623 153255
rect 384623 153221 384632 153255
rect 384580 153212 384632 153221
rect 423312 153144 423364 153196
rect 424692 153144 424744 153196
rect 424784 153144 424836 153196
rect 216864 151784 216916 151836
rect 3332 151716 3384 151768
rect 19984 151716 20036 151768
rect 219624 150424 219676 150476
rect 194784 150356 194836 150408
rect 198280 149107 198332 149116
rect 198280 149073 198289 149107
rect 198289 149073 198323 149107
rect 198323 149073 198332 149107
rect 198280 149064 198332 149073
rect 263784 148359 263836 148368
rect 263784 148325 263793 148359
rect 263793 148325 263827 148359
rect 263827 148325 263836 148359
rect 263784 148316 263836 148325
rect 162860 147636 162912 147688
rect 163044 147636 163096 147688
rect 173900 147636 173952 147688
rect 174084 147636 174136 147688
rect 252652 147636 252704 147688
rect 252836 147636 252888 147688
rect 284300 147636 284352 147688
rect 284484 147636 284536 147688
rect 307852 147636 307904 147688
rect 308036 147636 308088 147688
rect 346124 147636 346176 147688
rect 346308 147636 346360 147688
rect 357164 147636 357216 147688
rect 357348 147636 357400 147688
rect 238576 144916 238628 144968
rect 238668 144916 238720 144968
rect 379152 144916 379204 144968
rect 173992 144891 174044 144900
rect 173992 144857 174001 144891
rect 174001 144857 174035 144891
rect 174035 144857 174044 144891
rect 173992 144848 174044 144857
rect 178224 144848 178276 144900
rect 178408 144848 178460 144900
rect 190644 144848 190696 144900
rect 191840 144848 191892 144900
rect 191932 144848 191984 144900
rect 205916 144848 205968 144900
rect 206008 144848 206060 144900
rect 207112 144848 207164 144900
rect 207204 144848 207256 144900
rect 208492 144848 208544 144900
rect 208676 144848 208728 144900
rect 211252 144848 211304 144900
rect 211436 144848 211488 144900
rect 234896 144848 234948 144900
rect 234988 144848 235040 144900
rect 236276 144848 236328 144900
rect 236368 144848 236420 144900
rect 237564 144848 237616 144900
rect 237656 144848 237708 144900
rect 239036 144848 239088 144900
rect 239128 144848 239180 144900
rect 252744 144891 252796 144900
rect 252744 144857 252753 144891
rect 252753 144857 252787 144891
rect 252787 144857 252796 144891
rect 252744 144848 252796 144857
rect 284392 144891 284444 144900
rect 284392 144857 284401 144891
rect 284401 144857 284435 144891
rect 284435 144857 284444 144891
rect 284392 144848 284444 144857
rect 303896 144848 303948 144900
rect 303988 144848 304040 144900
rect 307944 144891 307996 144900
rect 307944 144857 307953 144891
rect 307953 144857 307987 144891
rect 307987 144857 307996 144891
rect 307944 144848 307996 144857
rect 346216 144891 346268 144900
rect 346216 144857 346225 144891
rect 346225 144857 346259 144891
rect 346259 144857 346268 144891
rect 346216 144848 346268 144857
rect 357256 144891 357308 144900
rect 357256 144857 357265 144891
rect 357265 144857 357299 144891
rect 357299 144857 357308 144891
rect 357256 144848 357308 144857
rect 190736 144780 190788 144832
rect 379152 144780 379204 144832
rect 384580 144780 384632 144832
rect 384856 144780 384908 144832
rect 423220 143599 423272 143608
rect 423220 143565 423229 143599
rect 423229 143565 423263 143599
rect 423263 143565 423272 143599
rect 423220 143556 423272 143565
rect 162952 143531 163004 143540
rect 162952 143497 162961 143531
rect 162961 143497 162995 143531
rect 162995 143497 163004 143531
rect 162952 143488 163004 143497
rect 189264 143531 189316 143540
rect 189264 143497 189273 143531
rect 189273 143497 189307 143531
rect 189307 143497 189316 143531
rect 189264 143488 189316 143497
rect 190368 143488 190420 143540
rect 190736 143488 190788 143540
rect 205916 143488 205968 143540
rect 206100 143488 206152 143540
rect 238668 143531 238720 143540
rect 238668 143497 238677 143531
rect 238677 143497 238711 143531
rect 238711 143497 238720 143531
rect 238668 143488 238720 143497
rect 245752 143488 245804 143540
rect 248328 143531 248380 143540
rect 248328 143497 248337 143531
rect 248337 143497 248371 143531
rect 248371 143497 248380 143531
rect 248328 143488 248380 143497
rect 374276 143531 374328 143540
rect 374276 143497 374285 143531
rect 374285 143497 374319 143531
rect 374319 143497 374328 143531
rect 374276 143488 374328 143497
rect 424692 143531 424744 143540
rect 424692 143497 424701 143531
rect 424701 143497 424735 143531
rect 424735 143497 424744 143531
rect 424692 143488 424744 143497
rect 245936 143420 245988 143472
rect 196256 142196 196308 142248
rect 217968 142128 218020 142180
rect 218428 142128 218480 142180
rect 152004 142060 152056 142112
rect 152188 142060 152240 142112
rect 196164 142060 196216 142112
rect 263784 142103 263836 142112
rect 263784 142069 263793 142103
rect 263793 142069 263827 142103
rect 263827 142069 263836 142103
rect 263784 142060 263836 142069
rect 379152 142103 379204 142112
rect 379152 142069 379161 142103
rect 379161 142069 379195 142103
rect 379195 142069 379204 142103
rect 379152 142060 379204 142069
rect 194692 140811 194744 140820
rect 194692 140777 194701 140811
rect 194701 140777 194735 140811
rect 194735 140777 194744 140811
rect 194692 140768 194744 140777
rect 150716 140700 150768 140752
rect 152188 140743 152240 140752
rect 152188 140709 152197 140743
rect 152197 140709 152231 140743
rect 152231 140709 152240 140743
rect 152188 140700 152240 140709
rect 198280 138048 198332 138100
rect 247224 137980 247276 138032
rect 162952 137955 163004 137964
rect 162952 137921 162961 137955
rect 162961 137921 162995 137955
rect 162995 137921 163004 137955
rect 162952 137912 163004 137921
rect 173992 137955 174044 137964
rect 173992 137921 174001 137955
rect 174001 137921 174035 137955
rect 174035 137921 174044 137955
rect 173992 137912 174044 137921
rect 198280 137912 198332 137964
rect 403624 138048 403676 138100
rect 423220 137980 423272 138032
rect 247316 137912 247368 137964
rect 252744 137955 252796 137964
rect 252744 137921 252753 137955
rect 252753 137921 252787 137955
rect 252787 137921 252796 137955
rect 252744 137912 252796 137921
rect 284392 137955 284444 137964
rect 284392 137921 284401 137955
rect 284401 137921 284435 137955
rect 284435 137921 284444 137955
rect 284392 137912 284444 137921
rect 307944 137955 307996 137964
rect 307944 137921 307953 137955
rect 307953 137921 307987 137955
rect 307987 137921 307996 137955
rect 307944 137912 307996 137921
rect 346216 137955 346268 137964
rect 346216 137921 346225 137955
rect 346225 137921 346259 137955
rect 346259 137921 346268 137955
rect 346216 137912 346268 137921
rect 357256 137955 357308 137964
rect 357256 137921 357265 137955
rect 357265 137921 357299 137955
rect 357299 137921 357308 137955
rect 357256 137912 357308 137921
rect 403532 137912 403584 137964
rect 423312 137912 423364 137964
rect 424692 137955 424744 137964
rect 424692 137921 424701 137955
rect 424701 137921 424735 137955
rect 424735 137921 424744 137955
rect 424692 137912 424744 137921
rect 216864 135192 216916 135244
rect 234804 135192 234856 135244
rect 234988 135192 235040 135244
rect 271880 135192 271932 135244
rect 272064 135192 272116 135244
rect 403256 135192 403308 135244
rect 403532 135192 403584 135244
rect 577872 135192 577924 135244
rect 580632 135192 580684 135244
rect 168748 133968 168800 134020
rect 168840 133968 168892 134020
rect 189264 133943 189316 133952
rect 189264 133909 189273 133943
rect 189273 133909 189307 133943
rect 189307 133909 189316 133943
rect 189264 133900 189316 133909
rect 248328 133943 248380 133952
rect 248328 133909 248337 133943
rect 248337 133909 248371 133943
rect 248371 133909 248380 133943
rect 248328 133900 248380 133909
rect 374276 133943 374328 133952
rect 374276 133909 374285 133943
rect 374285 133909 374319 133943
rect 374319 133909 374328 133943
rect 374276 133900 374328 133909
rect 153384 133875 153436 133884
rect 153384 133841 153393 133875
rect 153393 133841 153427 133875
rect 153427 133841 153436 133875
rect 153384 133832 153436 133841
rect 156144 133875 156196 133884
rect 156144 133841 156153 133875
rect 156153 133841 156187 133875
rect 156187 133841 156196 133875
rect 156144 133832 156196 133841
rect 168840 133875 168892 133884
rect 168840 133841 168849 133875
rect 168849 133841 168883 133875
rect 168883 133841 168892 133875
rect 168840 133832 168892 133841
rect 190460 133832 190512 133884
rect 190644 133832 190696 133884
rect 234988 133832 235040 133884
rect 245936 133832 245988 133884
rect 384672 133875 384724 133884
rect 384672 133841 384681 133875
rect 384681 133841 384715 133875
rect 384715 133841 384724 133875
rect 384672 133832 384724 133841
rect 424784 133832 424836 133884
rect 263784 132515 263836 132524
rect 263784 132481 263793 132515
rect 263793 132481 263827 132515
rect 263827 132481 263836 132515
rect 263784 132472 263836 132481
rect 379244 132472 379296 132524
rect 192024 132447 192076 132456
rect 192024 132413 192033 132447
rect 192033 132413 192067 132447
rect 192067 132413 192076 132447
rect 192024 132404 192076 132413
rect 379244 132336 379296 132388
rect 150808 131155 150860 131164
rect 150808 131121 150817 131155
rect 150817 131121 150851 131155
rect 150851 131121 150860 131155
rect 152188 131155 152240 131164
rect 150808 131112 150860 131121
rect 152188 131121 152197 131155
rect 152197 131121 152231 131155
rect 152231 131121 152240 131155
rect 152188 131112 152240 131121
rect 216772 129727 216824 129736
rect 216772 129693 216781 129727
rect 216781 129693 216815 129727
rect 216815 129693 216824 129727
rect 216772 129684 216824 129693
rect 423312 129004 423364 129056
rect 423496 129004 423548 129056
rect 162860 128324 162912 128376
rect 163044 128324 163096 128376
rect 173900 128324 173952 128376
rect 174084 128324 174136 128376
rect 218336 128392 218388 128444
rect 252652 128324 252704 128376
rect 252836 128324 252888 128376
rect 284300 128324 284352 128376
rect 284484 128324 284536 128376
rect 307852 128324 307904 128376
rect 308036 128324 308088 128376
rect 346124 128324 346176 128376
rect 346308 128324 346360 128376
rect 357164 128324 357216 128376
rect 357348 128324 357400 128376
rect 218244 128256 218296 128308
rect 384672 127823 384724 127832
rect 384672 127789 384681 127823
rect 384681 127789 384715 127823
rect 384715 127789 384724 127823
rect 384672 127780 384724 127789
rect 238668 125647 238720 125656
rect 238668 125613 238677 125647
rect 238677 125613 238711 125647
rect 238711 125613 238720 125647
rect 238668 125604 238720 125613
rect 173992 125579 174044 125588
rect 173992 125545 174001 125579
rect 174001 125545 174035 125579
rect 174035 125545 174044 125579
rect 173992 125536 174044 125545
rect 178224 125579 178276 125588
rect 178224 125545 178233 125579
rect 178233 125545 178267 125579
rect 178267 125545 178276 125579
rect 178224 125536 178276 125545
rect 205824 125536 205876 125588
rect 206008 125536 206060 125588
rect 208492 125536 208544 125588
rect 208676 125536 208728 125588
rect 211252 125536 211304 125588
rect 216772 125536 216824 125588
rect 216956 125536 217008 125588
rect 218244 125536 218296 125588
rect 218428 125536 218480 125588
rect 219532 125536 219584 125588
rect 219716 125536 219768 125588
rect 238944 125536 238996 125588
rect 239128 125536 239180 125588
rect 252744 125579 252796 125588
rect 252744 125545 252753 125579
rect 252753 125545 252787 125579
rect 252787 125545 252796 125579
rect 252744 125536 252796 125545
rect 284392 125579 284444 125588
rect 284392 125545 284401 125579
rect 284401 125545 284435 125579
rect 284435 125545 284444 125579
rect 284392 125536 284444 125545
rect 303896 125536 303948 125588
rect 303988 125536 304040 125588
rect 307944 125579 307996 125588
rect 307944 125545 307953 125579
rect 307953 125545 307987 125579
rect 307987 125545 307996 125579
rect 307944 125536 307996 125545
rect 346216 125579 346268 125588
rect 346216 125545 346225 125579
rect 346225 125545 346259 125579
rect 346259 125545 346268 125579
rect 346216 125536 346268 125545
rect 357256 125579 357308 125588
rect 357256 125545 357265 125579
rect 357265 125545 357299 125579
rect 357299 125545 357308 125579
rect 357256 125536 357308 125545
rect 211344 125468 211396 125520
rect 234804 124287 234856 124296
rect 234804 124253 234813 124287
rect 234813 124253 234847 124287
rect 234847 124253 234856 124287
rect 234804 124244 234856 124253
rect 424692 124287 424744 124296
rect 424692 124253 424701 124287
rect 424701 124253 424735 124287
rect 424735 124253 424744 124287
rect 424692 124244 424744 124253
rect 153384 124219 153436 124228
rect 153384 124185 153393 124219
rect 153393 124185 153427 124219
rect 153427 124185 153436 124219
rect 153384 124176 153436 124185
rect 156144 124219 156196 124228
rect 156144 124185 156153 124219
rect 156153 124185 156187 124219
rect 156187 124185 156196 124219
rect 156144 124176 156196 124185
rect 168840 124219 168892 124228
rect 168840 124185 168849 124219
rect 168849 124185 168883 124219
rect 168883 124185 168892 124219
rect 168840 124176 168892 124185
rect 245752 124219 245804 124228
rect 245752 124185 245761 124219
rect 245761 124185 245795 124219
rect 245795 124185 245804 124219
rect 245752 124176 245804 124185
rect 162952 124151 163004 124160
rect 162952 124117 162961 124151
rect 162961 124117 162995 124151
rect 162995 124117 163004 124151
rect 162952 124108 163004 124117
rect 189264 124151 189316 124160
rect 189264 124117 189273 124151
rect 189273 124117 189307 124151
rect 189307 124117 189316 124151
rect 189264 124108 189316 124117
rect 190644 124108 190696 124160
rect 192024 124151 192076 124160
rect 192024 124117 192033 124151
rect 192033 124117 192067 124151
rect 192067 124117 192076 124151
rect 192024 124108 192076 124117
rect 234804 124151 234856 124160
rect 234804 124117 234813 124151
rect 234813 124117 234847 124151
rect 234847 124117 234856 124151
rect 234804 124108 234856 124117
rect 238668 124108 238720 124160
rect 248328 124151 248380 124160
rect 248328 124117 248337 124151
rect 248337 124117 248371 124151
rect 248371 124117 248380 124151
rect 248328 124108 248380 124117
rect 374276 124151 374328 124160
rect 374276 124117 374285 124151
rect 374285 124117 374319 124151
rect 374319 124117 374328 124151
rect 374276 124108 374328 124117
rect 384396 124108 384448 124160
rect 384488 124108 384540 124160
rect 424692 124151 424744 124160
rect 424692 124117 424701 124151
rect 424701 124117 424735 124151
rect 424735 124117 424744 124151
rect 424692 124108 424744 124117
rect 190920 124040 190972 124092
rect 384488 123972 384540 124024
rect 384396 123904 384448 123956
rect 152004 122816 152056 122868
rect 152096 122816 152148 122868
rect 196164 122816 196216 122868
rect 196256 122816 196308 122868
rect 379152 122859 379204 122868
rect 379152 122825 379161 122859
rect 379161 122825 379195 122859
rect 379195 122825 379204 122859
rect 379152 122816 379204 122825
rect 263784 122791 263836 122800
rect 263784 122757 263793 122791
rect 263793 122757 263827 122791
rect 263827 122757 263836 122791
rect 263784 122748 263836 122757
rect 264980 122791 265032 122800
rect 264980 122757 264989 122791
rect 264989 122757 265023 122791
rect 265023 122757 265032 122791
rect 264980 122748 265032 122757
rect 423220 122791 423272 122800
rect 423220 122757 423229 122791
rect 423229 122757 423263 122791
rect 423263 122757 423272 122791
rect 423220 122748 423272 122757
rect 152004 121431 152056 121440
rect 152004 121397 152013 121431
rect 152013 121397 152047 121431
rect 152047 121397 152056 121431
rect 152004 121388 152056 121397
rect 208584 120504 208636 120556
rect 208676 120504 208728 120556
rect 156144 118736 156196 118788
rect 222568 118736 222620 118788
rect 223856 118736 223908 118788
rect 247224 118668 247276 118720
rect 403440 118668 403492 118720
rect 156144 118600 156196 118652
rect 173992 118643 174044 118652
rect 173992 118609 174001 118643
rect 174001 118609 174035 118643
rect 174035 118609 174044 118643
rect 173992 118600 174044 118609
rect 222568 118600 222620 118652
rect 223856 118600 223908 118652
rect 247316 118600 247368 118652
rect 252744 118643 252796 118652
rect 252744 118609 252753 118643
rect 252753 118609 252787 118643
rect 252787 118609 252796 118643
rect 252744 118600 252796 118609
rect 284392 118643 284444 118652
rect 284392 118609 284401 118643
rect 284401 118609 284435 118643
rect 284435 118609 284444 118643
rect 284392 118600 284444 118609
rect 307944 118643 307996 118652
rect 307944 118609 307953 118643
rect 307953 118609 307987 118643
rect 307987 118609 307996 118643
rect 307944 118600 307996 118609
rect 346216 118643 346268 118652
rect 346216 118609 346225 118643
rect 346225 118609 346259 118643
rect 346259 118609 346268 118643
rect 346216 118600 346268 118609
rect 357256 118643 357308 118652
rect 357256 118609 357265 118643
rect 357265 118609 357299 118643
rect 357299 118609 357308 118643
rect 357256 118600 357308 118609
rect 403532 118600 403584 118652
rect 150716 116331 150768 116340
rect 150716 116297 150725 116331
rect 150725 116297 150759 116331
rect 150759 116297 150768 116331
rect 150716 116288 150768 116297
rect 178224 115991 178276 116000
rect 178224 115957 178233 115991
rect 178233 115957 178267 115991
rect 178267 115957 178276 115991
rect 178224 115948 178276 115957
rect 236276 115880 236328 115932
rect 237564 115880 237616 115932
rect 403256 115880 403308 115932
rect 403532 115880 403584 115932
rect 168840 115812 168892 115864
rect 236368 115812 236420 115864
rect 237656 115812 237708 115864
rect 168748 115744 168800 115796
rect 153476 114588 153528 114640
rect 153292 114520 153344 114572
rect 216956 114588 217008 114640
rect 163044 114520 163096 114572
rect 189264 114563 189316 114572
rect 189264 114529 189273 114563
rect 189273 114529 189307 114563
rect 189307 114529 189316 114563
rect 189264 114520 189316 114529
rect 216864 114520 216916 114572
rect 234804 114563 234856 114572
rect 234804 114529 234813 114563
rect 234813 114529 234847 114563
rect 234847 114529 234856 114563
rect 234804 114520 234856 114529
rect 238576 114563 238628 114572
rect 238576 114529 238585 114563
rect 238585 114529 238619 114563
rect 238619 114529 238628 114563
rect 238576 114520 238628 114529
rect 248328 114563 248380 114572
rect 248328 114529 248337 114563
rect 248337 114529 248371 114563
rect 248371 114529 248380 114563
rect 248328 114520 248380 114529
rect 374276 114563 374328 114572
rect 374276 114529 374285 114563
rect 374285 114529 374319 114563
rect 374319 114529 374328 114563
rect 374276 114520 374328 114529
rect 384580 114520 384632 114572
rect 384672 114520 384724 114572
rect 424784 114520 424836 114572
rect 168840 114495 168892 114504
rect 168840 114461 168849 114495
rect 168849 114461 168883 114495
rect 168883 114461 168892 114495
rect 168840 114452 168892 114461
rect 207020 114495 207072 114504
rect 207020 114461 207029 114495
rect 207029 114461 207063 114495
rect 207063 114461 207072 114495
rect 207020 114452 207072 114461
rect 271972 114452 272024 114504
rect 272064 114452 272116 114504
rect 153292 114427 153344 114436
rect 153292 114393 153301 114427
rect 153301 114393 153335 114427
rect 153335 114393 153344 114427
rect 153292 114384 153344 114393
rect 384580 114427 384632 114436
rect 384580 114393 384589 114427
rect 384589 114393 384623 114427
rect 384623 114393 384632 114427
rect 384580 114384 384632 114393
rect 263784 114291 263836 114300
rect 263784 114257 263793 114291
rect 263793 114257 263827 114291
rect 263827 114257 263836 114291
rect 263784 114248 263836 114257
rect 192024 113228 192076 113280
rect 194692 113160 194744 113212
rect 194784 113160 194836 113212
rect 196164 113160 196216 113212
rect 196256 113160 196308 113212
rect 265072 113160 265124 113212
rect 423312 113160 423364 113212
rect 152004 111843 152056 111852
rect 152004 111809 152013 111843
rect 152013 111809 152047 111843
rect 152047 111809 152056 111843
rect 152004 111800 152056 111809
rect 191932 111843 191984 111852
rect 191932 111809 191941 111843
rect 191941 111809 191975 111843
rect 191975 111809 191984 111843
rect 191932 111800 191984 111809
rect 577780 111732 577832 111784
rect 580632 111732 580684 111784
rect 245936 109692 245988 109744
rect 423312 109692 423364 109744
rect 218336 109080 218388 109132
rect 219624 109080 219676 109132
rect 162860 109012 162912 109064
rect 163044 109012 163096 109064
rect 173900 109012 173952 109064
rect 174084 109012 174136 109064
rect 252652 109012 252704 109064
rect 252836 109012 252888 109064
rect 284300 109012 284352 109064
rect 284484 109012 284536 109064
rect 307852 109012 307904 109064
rect 308036 109012 308088 109064
rect 346124 109012 346176 109064
rect 346308 109012 346360 109064
rect 357164 109012 357216 109064
rect 357348 109012 357400 109064
rect 218336 108944 218388 108996
rect 219624 108944 219676 108996
rect 424784 107040 424836 107092
rect 208584 106292 208636 106344
rect 211344 106292 211396 106344
rect 238576 106292 238628 106344
rect 238668 106292 238720 106344
rect 168840 106267 168892 106276
rect 168840 106233 168849 106267
rect 168849 106233 168883 106267
rect 168883 106233 168892 106267
rect 168840 106224 168892 106233
rect 173992 106267 174044 106276
rect 173992 106233 174001 106267
rect 174001 106233 174035 106267
rect 174035 106233 174044 106267
rect 173992 106224 174044 106233
rect 178224 106267 178276 106276
rect 178224 106233 178233 106267
rect 178233 106233 178267 106267
rect 178267 106233 178276 106267
rect 178224 106224 178276 106233
rect 190644 106267 190696 106276
rect 190644 106233 190653 106267
rect 190653 106233 190687 106267
rect 190687 106233 190696 106267
rect 190644 106224 190696 106233
rect 154764 106199 154816 106208
rect 154764 106165 154773 106199
rect 154773 106165 154807 106199
rect 154807 106165 154816 106199
rect 154764 106156 154816 106165
rect 222476 106224 222528 106276
rect 222568 106224 222620 106276
rect 223764 106224 223816 106276
rect 223856 106224 223908 106276
rect 252744 106267 252796 106276
rect 252744 106233 252753 106267
rect 252753 106233 252787 106267
rect 252787 106233 252796 106267
rect 252744 106224 252796 106233
rect 284392 106267 284444 106276
rect 284392 106233 284401 106267
rect 284401 106233 284435 106267
rect 284435 106233 284444 106267
rect 284392 106224 284444 106233
rect 307944 106267 307996 106276
rect 307944 106233 307953 106267
rect 307953 106233 307987 106267
rect 307987 106233 307996 106267
rect 307944 106224 307996 106233
rect 346216 106267 346268 106276
rect 346216 106233 346225 106267
rect 346225 106233 346259 106267
rect 346259 106233 346268 106267
rect 346216 106224 346268 106233
rect 357256 106267 357308 106276
rect 357256 106233 357265 106267
rect 357265 106233 357299 106267
rect 357299 106233 357308 106267
rect 357256 106224 357308 106233
rect 211344 106088 211396 106140
rect 153384 104864 153436 104916
rect 189172 104864 189224 104916
rect 189264 104864 189316 104916
rect 205824 104864 205876 104916
rect 206008 104864 206060 104916
rect 207112 104864 207164 104916
rect 208400 104907 208452 104916
rect 208400 104873 208409 104907
rect 208409 104873 208443 104907
rect 208443 104873 208452 104907
rect 208400 104864 208452 104873
rect 245752 104907 245804 104916
rect 245752 104873 245761 104907
rect 245761 104873 245795 104907
rect 245795 104873 245804 104907
rect 245752 104864 245804 104873
rect 384856 104864 384908 104916
rect 423036 104907 423088 104916
rect 423036 104873 423045 104907
rect 423045 104873 423079 104907
rect 423079 104873 423088 104907
rect 423036 104864 423088 104873
rect 168840 104839 168892 104848
rect 168840 104805 168849 104839
rect 168849 104805 168883 104839
rect 168883 104805 168892 104839
rect 168840 104796 168892 104805
rect 222476 104796 222528 104848
rect 223764 104839 223816 104848
rect 223764 104805 223773 104839
rect 223773 104805 223807 104839
rect 223807 104805 223816 104839
rect 223764 104796 223816 104805
rect 238668 104839 238720 104848
rect 238668 104805 238677 104839
rect 238677 104805 238711 104839
rect 238711 104805 238720 104839
rect 238668 104796 238720 104805
rect 248328 104839 248380 104848
rect 248328 104805 248337 104839
rect 248337 104805 248371 104839
rect 248371 104805 248380 104839
rect 248328 104796 248380 104805
rect 263784 104839 263836 104848
rect 263784 104805 263793 104839
rect 263793 104805 263827 104839
rect 263827 104805 263836 104839
rect 263784 104796 263836 104805
rect 374276 104839 374328 104848
rect 374276 104805 374285 104839
rect 374285 104805 374319 104839
rect 374319 104805 374328 104839
rect 374276 104796 374328 104805
rect 222568 104728 222620 104780
rect 150808 103504 150860 103556
rect 206008 103479 206060 103488
rect 206008 103445 206017 103479
rect 206017 103445 206051 103479
rect 206051 103445 206060 103479
rect 206008 103436 206060 103445
rect 208400 103479 208452 103488
rect 208400 103445 208409 103479
rect 208409 103445 208443 103479
rect 208443 103445 208452 103479
rect 208400 103436 208452 103445
rect 270500 103479 270552 103488
rect 270500 103445 270509 103479
rect 270509 103445 270543 103479
rect 270543 103445 270552 103479
rect 270500 103436 270552 103445
rect 272064 103479 272116 103488
rect 272064 103445 272073 103479
rect 272073 103445 272107 103479
rect 272107 103445 272116 103479
rect 272064 103436 272116 103445
rect 191748 102144 191800 102196
rect 192208 102144 192260 102196
rect 152004 102119 152056 102128
rect 152004 102085 152013 102119
rect 152013 102085 152047 102119
rect 152047 102085 152056 102119
rect 152004 102076 152056 102085
rect 190644 101371 190696 101380
rect 190644 101337 190653 101371
rect 190653 101337 190687 101371
rect 190687 101337 190696 101371
rect 190644 101328 190696 101337
rect 379152 100079 379204 100088
rect 379152 100045 379161 100079
rect 379161 100045 379195 100079
rect 379195 100045 379204 100079
rect 379152 100036 379204 100045
rect 153384 99424 153436 99476
rect 156144 99424 156196 99476
rect 214104 99424 214156 99476
rect 162952 99356 163004 99408
rect 153384 99288 153436 99340
rect 156144 99288 156196 99340
rect 247224 99356 247276 99408
rect 403440 99356 403492 99408
rect 163044 99288 163096 99340
rect 173992 99331 174044 99340
rect 173992 99297 174001 99331
rect 174001 99297 174035 99331
rect 174035 99297 174044 99331
rect 173992 99288 174044 99297
rect 214104 99288 214156 99340
rect 247316 99288 247368 99340
rect 252744 99331 252796 99340
rect 252744 99297 252753 99331
rect 252753 99297 252787 99331
rect 252787 99297 252796 99331
rect 252744 99288 252796 99297
rect 284392 99331 284444 99340
rect 284392 99297 284401 99331
rect 284401 99297 284435 99331
rect 284435 99297 284444 99331
rect 284392 99288 284444 99297
rect 307944 99331 307996 99340
rect 307944 99297 307953 99331
rect 307953 99297 307987 99331
rect 307987 99297 307996 99331
rect 307944 99288 307996 99297
rect 346216 99331 346268 99340
rect 346216 99297 346225 99331
rect 346225 99297 346259 99331
rect 346259 99297 346268 99331
rect 346216 99288 346268 99297
rect 357256 99331 357308 99340
rect 357256 99297 357265 99331
rect 357265 99297 357299 99331
rect 357299 99297 357308 99331
rect 357256 99288 357308 99297
rect 403532 99288 403584 99340
rect 424692 99331 424744 99340
rect 424692 99297 424701 99331
rect 424701 99297 424735 99331
rect 424735 99297 424744 99331
rect 424692 99288 424744 99297
rect 198280 98676 198332 98728
rect 198280 98540 198332 98592
rect 263784 96883 263836 96892
rect 263784 96849 263793 96883
rect 263793 96849 263827 96883
rect 263827 96849 263836 96883
rect 263784 96840 263836 96849
rect 154764 96747 154816 96756
rect 154764 96713 154773 96747
rect 154773 96713 154807 96747
rect 154807 96713 154816 96747
rect 154764 96704 154816 96713
rect 178224 96679 178276 96688
rect 178224 96645 178233 96679
rect 178233 96645 178267 96679
rect 178267 96645 178276 96679
rect 178224 96636 178276 96645
rect 154764 96568 154816 96620
rect 154948 96568 155000 96620
rect 162860 96568 162912 96620
rect 163044 96568 163096 96620
rect 303620 96568 303672 96620
rect 303712 96568 303764 96620
rect 384672 96568 384724 96620
rect 384856 96568 384908 96620
rect 403256 96568 403308 96620
rect 403532 96568 403584 96620
rect 423036 96568 423088 96620
rect 423128 96568 423180 96620
rect 168840 95251 168892 95260
rect 168840 95217 168849 95251
rect 168849 95217 168883 95251
rect 168883 95217 168892 95251
rect 168840 95208 168892 95217
rect 207112 95208 207164 95260
rect 224040 95208 224092 95260
rect 238668 95251 238720 95260
rect 238668 95217 238677 95251
rect 238677 95217 238711 95251
rect 238711 95217 238720 95251
rect 238668 95208 238720 95217
rect 248328 95251 248380 95260
rect 248328 95217 248337 95251
rect 248337 95217 248371 95251
rect 248371 95217 248380 95251
rect 248328 95208 248380 95217
rect 374276 95251 374328 95260
rect 374276 95217 374285 95251
rect 374285 95217 374319 95251
rect 374319 95217 374328 95251
rect 374276 95208 374328 95217
rect 188988 95183 189040 95192
rect 188988 95149 188997 95183
rect 188997 95149 189031 95183
rect 189031 95149 189040 95183
rect 188988 95140 189040 95149
rect 211344 95183 211396 95192
rect 211344 95149 211353 95183
rect 211353 95149 211387 95183
rect 211387 95149 211396 95183
rect 211344 95140 211396 95149
rect 216864 95183 216916 95192
rect 216864 95149 216873 95183
rect 216873 95149 216907 95183
rect 216907 95149 216916 95183
rect 216864 95140 216916 95149
rect 218336 95183 218388 95192
rect 218336 95149 218345 95183
rect 218345 95149 218379 95183
rect 218379 95149 218388 95183
rect 218336 95140 218388 95149
rect 219624 95183 219676 95192
rect 219624 95149 219633 95183
rect 219633 95149 219667 95183
rect 219667 95149 219676 95183
rect 219624 95140 219676 95149
rect 207204 95072 207256 95124
rect 208768 95072 208820 95124
rect 206008 93891 206060 93900
rect 206008 93857 206017 93891
rect 206017 93857 206051 93891
rect 206051 93857 206060 93891
rect 206008 93848 206060 93857
rect 270592 93848 270644 93900
rect 272064 93891 272116 93900
rect 272064 93857 272073 93891
rect 272073 93857 272107 93891
rect 272107 93857 272116 93891
rect 272064 93848 272116 93857
rect 226616 93823 226668 93832
rect 226616 93789 226625 93823
rect 226625 93789 226659 93823
rect 226659 93789 226668 93823
rect 226616 93780 226668 93789
rect 152004 92531 152056 92540
rect 152004 92497 152013 92531
rect 152013 92497 152047 92531
rect 152047 92497 152056 92531
rect 152004 92488 152056 92497
rect 192024 92488 192076 92540
rect 192116 92488 192168 92540
rect 226616 92531 226668 92540
rect 226616 92497 226625 92531
rect 226625 92497 226659 92531
rect 226659 92497 226668 92531
rect 226616 92488 226668 92497
rect 150716 92420 150768 92472
rect 150992 92420 151044 92472
rect 168472 91740 168524 91792
rect 168840 91740 168892 91792
rect 190644 91740 190696 91792
rect 190828 91740 190880 91792
rect 245936 90380 245988 90432
rect 173900 89700 173952 89752
rect 174084 89700 174136 89752
rect 252652 89700 252704 89752
rect 252836 89700 252888 89752
rect 264980 89700 265032 89752
rect 284300 89700 284352 89752
rect 284484 89700 284536 89752
rect 307852 89700 307904 89752
rect 308036 89700 308088 89752
rect 346124 89700 346176 89752
rect 346308 89700 346360 89752
rect 357164 89700 357216 89752
rect 357348 89700 357400 89752
rect 265072 89632 265124 89684
rect 379152 89403 379204 89412
rect 379152 89369 379161 89403
rect 379161 89369 379195 89403
rect 379195 89369 379204 89403
rect 379152 89360 379204 89369
rect 189080 86980 189132 87032
rect 206008 87023 206060 87032
rect 206008 86989 206017 87023
rect 206017 86989 206051 87023
rect 206051 86989 206060 87023
rect 206008 86980 206060 86989
rect 229192 86980 229244 87032
rect 229284 86980 229336 87032
rect 236184 86980 236236 87032
rect 236276 86980 236328 87032
rect 169852 86912 169904 86964
rect 173992 86955 174044 86964
rect 173992 86921 174001 86955
rect 174001 86921 174035 86955
rect 174035 86921 174044 86955
rect 173992 86912 174044 86921
rect 178224 86955 178276 86964
rect 178224 86921 178233 86955
rect 178233 86921 178267 86955
rect 178267 86921 178276 86955
rect 178224 86912 178276 86921
rect 190644 86955 190696 86964
rect 190644 86921 190653 86955
rect 190653 86921 190687 86955
rect 190687 86921 190696 86955
rect 190644 86912 190696 86921
rect 191932 86955 191984 86964
rect 191932 86921 191941 86955
rect 191941 86921 191975 86955
rect 191975 86921 191984 86955
rect 191932 86912 191984 86921
rect 222476 86912 222528 86964
rect 222568 86912 222620 86964
rect 223764 86912 223816 86964
rect 223856 86912 223908 86964
rect 247132 86912 247184 86964
rect 252744 86955 252796 86964
rect 252744 86921 252753 86955
rect 252753 86921 252787 86955
rect 252787 86921 252796 86955
rect 252744 86912 252796 86921
rect 258172 86912 258224 86964
rect 284392 86955 284444 86964
rect 284392 86921 284401 86955
rect 284401 86921 284435 86955
rect 284435 86921 284444 86955
rect 284392 86912 284444 86921
rect 307944 86955 307996 86964
rect 307944 86921 307953 86955
rect 307953 86921 307987 86955
rect 307987 86921 307996 86955
rect 307944 86912 307996 86921
rect 346216 86955 346268 86964
rect 346216 86921 346225 86955
rect 346225 86921 346259 86955
rect 346259 86921 346268 86955
rect 346216 86912 346268 86921
rect 357256 86955 357308 86964
rect 357256 86921 357265 86955
rect 357265 86921 357299 86955
rect 357299 86921 357308 86955
rect 357256 86912 357308 86921
rect 423220 86912 423272 86964
rect 423404 86912 423456 86964
rect 424692 86955 424744 86964
rect 424692 86921 424701 86955
rect 424701 86921 424735 86955
rect 424735 86921 424744 86955
rect 424692 86912 424744 86921
rect 189080 86844 189132 86896
rect 189172 85552 189224 85604
rect 194692 85552 194744 85604
rect 194784 85552 194836 85604
rect 206008 85595 206060 85604
rect 206008 85561 206017 85595
rect 206017 85561 206051 85595
rect 206051 85561 206060 85595
rect 206008 85552 206060 85561
rect 207020 85552 207072 85604
rect 207204 85552 207256 85604
rect 211344 85595 211396 85604
rect 211344 85561 211353 85595
rect 211353 85561 211387 85595
rect 211387 85561 211396 85595
rect 211344 85552 211396 85561
rect 216864 85595 216916 85604
rect 216864 85561 216873 85595
rect 216873 85561 216907 85595
rect 216907 85561 216916 85595
rect 216864 85552 216916 85561
rect 218336 85595 218388 85604
rect 218336 85561 218345 85595
rect 218345 85561 218379 85595
rect 218379 85561 218388 85595
rect 218336 85552 218388 85561
rect 219624 85595 219676 85604
rect 219624 85561 219633 85595
rect 219633 85561 219667 85595
rect 219667 85561 219676 85595
rect 219624 85552 219676 85561
rect 162952 85527 163004 85536
rect 162952 85493 162961 85527
rect 162961 85493 162995 85527
rect 162995 85493 163004 85527
rect 162952 85484 163004 85493
rect 223764 85527 223816 85536
rect 223764 85493 223773 85527
rect 223773 85493 223807 85527
rect 223807 85493 223816 85527
rect 223764 85484 223816 85493
rect 229192 85484 229244 85536
rect 238668 85527 238720 85536
rect 238668 85493 238677 85527
rect 238677 85493 238711 85527
rect 238711 85493 238720 85527
rect 238668 85484 238720 85493
rect 248328 85527 248380 85536
rect 248328 85493 248337 85527
rect 248337 85493 248371 85527
rect 248371 85493 248380 85527
rect 248328 85484 248380 85493
rect 270500 85527 270552 85536
rect 270500 85493 270509 85527
rect 270509 85493 270543 85527
rect 270543 85493 270552 85527
rect 270500 85484 270552 85493
rect 272064 85527 272116 85536
rect 272064 85493 272073 85527
rect 272073 85493 272107 85527
rect 272107 85493 272116 85527
rect 272064 85484 272116 85493
rect 374276 85527 374328 85536
rect 374276 85493 374285 85527
rect 374285 85493 374319 85527
rect 374319 85493 374328 85527
rect 374276 85484 374328 85493
rect 229376 85416 229428 85468
rect 194784 84124 194836 84176
rect 207020 84167 207072 84176
rect 207020 84133 207029 84167
rect 207029 84133 207063 84167
rect 207063 84133 207072 84167
rect 207020 84124 207072 84133
rect 208584 84124 208636 84176
rect 246212 83172 246264 83224
rect 152004 82807 152056 82816
rect 152004 82773 152013 82807
rect 152013 82773 152047 82807
rect 152047 82773 152056 82807
rect 152004 82764 152056 82773
rect 226616 82764 226668 82816
rect 190644 80699 190696 80708
rect 190644 80665 190653 80699
rect 190653 80665 190687 80699
rect 190687 80665 190696 80699
rect 190644 80656 190696 80665
rect 403440 80044 403492 80096
rect 403532 79908 403584 79960
rect 168472 77324 168524 77376
rect 168656 77324 168708 77376
rect 169760 77299 169812 77308
rect 169760 77265 169769 77299
rect 169769 77265 169803 77299
rect 169803 77265 169812 77299
rect 169760 77256 169812 77265
rect 174084 77256 174136 77308
rect 178224 77299 178276 77308
rect 178224 77265 178233 77299
rect 178233 77265 178267 77299
rect 178267 77265 178276 77299
rect 178224 77256 178276 77265
rect 234712 77256 234764 77308
rect 234804 77256 234856 77308
rect 236184 77256 236236 77308
rect 236276 77256 236328 77308
rect 237472 77256 237524 77308
rect 237564 77256 237616 77308
rect 247040 77299 247092 77308
rect 247040 77265 247049 77299
rect 247049 77265 247083 77299
rect 247083 77265 247092 77299
rect 247040 77256 247092 77265
rect 252836 77256 252888 77308
rect 258080 77299 258132 77308
rect 258080 77265 258089 77299
rect 258089 77265 258123 77299
rect 258123 77265 258132 77299
rect 258080 77256 258132 77265
rect 265072 77256 265124 77308
rect 284484 77256 284536 77308
rect 308036 77256 308088 77308
rect 346308 77256 346360 77308
rect 357348 77256 357400 77308
rect 424784 77256 424836 77308
rect 154764 77231 154816 77240
rect 154764 77197 154773 77231
rect 154773 77197 154807 77231
rect 154807 77197 154816 77231
rect 154764 77188 154816 77197
rect 303896 77231 303948 77240
rect 303896 77197 303905 77231
rect 303905 77197 303939 77231
rect 303939 77197 303948 77231
rect 303896 77188 303948 77197
rect 577688 77188 577740 77240
rect 579620 77188 579672 77240
rect 265072 77120 265124 77172
rect 357348 77120 357400 77172
rect 198280 75964 198332 76016
rect 163228 75896 163280 75948
rect 192024 75896 192076 75948
rect 198188 75896 198240 75948
rect 238668 75939 238720 75948
rect 238668 75905 238677 75939
rect 238677 75905 238711 75939
rect 238711 75905 238720 75939
rect 238668 75896 238720 75905
rect 248328 75939 248380 75948
rect 248328 75905 248337 75939
rect 248337 75905 248371 75939
rect 248371 75905 248380 75939
rect 248328 75896 248380 75905
rect 270592 75896 270644 75948
rect 272064 75939 272116 75948
rect 272064 75905 272073 75939
rect 272073 75905 272107 75939
rect 272107 75905 272116 75939
rect 272064 75896 272116 75905
rect 374276 75939 374328 75948
rect 374276 75905 374285 75939
rect 374285 75905 374319 75939
rect 374319 75905 374328 75939
rect 374276 75896 374328 75905
rect 196256 75828 196308 75880
rect 196348 75828 196400 75880
rect 384672 75871 384724 75880
rect 384672 75837 384681 75871
rect 384681 75837 384715 75871
rect 384715 75837 384724 75871
rect 384672 75828 384724 75837
rect 194784 74536 194836 74588
rect 223764 74579 223816 74588
rect 223764 74545 223773 74579
rect 223773 74545 223807 74579
rect 223807 74545 223816 74579
rect 223764 74536 223816 74545
rect 198188 74468 198240 74520
rect 198280 74468 198332 74520
rect 211252 74511 211304 74520
rect 211252 74477 211261 74511
rect 211261 74477 211295 74511
rect 211295 74477 211304 74511
rect 211252 74468 211304 74477
rect 246212 74468 246264 74520
rect 152004 73219 152056 73228
rect 152004 73185 152013 73219
rect 152013 73185 152047 73219
rect 152047 73185 152056 73219
rect 152004 73176 152056 73185
rect 190644 70499 190696 70508
rect 190644 70465 190653 70499
rect 190653 70465 190687 70499
rect 190687 70465 190696 70499
rect 190644 70456 190696 70465
rect 192024 70456 192076 70508
rect 194784 70456 194836 70508
rect 216864 70456 216916 70508
rect 219624 70524 219676 70576
rect 346124 70388 346176 70440
rect 191932 70320 191984 70372
rect 194692 70320 194744 70372
rect 216772 70320 216824 70372
rect 219532 70320 219584 70372
rect 346216 70320 346268 70372
rect 150716 70295 150768 70304
rect 150716 70261 150725 70295
rect 150725 70261 150759 70295
rect 150759 70261 150768 70295
rect 150716 70252 150768 70261
rect 303896 70227 303948 70236
rect 303896 70193 303905 70227
rect 303905 70193 303939 70227
rect 303939 70193 303948 70227
rect 303896 70184 303948 70193
rect 248328 67736 248380 67788
rect 265072 67736 265124 67788
rect 162952 67668 163004 67720
rect 163228 67668 163280 67720
rect 252836 67668 252888 67720
rect 307944 67668 307996 67720
rect 308036 67668 308088 67720
rect 154764 67643 154816 67652
rect 154764 67609 154773 67643
rect 154773 67609 154807 67643
rect 154807 67609 154816 67643
rect 154764 67600 154816 67609
rect 173992 67600 174044 67652
rect 174084 67600 174136 67652
rect 222476 67600 222528 67652
rect 222568 67600 222620 67652
rect 248328 67600 248380 67652
rect 265072 67600 265124 67652
rect 357256 67643 357308 67652
rect 357256 67609 357265 67643
rect 357265 67609 357299 67643
rect 357299 67609 357308 67643
rect 357256 67600 357308 67609
rect 423220 67600 423272 67652
rect 423312 67600 423364 67652
rect 236276 67532 236328 67584
rect 236368 67532 236420 67584
rect 237564 67532 237616 67584
rect 237656 67532 237708 67584
rect 307668 67532 307720 67584
rect 307944 67532 307996 67584
rect 424692 67575 424744 67584
rect 424692 67541 424701 67575
rect 424701 67541 424735 67575
rect 424735 67541 424744 67575
rect 424692 67532 424744 67541
rect 208492 66351 208544 66360
rect 208492 66317 208501 66351
rect 208501 66317 208535 66351
rect 208535 66317 208544 66351
rect 208492 66308 208544 66317
rect 190644 66283 190696 66292
rect 190644 66249 190653 66283
rect 190653 66249 190687 66283
rect 190687 66249 190696 66283
rect 190644 66240 190696 66249
rect 207112 66240 207164 66292
rect 252744 66283 252796 66292
rect 252744 66249 252753 66283
rect 252753 66249 252787 66283
rect 252787 66249 252796 66283
rect 252744 66240 252796 66249
rect 284392 66240 284444 66292
rect 284484 66240 284536 66292
rect 384764 66240 384816 66292
rect 162952 66172 163004 66224
rect 168564 66172 168616 66224
rect 191932 66172 191984 66224
rect 192116 66172 192168 66224
rect 219532 66215 219584 66224
rect 219532 66181 219541 66215
rect 219541 66181 219575 66215
rect 219575 66181 219584 66215
rect 219532 66172 219584 66181
rect 238668 66215 238720 66224
rect 238668 66181 238677 66215
rect 238677 66181 238711 66215
rect 238711 66181 238720 66215
rect 238668 66172 238720 66181
rect 248328 66215 248380 66224
rect 248328 66181 248337 66215
rect 248337 66181 248371 66215
rect 248371 66181 248380 66215
rect 248328 66172 248380 66181
rect 263784 66172 263836 66224
rect 265072 66215 265124 66224
rect 265072 66181 265081 66215
rect 265081 66181 265115 66215
rect 265115 66181 265124 66215
rect 265072 66172 265124 66181
rect 374276 66215 374328 66224
rect 374276 66181 374285 66215
rect 374285 66181 374319 66215
rect 374319 66181 374328 66215
rect 374276 66172 374328 66181
rect 379152 66215 379204 66224
rect 379152 66181 379161 66215
rect 379161 66181 379195 66215
rect 379195 66181 379204 66215
rect 379152 66172 379204 66181
rect 211344 64948 211396 65000
rect 246028 64923 246080 64932
rect 246028 64889 246037 64923
rect 246037 64889 246071 64923
rect 246071 64889 246080 64923
rect 246028 64880 246080 64889
rect 3332 64812 3384 64864
rect 21364 64812 21416 64864
rect 150716 64855 150768 64864
rect 150716 64821 150725 64855
rect 150725 64821 150759 64855
rect 150759 64821 150768 64855
rect 150716 64812 150768 64821
rect 189172 64855 189224 64864
rect 189172 64821 189181 64855
rect 189181 64821 189215 64855
rect 189215 64821 189224 64855
rect 189172 64812 189224 64821
rect 207112 64855 207164 64864
rect 207112 64821 207121 64855
rect 207121 64821 207155 64855
rect 207155 64821 207164 64855
rect 207112 64812 207164 64821
rect 208492 64855 208544 64864
rect 208492 64821 208501 64855
rect 208501 64821 208535 64855
rect 208535 64821 208544 64855
rect 208492 64812 208544 64821
rect 211344 64855 211396 64864
rect 211344 64821 211353 64855
rect 211353 64821 211387 64855
rect 211387 64821 211396 64855
rect 211344 64812 211396 64821
rect 218244 64855 218296 64864
rect 218244 64821 218253 64855
rect 218253 64821 218287 64855
rect 218287 64821 218296 64855
rect 218244 64812 218296 64821
rect 223764 64812 223816 64864
rect 577596 64676 577648 64728
rect 580356 64676 580408 64728
rect 190644 64651 190696 64660
rect 190644 64617 190653 64651
rect 190653 64617 190687 64651
rect 190687 64617 190696 64651
rect 190644 64608 190696 64617
rect 198188 63495 198240 63504
rect 198188 63461 198197 63495
rect 198197 63461 198231 63495
rect 198231 63461 198240 63495
rect 198188 63452 198240 63461
rect 177948 62772 178000 62824
rect 178224 62772 178276 62824
rect 403440 62092 403492 62144
rect 403532 62092 403584 62144
rect 284392 60800 284444 60852
rect 169852 60664 169904 60716
rect 170036 60664 170088 60716
rect 258172 60664 258224 60716
rect 258356 60664 258408 60716
rect 265072 60707 265124 60716
rect 265072 60673 265081 60707
rect 265081 60673 265115 60707
rect 265115 60673 265124 60707
rect 265072 60664 265124 60673
rect 278872 60664 278924 60716
rect 284392 60664 284444 60716
rect 278964 60596 279016 60648
rect 252468 58012 252520 58064
rect 423220 58012 423272 58064
rect 423496 58012 423548 58064
rect 214104 57944 214156 57996
rect 214196 57944 214248 57996
rect 229284 57944 229336 57996
rect 229376 57944 229428 57996
rect 303620 57944 303672 57996
rect 303896 57944 303948 57996
rect 424784 57944 424836 57996
rect 154764 57919 154816 57928
rect 154764 57885 154773 57919
rect 154773 57885 154807 57919
rect 154807 57885 154816 57919
rect 154764 57876 154816 57885
rect 174084 57876 174136 57928
rect 178224 57919 178276 57928
rect 178224 57885 178233 57919
rect 178233 57885 178267 57919
rect 178267 57885 178276 57919
rect 178224 57876 178276 57885
rect 252468 57876 252520 57928
rect 258356 57876 258408 57928
rect 307852 57919 307904 57928
rect 307852 57885 307861 57919
rect 307861 57885 307895 57919
rect 307895 57885 307904 57919
rect 307852 57876 307904 57885
rect 357348 57876 357400 57928
rect 252376 56992 252428 57044
rect 252836 56992 252888 57044
rect 162860 56627 162912 56636
rect 162860 56593 162869 56627
rect 162869 56593 162903 56627
rect 162903 56593 162912 56627
rect 168472 56627 168524 56636
rect 162860 56584 162912 56593
rect 168472 56593 168481 56627
rect 168481 56593 168515 56627
rect 168515 56593 168524 56627
rect 168472 56584 168524 56593
rect 190736 56584 190788 56636
rect 246028 56652 246080 56704
rect 379152 56695 379204 56704
rect 379152 56661 379161 56695
rect 379161 56661 379195 56695
rect 379195 56661 379204 56695
rect 379152 56652 379204 56661
rect 247132 56584 247184 56636
rect 247316 56584 247368 56636
rect 248328 56627 248380 56636
rect 248328 56593 248337 56627
rect 248337 56593 248371 56627
rect 248371 56593 248380 56627
rect 248328 56584 248380 56593
rect 374276 56627 374328 56636
rect 374276 56593 374285 56627
rect 374285 56593 374319 56627
rect 374319 56593 374328 56627
rect 374276 56584 374328 56593
rect 216864 56516 216916 56568
rect 216956 56516 217008 56568
rect 245844 56516 245896 56568
rect 379152 56559 379204 56568
rect 379152 56525 379161 56559
rect 379161 56525 379195 56559
rect 379195 56525 379204 56559
rect 379152 56516 379204 56525
rect 207112 56355 207164 56364
rect 207112 56321 207121 56355
rect 207121 56321 207155 56355
rect 207155 56321 207164 56355
rect 207112 56312 207164 56321
rect 192116 55292 192168 55344
rect 194692 55267 194744 55276
rect 194692 55233 194701 55267
rect 194701 55233 194735 55267
rect 194735 55233 194744 55267
rect 194692 55224 194744 55233
rect 208492 55267 208544 55276
rect 208492 55233 208501 55267
rect 208501 55233 208535 55267
rect 208535 55233 208544 55267
rect 208492 55224 208544 55233
rect 211528 55224 211580 55276
rect 223672 55267 223724 55276
rect 223672 55233 223681 55267
rect 223681 55233 223715 55267
rect 223715 55233 223724 55267
rect 223672 55224 223724 55233
rect 226708 55224 226760 55276
rect 216956 55199 217008 55208
rect 216956 55165 216965 55199
rect 216965 55165 216999 55199
rect 216999 55165 217008 55199
rect 216956 55156 217008 55165
rect 192024 53839 192076 53848
rect 192024 53805 192033 53839
rect 192033 53805 192067 53839
rect 192067 53805 192076 53839
rect 192024 53796 192076 53805
rect 194692 53839 194744 53848
rect 194692 53805 194701 53839
rect 194701 53805 194735 53839
rect 194735 53805 194744 53839
rect 194692 53796 194744 53805
rect 198188 53839 198240 53848
rect 198188 53805 198197 53839
rect 198197 53805 198231 53839
rect 198231 53805 198240 53839
rect 198188 53796 198240 53805
rect 403624 52436 403676 52488
rect 403716 52436 403768 52488
rect 179512 51144 179564 51196
rect 270592 51187 270644 51196
rect 270592 51153 270601 51187
rect 270601 51153 270635 51187
rect 270635 51153 270644 51187
rect 270592 51144 270644 51153
rect 196256 51076 196308 51128
rect 272064 51076 272116 51128
rect 284392 51076 284444 51128
rect 179512 51008 179564 51060
rect 196164 51008 196216 51060
rect 252376 51008 252428 51060
rect 252744 51008 252796 51060
rect 284300 51008 284352 51060
rect 154764 48399 154816 48408
rect 154764 48365 154773 48399
rect 154773 48365 154807 48399
rect 154807 48365 154816 48399
rect 154764 48356 154816 48365
rect 173992 48331 174044 48340
rect 173992 48297 174001 48331
rect 174001 48297 174035 48331
rect 174035 48297 174044 48331
rect 173992 48288 174044 48297
rect 178316 48288 178368 48340
rect 190644 48288 190696 48340
rect 190736 48288 190788 48340
rect 238668 48331 238720 48340
rect 238668 48297 238677 48331
rect 238677 48297 238711 48331
rect 238711 48297 238720 48331
rect 238668 48288 238720 48297
rect 258172 48331 258224 48340
rect 258172 48297 258181 48331
rect 258181 48297 258215 48331
rect 258215 48297 258224 48331
rect 258172 48288 258224 48297
rect 263692 48331 263744 48340
rect 263692 48297 263701 48331
rect 263701 48297 263735 48331
rect 263735 48297 263744 48331
rect 263692 48288 263744 48297
rect 270592 48331 270644 48340
rect 270592 48297 270601 48331
rect 270601 48297 270635 48331
rect 270635 48297 270644 48331
rect 270592 48288 270644 48297
rect 271880 48331 271932 48340
rect 271880 48297 271889 48331
rect 271889 48297 271923 48331
rect 271923 48297 271932 48331
rect 271880 48288 271932 48297
rect 307944 48288 307996 48340
rect 346216 48288 346268 48340
rect 346308 48288 346360 48340
rect 357256 48331 357308 48340
rect 357256 48297 357265 48331
rect 357265 48297 357299 48331
rect 357299 48297 357308 48331
rect 357256 48288 357308 48297
rect 384764 48288 384816 48340
rect 384856 48288 384908 48340
rect 403716 48288 403768 48340
rect 403808 48288 403860 48340
rect 154764 48263 154816 48272
rect 154764 48229 154773 48263
rect 154773 48229 154807 48263
rect 154807 48229 154816 48263
rect 154764 48220 154816 48229
rect 225052 48220 225104 48272
rect 225144 48220 225196 48272
rect 234896 48220 234948 48272
rect 236276 48220 236328 48272
rect 236368 48220 236420 48272
rect 237564 48220 237616 48272
rect 237656 48220 237708 48272
rect 284300 48220 284352 48272
rect 424692 48263 424744 48272
rect 424692 48229 424701 48263
rect 424701 48229 424735 48263
rect 424735 48229 424744 48263
rect 424692 48220 424744 48229
rect 211528 47268 211580 47320
rect 189356 46928 189408 46980
rect 218244 46971 218296 46980
rect 218244 46937 218253 46971
rect 218253 46937 218287 46971
rect 218287 46937 218296 46971
rect 218244 46928 218296 46937
rect 219532 46971 219584 46980
rect 219532 46937 219541 46971
rect 219541 46937 219575 46971
rect 219575 46937 219584 46971
rect 219532 46928 219584 46937
rect 379244 46928 379296 46980
rect 168564 46903 168616 46912
rect 168564 46869 168573 46903
rect 168573 46869 168607 46903
rect 168607 46869 168616 46903
rect 168564 46860 168616 46869
rect 169852 46903 169904 46912
rect 169852 46869 169861 46903
rect 169861 46869 169895 46903
rect 169895 46869 169904 46903
rect 169852 46860 169904 46869
rect 207112 46903 207164 46912
rect 207112 46869 207121 46903
rect 207121 46869 207155 46903
rect 207155 46869 207164 46903
rect 207112 46860 207164 46869
rect 214012 46860 214064 46912
rect 238668 46860 238720 46912
rect 245844 46860 245896 46912
rect 247132 46860 247184 46912
rect 247408 46860 247460 46912
rect 248328 46903 248380 46912
rect 248328 46869 248337 46903
rect 248337 46869 248371 46903
rect 248371 46869 248380 46903
rect 248328 46860 248380 46869
rect 374276 46903 374328 46912
rect 374276 46869 374285 46903
rect 374285 46869 374319 46903
rect 374319 46869 374328 46903
rect 374276 46860 374328 46869
rect 245752 46792 245804 46844
rect 194692 45772 194744 45824
rect 150532 45636 150584 45688
rect 150716 45636 150768 45688
rect 194784 45568 194836 45620
rect 211252 45611 211304 45620
rect 211252 45577 211261 45611
rect 211261 45577 211295 45611
rect 211295 45577 211304 45611
rect 211252 45568 211304 45577
rect 216956 45611 217008 45620
rect 216956 45577 216965 45611
rect 216965 45577 216999 45611
rect 216999 45577 217008 45611
rect 216956 45568 217008 45577
rect 196164 45500 196216 45552
rect 196348 45500 196400 45552
rect 218244 45500 218296 45552
rect 218336 45500 218388 45552
rect 219532 45500 219584 45552
rect 245752 45543 245804 45552
rect 245752 45509 245761 45543
rect 245761 45509 245795 45543
rect 245795 45509 245804 45543
rect 245752 45500 245804 45509
rect 247408 45543 247460 45552
rect 247408 45509 247417 45543
rect 247417 45509 247451 45543
rect 247451 45509 247460 45543
rect 247408 45500 247460 45509
rect 155040 43664 155092 43716
rect 208584 42075 208636 42084
rect 208584 42041 208593 42075
rect 208593 42041 208627 42075
rect 208627 42041 208636 42075
rect 208584 42032 208636 42041
rect 222476 42075 222528 42084
rect 222476 42041 222485 42075
rect 222485 42041 222519 42075
rect 222519 42041 222528 42075
rect 222476 42032 222528 42041
rect 223764 42075 223816 42084
rect 223764 42041 223773 42075
rect 223773 42041 223807 42075
rect 223807 42041 223816 42075
rect 223764 42032 223816 42041
rect 178132 41352 178184 41404
rect 178316 41352 178368 41404
rect 284484 41395 284536 41404
rect 284484 41361 284493 41395
rect 284493 41361 284527 41395
rect 284527 41361 284536 41395
rect 284484 41352 284536 41361
rect 340696 40196 340748 40248
rect 340972 40196 341024 40248
rect 201500 40128 201552 40180
rect 219348 40128 219400 40180
rect 321284 40128 321336 40180
rect 321560 40128 321612 40180
rect 359924 40128 359976 40180
rect 360200 40128 360252 40180
rect 444380 40060 444432 40112
rect 447232 40060 447284 40112
rect 476028 40060 476080 40112
rect 482928 40060 482980 40112
rect 258264 38768 258316 38820
rect 423312 38700 423364 38752
rect 423496 38700 423548 38752
rect 189264 38632 189316 38684
rect 189356 38632 189408 38684
rect 190644 38632 190696 38684
rect 190736 38632 190788 38684
rect 234804 38675 234856 38684
rect 234804 38641 234813 38675
rect 234813 38641 234847 38675
rect 234847 38641 234856 38675
rect 234804 38632 234856 38641
rect 252652 38632 252704 38684
rect 252836 38632 252888 38684
rect 258264 38632 258316 38684
rect 264980 38632 265032 38684
rect 265072 38632 265124 38684
rect 384672 38632 384724 38684
rect 384764 38632 384816 38684
rect 424784 38632 424836 38684
rect 284484 38564 284536 38616
rect 308036 38564 308088 38616
rect 357348 38564 357400 38616
rect 403808 38607 403860 38616
rect 403808 38573 403817 38607
rect 403817 38573 403851 38607
rect 403851 38573 403860 38607
rect 403808 38564 403860 38573
rect 168656 37272 168708 37324
rect 169944 37272 169996 37324
rect 190736 37204 190788 37256
rect 238668 37272 238720 37324
rect 248328 37315 248380 37324
rect 248328 37281 248337 37315
rect 248337 37281 248371 37315
rect 248371 37281 248380 37315
rect 248328 37272 248380 37281
rect 374276 37315 374328 37324
rect 374276 37281 374285 37315
rect 374285 37281 374319 37315
rect 374319 37281 374328 37315
rect 374276 37272 374328 37281
rect 379152 37272 379204 37324
rect 379244 37272 379296 37324
rect 219532 37204 219584 37256
rect 247408 37247 247460 37256
rect 247408 37213 247417 37247
rect 247417 37213 247451 37247
rect 247451 37213 247460 37247
rect 247408 37204 247460 37213
rect 194508 34484 194560 34536
rect 194692 34484 194744 34536
rect 174084 33804 174136 33856
rect 213920 32376 213972 32428
rect 270592 31875 270644 31884
rect 270592 31841 270601 31875
rect 270601 31841 270635 31875
rect 270635 31841 270644 31875
rect 270592 31832 270644 31841
rect 273352 31875 273404 31884
rect 273352 31841 273361 31875
rect 273361 31841 273395 31875
rect 273395 31841 273404 31875
rect 273352 31832 273404 31841
rect 168656 31764 168708 31816
rect 169944 31764 169996 31816
rect 346124 31764 346176 31816
rect 168748 31628 168800 31680
rect 169944 31628 169996 31680
rect 357256 31739 357308 31748
rect 357256 31705 357265 31739
rect 357265 31705 357299 31739
rect 357299 31705 357308 31739
rect 357256 31696 357308 31705
rect 379336 31764 379388 31816
rect 423312 31764 423364 31816
rect 424784 31764 424836 31816
rect 424968 31764 425020 31816
rect 384672 31696 384724 31748
rect 384856 31696 384908 31748
rect 393964 31696 394016 31748
rect 394148 31696 394200 31748
rect 346216 31628 346268 31680
rect 379244 31628 379296 31680
rect 423404 31628 423456 31680
rect 247408 31331 247460 31340
rect 247408 31297 247417 31331
rect 247417 31297 247451 31331
rect 247451 31297 247460 31331
rect 247408 31288 247460 31297
rect 178316 31220 178368 31272
rect 178316 31084 178368 31136
rect 577504 30268 577556 30320
rect 579620 30268 579672 30320
rect 179604 29044 179656 29096
rect 236276 29044 236328 29096
rect 264980 29044 265032 29096
rect 265072 29044 265124 29096
rect 173992 29019 174044 29028
rect 173992 28985 174001 29019
rect 174001 28985 174035 29019
rect 174035 28985 174044 29019
rect 173992 28976 174044 28985
rect 179512 28976 179564 29028
rect 205732 28976 205784 29028
rect 205824 28976 205876 29028
rect 208584 29019 208636 29028
rect 208584 28985 208593 29019
rect 208593 28985 208627 29019
rect 208627 28985 208636 29019
rect 208584 28976 208636 28985
rect 222660 28976 222712 29028
rect 223764 29019 223816 29028
rect 223764 28985 223773 29019
rect 223773 28985 223807 29019
rect 223807 28985 223816 29019
rect 223764 28976 223816 28985
rect 229376 28976 229428 29028
rect 229468 28976 229520 29028
rect 236184 28976 236236 29028
rect 238668 29019 238720 29028
rect 238668 28985 238677 29019
rect 238677 28985 238711 29019
rect 238711 28985 238720 29019
rect 238668 28976 238720 28985
rect 284392 29019 284444 29028
rect 284392 28985 284401 29019
rect 284401 28985 284435 29019
rect 284435 28985 284444 29019
rect 284392 28976 284444 28985
rect 307944 29019 307996 29028
rect 307944 28985 307953 29019
rect 307953 28985 307987 29019
rect 307987 28985 307996 29019
rect 307944 28976 307996 28985
rect 403900 28976 403952 29028
rect 271972 28908 272024 28960
rect 272064 28908 272116 28960
rect 394148 28908 394200 28960
rect 150532 28296 150584 28348
rect 150716 28296 150768 28348
rect 190644 27727 190696 27736
rect 190644 27693 190653 27727
rect 190653 27693 190687 27727
rect 190687 27693 190696 27727
rect 190644 27684 190696 27693
rect 207112 27684 207164 27736
rect 238668 27727 238720 27736
rect 238668 27693 238677 27727
rect 238677 27693 238711 27727
rect 238711 27693 238720 27727
rect 238668 27684 238720 27693
rect 191932 27659 191984 27668
rect 191932 27625 191941 27659
rect 191941 27625 191975 27659
rect 191975 27625 191984 27659
rect 191932 27616 191984 27625
rect 198188 27616 198240 27668
rect 198280 27616 198332 27668
rect 245844 27616 245896 27668
rect 247408 27659 247460 27668
rect 247408 27625 247417 27659
rect 247417 27625 247451 27659
rect 247451 27625 247460 27659
rect 247408 27616 247460 27625
rect 270592 27659 270644 27668
rect 270592 27625 270601 27659
rect 270601 27625 270635 27659
rect 270635 27625 270644 27659
rect 270592 27616 270644 27625
rect 273352 27659 273404 27668
rect 273352 27625 273361 27659
rect 273361 27625 273395 27659
rect 273395 27625 273404 27659
rect 273352 27616 273404 27625
rect 168564 27548 168616 27600
rect 168748 27548 168800 27600
rect 173992 27591 174044 27600
rect 173992 27557 174001 27591
rect 174001 27557 174035 27591
rect 174035 27557 174044 27591
rect 173992 27548 174044 27557
rect 179512 27591 179564 27600
rect 179512 27557 179521 27591
rect 179521 27557 179555 27591
rect 179555 27557 179564 27591
rect 179512 27548 179564 27557
rect 205824 27548 205876 27600
rect 205916 27548 205968 27600
rect 207112 27591 207164 27600
rect 207112 27557 207121 27591
rect 207121 27557 207155 27591
rect 207155 27557 207164 27591
rect 207112 27548 207164 27557
rect 211252 27548 211304 27600
rect 223764 27548 223816 27600
rect 238668 27548 238720 27600
rect 252744 27591 252796 27600
rect 252744 27557 252753 27591
rect 252753 27557 252787 27591
rect 252787 27557 252796 27591
rect 252744 27548 252796 27557
rect 264980 27591 265032 27600
rect 264980 27557 264989 27591
rect 264989 27557 265023 27591
rect 265023 27557 265032 27591
rect 264980 27548 265032 27557
rect 346216 27591 346268 27600
rect 346216 27557 346225 27591
rect 346225 27557 346259 27591
rect 346259 27557 346268 27591
rect 346216 27548 346268 27557
rect 374276 27591 374328 27600
rect 374276 27557 374285 27591
rect 374285 27557 374319 27591
rect 374319 27557 374328 27591
rect 374276 27548 374328 27557
rect 384856 27548 384908 27600
rect 379244 27523 379296 27532
rect 379244 27489 379253 27523
rect 379253 27489 379287 27523
rect 379287 27489 379296 27523
rect 379244 27480 379296 27489
rect 245844 27251 245896 27260
rect 245844 27217 245853 27251
rect 245853 27217 245887 27251
rect 245887 27217 245896 27251
rect 245844 27208 245896 27217
rect 152004 26256 152056 26308
rect 152096 26256 152148 26308
rect 191932 26299 191984 26308
rect 191932 26265 191941 26299
rect 191941 26265 191975 26299
rect 191975 26265 191984 26299
rect 191932 26256 191984 26265
rect 189172 26231 189224 26240
rect 189172 26197 189181 26231
rect 189181 26197 189215 26231
rect 189215 26197 189224 26231
rect 189172 26188 189224 26197
rect 194692 26231 194744 26240
rect 194692 26197 194701 26231
rect 194701 26197 194735 26231
rect 194735 26197 194744 26231
rect 194692 26188 194744 26197
rect 190644 22108 190696 22160
rect 173992 22083 174044 22092
rect 173992 22049 174001 22083
rect 174001 22049 174035 22083
rect 174035 22049 174044 22083
rect 173992 22040 174044 22049
rect 198280 22108 198332 22160
rect 196164 22040 196216 22092
rect 196348 22040 196400 22092
rect 198188 22040 198240 22092
rect 346216 22083 346268 22092
rect 346216 22049 346225 22083
rect 346225 22049 346259 22083
rect 346259 22049 346268 22083
rect 346216 22040 346268 22049
rect 379336 22040 379388 22092
rect 190736 21972 190788 22024
rect 191748 21360 191800 21412
rect 218244 19388 218296 19440
rect 219532 19388 219584 19440
rect 211344 19363 211396 19372
rect 211344 19329 211353 19363
rect 211353 19329 211387 19363
rect 211387 19329 211396 19363
rect 211344 19320 211396 19329
rect 229284 19320 229336 19372
rect 229376 19320 229428 19372
rect 234712 19320 234764 19372
rect 234804 19320 234856 19372
rect 236184 19320 236236 19372
rect 236276 19320 236328 19372
rect 237472 19320 237524 19372
rect 237564 19320 237616 19372
rect 239036 19320 239088 19372
rect 239128 19320 239180 19372
rect 245936 19320 245988 19372
rect 270592 19320 270644 19372
rect 394056 19363 394108 19372
rect 394056 19329 394065 19363
rect 394065 19329 394099 19363
rect 394099 19329 394108 19363
rect 394056 19320 394108 19329
rect 403716 19320 403768 19372
rect 403808 19320 403860 19372
rect 218244 19252 218296 19304
rect 219532 19252 219584 19304
rect 248328 19252 248380 19304
rect 179512 18003 179564 18012
rect 179512 17969 179521 18003
rect 179521 17969 179555 18003
rect 179555 17969 179564 18003
rect 179512 17960 179564 17969
rect 207204 17960 207256 18012
rect 252836 17960 252888 18012
rect 265072 17960 265124 18012
rect 374276 18003 374328 18012
rect 374276 17969 374285 18003
rect 374285 17969 374319 18003
rect 374319 17969 374328 18003
rect 374276 17960 374328 17969
rect 384580 18003 384632 18012
rect 384580 17969 384589 18003
rect 384589 17969 384623 18003
rect 384623 17969 384632 18003
rect 384580 17960 384632 17969
rect 154856 17935 154908 17944
rect 154856 17901 154865 17935
rect 154865 17901 154899 17935
rect 154899 17901 154908 17935
rect 154856 17892 154908 17901
rect 338212 16804 338264 16856
rect 342628 16804 342680 16856
rect 359924 16804 359976 16856
rect 362224 16804 362276 16856
rect 379244 16804 379296 16856
rect 379612 16804 379664 16856
rect 318800 16736 318852 16788
rect 321560 16736 321612 16788
rect 398656 16736 398708 16788
rect 400864 16736 400916 16788
rect 417976 16736 418028 16788
rect 418252 16736 418304 16788
rect 173900 16668 173952 16720
rect 183468 16668 183520 16720
rect 444380 16668 444432 16720
rect 447232 16668 447284 16720
rect 476028 16668 476080 16720
rect 482928 16668 482980 16720
rect 189172 16643 189224 16652
rect 189172 16609 189181 16643
rect 189181 16609 189215 16643
rect 189215 16609 189224 16643
rect 189172 16600 189224 16609
rect 194692 16643 194744 16652
rect 194692 16609 194701 16643
rect 194701 16609 194735 16643
rect 194735 16609 194744 16643
rect 194692 16600 194744 16609
rect 190460 13472 190512 13524
rect 190736 13472 190788 13524
rect 374276 12520 374328 12572
rect 168564 12452 168616 12504
rect 216864 12452 216916 12504
rect 424784 12452 424836 12504
rect 424968 12452 425020 12504
rect 154856 12427 154908 12436
rect 154856 12393 154865 12427
rect 154865 12393 154899 12427
rect 154899 12393 154908 12427
rect 154856 12384 154908 12393
rect 168472 12384 168524 12436
rect 216772 12384 216824 12436
rect 356336 12384 356388 12436
rect 357440 12384 357492 12436
rect 358544 12384 358596 12436
rect 375564 12384 375616 12436
rect 376392 12384 376444 12436
rect 357348 12316 357400 12368
rect 169852 9664 169904 9716
rect 170128 9664 170180 9716
rect 191932 9707 191984 9716
rect 191932 9673 191941 9707
rect 191941 9673 191975 9707
rect 191975 9673 191984 9707
rect 191932 9664 191984 9673
rect 223672 9707 223724 9716
rect 223672 9673 223681 9707
rect 223681 9673 223715 9707
rect 223715 9673 223724 9707
rect 223672 9664 223724 9673
rect 238576 9707 238628 9716
rect 238576 9673 238585 9707
rect 238585 9673 238619 9707
rect 238619 9673 238628 9707
rect 238576 9664 238628 9673
rect 247960 9707 248012 9716
rect 247960 9673 247969 9707
rect 247969 9673 248003 9707
rect 248003 9673 248012 9707
rect 247960 9664 248012 9673
rect 270592 9664 270644 9716
rect 309416 9664 309468 9716
rect 309784 9664 309836 9716
rect 374184 9707 374236 9716
rect 374184 9673 374193 9707
rect 374193 9673 374227 9707
rect 374227 9673 374236 9707
rect 374184 9664 374236 9673
rect 384580 9664 384632 9716
rect 384856 9664 384908 9716
rect 109960 9596 110012 9648
rect 205824 9596 205876 9648
rect 106372 9528 106424 9580
rect 204352 9528 204404 9580
rect 102784 9460 102836 9512
rect 201592 9460 201644 9512
rect 383568 9460 383620 9512
rect 452476 9460 452528 9512
rect 95700 9392 95752 9444
rect 198832 9392 198884 9444
rect 380716 9392 380768 9444
rect 448980 9392 449032 9444
rect 92112 9324 92164 9376
rect 196072 9324 196124 9376
rect 384856 9324 384908 9376
rect 456064 9324 456116 9376
rect 88524 9256 88576 9308
rect 194784 9256 194836 9308
rect 386236 9256 386288 9308
rect 459652 9256 459704 9308
rect 84936 9188 84988 9240
rect 193312 9188 193364 9240
rect 388996 9188 389048 9240
rect 463240 9188 463292 9240
rect 81440 9120 81492 9172
rect 190552 9120 190604 9172
rect 391756 9120 391808 9172
rect 470324 9120 470376 9172
rect 77852 9052 77904 9104
rect 189172 9052 189224 9104
rect 445576 9052 445628 9104
rect 573824 9052 573876 9104
rect 74264 8984 74316 9036
rect 187792 8984 187844 9036
rect 446956 8984 447008 9036
rect 577412 8984 577464 9036
rect 31484 8916 31536 8968
rect 165712 8916 165764 8968
rect 448336 8916 448388 8968
rect 581000 8916 581052 8968
rect 117136 8848 117188 8900
rect 209872 8848 209924 8900
rect 120632 8780 120684 8832
rect 211344 8780 211396 8832
rect 124220 8712 124272 8764
rect 212632 8712 212684 8764
rect 131396 8644 131448 8696
rect 216772 8644 216824 8696
rect 134892 8576 134944 8628
rect 218244 8576 218296 8628
rect 138480 8508 138532 8560
rect 220912 8508 220964 8560
rect 142068 8440 142120 8492
rect 222384 8440 222436 8492
rect 145656 8372 145708 8424
rect 223672 8372 223724 8424
rect 156328 8304 156380 8356
rect 229284 8304 229336 8356
rect 119436 8236 119488 8288
rect 211160 8236 211212 8288
rect 422116 8236 422168 8288
rect 527456 8236 527508 8288
rect 2780 8168 2832 8220
rect 4804 8168 4856 8220
rect 115940 8168 115992 8220
rect 208584 8168 208636 8220
rect 423404 8168 423456 8220
rect 531044 8168 531096 8220
rect 112352 8100 112404 8152
rect 207204 8100 207256 8152
rect 420828 8100 420880 8152
rect 424876 8100 424928 8152
rect 534540 8100 534592 8152
rect 108764 8032 108816 8084
rect 205640 8032 205692 8084
rect 426256 8032 426308 8084
rect 538128 8032 538180 8084
rect 105176 7964 105228 8016
rect 202972 7964 203024 8016
rect 429108 7964 429160 8016
rect 541716 7964 541768 8016
rect 101588 7896 101640 7948
rect 201684 7896 201736 7948
rect 430396 7896 430448 7948
rect 545304 7896 545356 7948
rect 98092 7828 98144 7880
rect 200212 7828 200264 7880
rect 431684 7828 431736 7880
rect 548892 7828 548944 7880
rect 94504 7760 94556 7812
rect 197452 7760 197504 7812
rect 434536 7760 434588 7812
rect 552388 7760 552440 7812
rect 90916 7692 90968 7744
rect 196348 7692 196400 7744
rect 435916 7692 435968 7744
rect 555976 7692 556028 7744
rect 87328 7624 87380 7676
rect 194600 7624 194652 7676
rect 369676 7624 369728 7676
rect 427544 7624 427596 7676
rect 437296 7624 437348 7676
rect 559564 7624 559616 7676
rect 23112 7556 23164 7608
rect 161572 7556 161624 7608
rect 162308 7556 162360 7608
rect 233424 7556 233476 7608
rect 123024 7488 123076 7540
rect 212724 7488 212776 7540
rect 127808 7420 127860 7472
rect 215392 7420 215444 7472
rect 373724 7420 373776 7472
rect 434536 7556 434588 7608
rect 441436 7556 441488 7608
rect 566740 7556 566792 7608
rect 419356 7488 419408 7540
rect 523868 7488 523920 7540
rect 411076 7420 411128 7472
rect 508412 7420 508464 7472
rect 126612 7352 126664 7404
rect 214104 7352 214156 7404
rect 409788 7352 409840 7404
rect 504824 7352 504876 7404
rect 130200 7284 130252 7336
rect 216680 7284 216732 7336
rect 408316 7284 408368 7336
rect 501236 7284 501288 7336
rect 133788 7216 133840 7268
rect 218152 7216 218204 7268
rect 405556 7216 405608 7268
rect 497740 7216 497792 7268
rect 137284 7148 137336 7200
rect 219532 7148 219584 7200
rect 404268 7148 404320 7200
rect 494152 7148 494204 7200
rect 140872 7080 140924 7132
rect 222292 7080 222344 7132
rect 402796 7080 402848 7132
rect 490564 7080 490616 7132
rect 144460 7012 144512 7064
rect 223580 7012 223632 7064
rect 400036 7012 400088 7064
rect 486976 7012 487028 7064
rect 148048 6944 148100 6996
rect 225144 6944 225196 6996
rect 258172 6944 258224 6996
rect 379244 6944 379296 6996
rect 445392 6944 445444 6996
rect 150808 6876 150860 6928
rect 150900 6876 150952 6928
rect 258080 6876 258132 6928
rect 67180 6808 67232 6860
rect 183744 6808 183796 6860
rect 398748 6808 398800 6860
rect 483480 6808 483532 6860
rect 63592 6740 63644 6792
rect 182272 6740 182324 6792
rect 401508 6740 401560 6792
rect 488172 6740 488224 6792
rect 60004 6672 60056 6724
rect 180892 6672 180944 6724
rect 402888 6672 402940 6724
rect 491760 6672 491812 6724
rect 56416 6604 56468 6656
rect 178224 6604 178276 6656
rect 405648 6604 405700 6656
rect 495348 6604 495400 6656
rect 52828 6536 52880 6588
rect 176752 6536 176804 6588
rect 178960 6536 179012 6588
rect 241612 6536 241664 6588
rect 407028 6536 407080 6588
rect 498936 6536 498988 6588
rect 49332 6468 49384 6520
rect 175280 6468 175332 6520
rect 175372 6468 175424 6520
rect 239036 6468 239088 6520
rect 408408 6468 408460 6520
rect 502432 6468 502484 6520
rect 40960 6400 41012 6452
rect 169852 6400 169904 6452
rect 171784 6400 171836 6452
rect 237564 6400 237616 6452
rect 353116 6400 353168 6452
rect 395344 6400 395396 6452
rect 411168 6400 411220 6452
rect 506020 6400 506072 6452
rect 18328 6332 18380 6384
rect 158904 6332 158956 6384
rect 161112 6332 161164 6384
rect 231860 6332 231912 6384
rect 355876 6332 355928 6384
rect 399024 6332 399076 6384
rect 412548 6332 412600 6384
rect 509608 6332 509660 6384
rect 13636 6264 13688 6316
rect 156144 6264 156196 6316
rect 159916 6264 159968 6316
rect 231952 6264 232004 6316
rect 358636 6264 358688 6316
rect 406108 6264 406160 6316
rect 413836 6264 413888 6316
rect 513196 6264 513248 6316
rect 8852 6196 8904 6248
rect 153384 6196 153436 6248
rect 157524 6196 157576 6248
rect 230572 6196 230624 6248
rect 362684 6196 362736 6248
rect 413284 6196 413336 6248
rect 416504 6196 416556 6248
rect 516784 6196 516836 6248
rect 4068 6128 4120 6180
rect 151912 6128 151964 6180
rect 153936 6128 153988 6180
rect 227812 6128 227864 6180
rect 364156 6128 364208 6180
rect 416872 6128 416924 6180
rect 418068 6128 418120 6180
rect 520280 6128 520332 6180
rect 129004 6060 129056 6112
rect 215300 6060 215352 6112
rect 400128 6060 400180 6112
rect 484584 6060 484636 6112
rect 132592 5992 132644 6044
rect 218060 5992 218112 6044
rect 397368 5992 397420 6044
rect 479892 5992 479944 6044
rect 136088 5924 136140 5976
rect 219440 5924 219492 5976
rect 394608 5924 394660 5976
rect 476304 5924 476356 5976
rect 139676 5856 139728 5908
rect 220820 5856 220872 5908
rect 393228 5856 393280 5908
rect 472716 5856 472768 5908
rect 143264 5788 143316 5840
rect 222200 5788 222252 5840
rect 391848 5788 391900 5840
rect 469128 5788 469180 5840
rect 146852 5720 146904 5772
rect 224960 5720 225012 5772
rect 389088 5720 389140 5772
rect 465632 5720 465684 5772
rect 150440 5652 150492 5704
rect 226524 5652 226576 5704
rect 387708 5652 387760 5704
rect 462044 5652 462096 5704
rect 99288 5584 99340 5636
rect 163504 5584 163556 5636
rect 164700 5584 164752 5636
rect 233332 5584 233384 5636
rect 386328 5584 386380 5636
rect 458456 5584 458508 5636
rect 113548 5516 113600 5568
rect 160744 5516 160796 5568
rect 168196 5516 168248 5568
rect 236092 5516 236144 5568
rect 384948 5516 385000 5568
rect 454868 5516 454920 5568
rect 51632 5448 51684 5500
rect 175464 5448 175516 5500
rect 183468 5448 183520 5500
rect 187240 5448 187292 5500
rect 245660 5448 245712 5500
rect 362776 5448 362828 5500
rect 412088 5448 412140 5500
rect 416596 5448 416648 5500
rect 48136 5380 48188 5432
rect 173992 5380 174044 5432
rect 174176 5380 174228 5432
rect 181536 5380 181588 5432
rect 33876 5312 33928 5364
rect 93860 5312 93912 5364
rect 103428 5312 103480 5364
rect 113180 5312 113232 5364
rect 122656 5312 122708 5364
rect 132500 5312 132552 5364
rect 141976 5312 142028 5364
rect 30288 5244 30340 5296
rect 26700 5176 26752 5228
rect 152740 5312 152792 5364
rect 167092 5312 167144 5364
rect 244372 5380 244424 5432
rect 360016 5380 360068 5432
rect 408500 5380 408552 5432
rect 419448 5448 419500 5500
rect 424140 5380 424192 5432
rect 429936 5380 429988 5432
rect 431776 5380 431828 5432
rect 432604 5448 432656 5500
rect 540520 5448 540572 5500
rect 432788 5380 432840 5432
rect 242992 5312 243044 5364
rect 364248 5312 364300 5364
rect 415676 5312 415728 5364
rect 430488 5312 430540 5364
rect 544108 5380 544160 5432
rect 433248 5312 433300 5364
rect 178684 5244 178736 5296
rect 238852 5244 238904 5296
rect 365628 5244 365680 5296
rect 419172 5244 419224 5296
rect 547696 5312 547748 5364
rect 21916 5108 21968 5160
rect 170588 5176 170640 5228
rect 237380 5176 237432 5228
rect 368388 5176 368440 5228
rect 422760 5176 422812 5228
rect 162860 5108 162912 5160
rect 17316 5040 17368 5092
rect 158812 5040 158864 5092
rect 7656 4972 7708 5024
rect 142160 4972 142212 5024
rect 160192 5040 160244 5092
rect 164332 5108 164384 5160
rect 167184 5108 167236 5160
rect 234804 5108 234856 5160
rect 369768 5108 369820 5160
rect 426348 5176 426400 5228
rect 163504 5040 163556 5092
rect 233240 5040 233292 5092
rect 371056 5040 371108 5092
rect 403624 5040 403676 5092
rect 158996 4972 159048 5024
rect 230480 4972 230532 5024
rect 373816 4972 373868 5024
rect 379336 4972 379388 5024
rect 379520 4972 379572 5024
rect 398748 4972 398800 5024
rect 420092 5040 420144 5092
rect 427636 5108 427688 5160
rect 432604 5108 432656 5160
rect 551192 5244 551244 5296
rect 437388 5176 437440 5228
rect 433524 5108 433576 5160
rect 436008 5108 436060 5160
rect 441528 5108 441580 5160
rect 554780 5176 554832 5228
rect 2872 4904 2924 4956
rect 150808 4904 150860 4956
rect 150900 4904 150952 4956
rect 153200 4904 153252 4956
rect 155224 4904 155276 4956
rect 229100 4904 229152 4956
rect 375288 4904 375340 4956
rect 572 4836 624 4888
rect 149060 4836 149112 4888
rect 149244 4836 149296 4888
rect 226340 4836 226392 4888
rect 237196 4836 237248 4888
rect 270592 4836 270644 4888
rect 379428 4836 379480 4888
rect 398840 4836 398892 4888
rect 1676 4768 1728 4820
rect 150532 4768 150584 4820
rect 151544 4768 151596 4820
rect 227904 4768 227956 4820
rect 233700 4768 233752 4820
rect 269212 4768 269264 4820
rect 376668 4768 376720 4820
rect 55220 4700 55272 4752
rect 178040 4700 178092 4752
rect 188436 4700 188488 4752
rect 245936 4700 245988 4752
rect 358728 4700 358780 4752
rect 404912 4768 404964 4820
rect 405004 4768 405056 4820
rect 432420 4836 432472 4888
rect 432788 5040 432840 5092
rect 558368 5108 558420 5160
rect 565544 5040 565596 5092
rect 432696 4972 432748 5024
rect 437020 4972 437072 5024
rect 438676 4972 438728 5024
rect 561956 4972 562008 5024
rect 440608 4904 440660 4956
rect 569040 4904 569092 4956
rect 427636 4768 427688 4820
rect 431132 4768 431184 4820
rect 438216 4836 438268 4888
rect 444196 4836 444248 4888
rect 444288 4836 444340 4888
rect 572628 4836 572680 4888
rect 422208 4700 422260 4752
rect 441804 4768 441856 4820
rect 442816 4768 442868 4820
rect 447048 4768 447100 4820
rect 576216 4768 576268 4820
rect 58808 4632 58860 4684
rect 179512 4632 179564 4684
rect 184848 4632 184900 4684
rect 194416 4632 194468 4684
rect 249984 4632 250036 4684
rect 354588 4632 354640 4684
rect 397828 4632 397880 4684
rect 398104 4632 398156 4684
rect 398840 4632 398892 4684
rect 65984 4564 66036 4616
rect 183560 4564 183612 4616
rect 192024 4564 192076 4616
rect 248512 4564 248564 4616
rect 353208 4564 353260 4616
rect 394240 4564 394292 4616
rect 394424 4564 394476 4616
rect 403716 4564 403768 4616
rect 536932 4700 536984 4752
rect 424784 4632 424836 4684
rect 533436 4632 533488 4684
rect 529848 4564 529900 4616
rect 62396 4496 62448 4548
rect 180984 4496 181036 4548
rect 190828 4496 190880 4548
rect 247316 4496 247368 4548
rect 357164 4496 357216 4548
rect 401324 4496 401376 4548
rect 401416 4496 401468 4548
rect 403440 4496 403492 4548
rect 426348 4496 426400 4548
rect 526260 4496 526312 4548
rect 69480 4428 69532 4480
rect 185216 4428 185268 4480
rect 195612 4428 195664 4480
rect 249892 4428 249944 4480
rect 351828 4428 351880 4480
rect 391848 4428 391900 4480
rect 73068 4360 73120 4412
rect 186412 4360 186464 4412
rect 76656 4292 76708 4344
rect 189080 4292 189132 4344
rect 198096 4360 198148 4412
rect 251272 4360 251324 4412
rect 351736 4360 351788 4412
rect 390652 4360 390704 4412
rect 391388 4360 391440 4412
rect 394700 4428 394752 4480
rect 423956 4428 424008 4480
rect 519084 4428 519136 4480
rect 200764 4292 200816 4344
rect 201500 4292 201552 4344
rect 252836 4292 252888 4344
rect 350448 4292 350500 4344
rect 388260 4292 388312 4344
rect 427912 4360 427964 4412
rect 522672 4360 522724 4412
rect 80244 4224 80296 4276
rect 190460 4224 190512 4276
rect 205088 4224 205140 4276
rect 255412 4224 255464 4276
rect 347688 4224 347740 4276
rect 384672 4224 384724 4276
rect 83832 4156 83884 4208
rect 191840 4156 191892 4208
rect 212264 4156 212316 4208
rect 258080 4156 258132 4208
rect 346216 4156 346268 4208
rect 381176 4156 381228 4208
rect 382188 4156 382240 4208
rect 39764 4088 39816 4140
rect 42064 4088 42116 4140
rect 61200 4088 61252 4140
rect 175924 4088 175976 4140
rect 196808 4088 196860 4140
rect 197268 4088 197320 4140
rect 199200 4088 199252 4140
rect 203524 4088 203576 4140
rect 207480 4088 207532 4140
rect 208308 4088 208360 4140
rect 211068 4088 211120 4140
rect 211804 4088 211856 4140
rect 214656 4088 214708 4140
rect 215208 4088 215260 4140
rect 222936 4088 222988 4140
rect 263692 4088 263744 4140
rect 265808 4088 265860 4140
rect 266268 4088 266320 4140
rect 268108 4088 268160 4140
rect 269028 4088 269080 4140
rect 269304 4088 269356 4140
rect 270408 4088 270460 4140
rect 274088 4088 274140 4140
rect 274548 4088 274600 4140
rect 291936 4088 291988 4140
rect 292488 4088 292540 4140
rect 295524 4088 295576 4140
rect 298744 4088 298796 4140
rect 303804 4088 303856 4140
rect 304908 4088 304960 4140
rect 305000 4088 305052 4140
rect 306196 4088 306248 4140
rect 308036 4088 308088 4140
rect 308588 4088 308640 4140
rect 310428 4088 310480 4140
rect 310980 4088 311032 4140
rect 324136 4088 324188 4140
rect 337108 4088 337160 4140
rect 338856 4088 338908 4140
rect 54024 4020 54076 4072
rect 174544 4020 174596 4072
rect 189632 4020 189684 4072
rect 198188 4020 198240 4072
rect 220544 4020 220596 4072
rect 261484 4020 261536 4072
rect 14832 3952 14884 4004
rect 17224 3952 17276 4004
rect 43352 3952 43404 4004
rect 171140 3952 171192 4004
rect 186044 3952 186096 4004
rect 199384 3952 199436 4004
rect 202696 3952 202748 4004
rect 24308 3884 24360 3936
rect 28264 3884 28316 3936
rect 42156 3884 42208 3936
rect 171232 3884 171284 3936
rect 177764 3884 177816 3936
rect 36176 3816 36228 3868
rect 168380 3816 168432 3868
rect 180156 3816 180208 3868
rect 182548 3884 182600 3936
rect 202144 3884 202196 3936
rect 219348 3952 219400 4004
rect 262404 3952 262456 4004
rect 211896 3884 211948 3936
rect 215852 3884 215904 3936
rect 261024 3884 261076 3936
rect 268292 4020 268344 4072
rect 276020 4020 276072 4072
rect 302608 4020 302660 4072
rect 304264 4020 304316 4072
rect 321468 4020 321520 4072
rect 332416 4020 332468 4072
rect 333244 4020 333296 4072
rect 342904 4088 342956 4140
rect 344284 4088 344336 4140
rect 345664 4088 345716 4140
rect 360936 4088 360988 4140
rect 376024 4088 376076 4140
rect 377588 4088 377640 4140
rect 384856 4156 384908 4208
rect 388628 4224 388680 4276
rect 409696 4292 409748 4344
rect 415308 4292 415360 4344
rect 515588 4292 515640 4344
rect 402520 4224 402572 4276
rect 413928 4224 413980 4276
rect 512000 4224 512052 4276
rect 451280 4156 451332 4208
rect 385684 4088 385736 4140
rect 387064 4088 387116 4140
rect 395436 4088 395488 4140
rect 475108 4088 475160 4140
rect 507124 4088 507176 4140
rect 514392 4088 514444 4140
rect 525064 4088 525116 4140
rect 557172 4088 557224 4140
rect 349068 4020 349120 4072
rect 385868 4020 385920 4072
rect 395252 4020 395304 4072
rect 410892 4020 410944 4072
rect 423220 4020 423272 4072
rect 510804 4020 510856 4072
rect 511264 4020 511316 4072
rect 521476 4020 521528 4072
rect 527824 4020 527876 4072
rect 564348 4020 564400 4072
rect 264612 3952 264664 4004
rect 285772 3952 285824 4004
rect 328368 3952 328420 4004
rect 345480 3952 345532 4004
rect 355968 3952 356020 4004
rect 400220 3952 400272 4004
rect 416688 3952 416740 4004
rect 517888 3952 517940 4004
rect 529204 3952 529256 4004
rect 571432 3952 571484 4004
rect 25504 3748 25556 3800
rect 31024 3748 31076 3800
rect 34980 3748 35032 3800
rect 167000 3748 167052 3800
rect 176568 3748 176620 3800
rect 16028 3680 16080 3732
rect 24124 3680 24176 3732
rect 29092 3680 29144 3732
rect 164240 3680 164292 3732
rect 20720 3612 20772 3664
rect 160100 3612 160152 3664
rect 172980 3612 173032 3664
rect 204904 3816 204956 3868
rect 208676 3816 208728 3868
rect 256792 3816 256844 3868
rect 263416 3884 263468 3936
rect 284484 3884 284536 3936
rect 328276 3884 328328 3936
rect 346676 3884 346728 3936
rect 360108 3884 360160 3936
rect 407304 3884 407356 3936
rect 409144 3884 409196 3936
rect 417976 3884 418028 3936
rect 421656 3884 421708 3936
rect 525064 3884 525116 3936
rect 530584 3884 530636 3936
rect 578608 3884 578660 3936
rect 225328 3612 225380 3664
rect 226248 3612 226300 3664
rect 6460 3544 6512 3596
rect 13084 3544 13136 3596
rect 19524 3544 19576 3596
rect 158720 3544 158772 3596
rect 228916 3612 228968 3664
rect 231216 3612 231268 3664
rect 231308 3612 231360 3664
rect 231768 3612 231820 3664
rect 238760 3680 238812 3732
rect 240232 3748 240284 3800
rect 240784 3748 240836 3800
rect 241428 3748 241480 3800
rect 243176 3748 243228 3800
rect 244188 3748 244240 3800
rect 249156 3748 249208 3800
rect 249708 3748 249760 3800
rect 250352 3748 250404 3800
rect 251088 3748 251140 3800
rect 251456 3748 251508 3800
rect 252468 3748 252520 3800
rect 261024 3748 261076 3800
rect 283012 3816 283064 3868
rect 319996 3816 320048 3868
rect 330024 3816 330076 3868
rect 331128 3816 331180 3868
rect 352564 3816 352616 3868
rect 362868 3816 362920 3868
rect 414480 3816 414532 3868
rect 423588 3816 423640 3868
rect 532240 3816 532292 3868
rect 320088 3748 320140 3800
rect 331220 3748 331272 3800
rect 333888 3748 333940 3800
rect 356152 3748 356204 3800
rect 356704 3748 356756 3800
rect 364524 3748 364576 3800
rect 367008 3748 367060 3800
rect 420368 3748 420420 3800
rect 427728 3748 427780 3800
rect 539324 3748 539376 3800
rect 244464 3680 244516 3732
rect 236000 3612 236052 3664
rect 243544 3612 243596 3664
rect 250444 3680 250496 3732
rect 252652 3680 252704 3732
rect 278872 3680 278924 3732
rect 285956 3680 286008 3732
rect 294604 3680 294656 3732
rect 321376 3680 321428 3732
rect 333612 3680 333664 3732
rect 335268 3680 335320 3732
rect 359740 3680 359792 3732
rect 366916 3680 366968 3732
rect 421564 3680 421616 3732
rect 431868 3680 431920 3732
rect 546500 3680 546552 3732
rect 246764 3612 246816 3664
rect 273260 3612 273312 3664
rect 282460 3612 282512 3664
rect 294144 3612 294196 3664
rect 300308 3612 300360 3664
rect 303620 3612 303672 3664
rect 316776 3612 316828 3664
rect 320456 3612 320508 3664
rect 322756 3612 322808 3664
rect 335912 3612 335964 3664
rect 339408 3612 339460 3664
rect 11244 3476 11296 3528
rect 154856 3476 154908 3528
rect 169392 3476 169444 3528
rect 236276 3544 236328 3596
rect 241520 3544 241572 3596
rect 241980 3544 242032 3596
rect 277676 3544 277728 3596
rect 286324 3544 286376 3596
rect 316684 3544 316736 3596
rect 318064 3544 318116 3596
rect 324228 3544 324280 3596
rect 338304 3544 338356 3596
rect 340788 3544 340840 3596
rect 363328 3612 363380 3664
rect 371148 3612 371200 3664
rect 428740 3612 428792 3664
rect 434628 3612 434680 3664
rect 553584 3612 553636 3664
rect 366916 3544 366968 3596
rect 372528 3544 372580 3596
rect 432328 3544 432380 3596
rect 438768 3544 438820 3596
rect 560760 3544 560812 3596
rect 239588 3476 239640 3528
rect 271972 3476 272024 3528
rect 301412 3476 301464 3528
rect 302884 3476 302936 3528
rect 312544 3476 312596 3528
rect 313372 3476 313424 3528
rect 322204 3476 322256 3528
rect 325240 3476 325292 3528
rect 325608 3476 325660 3528
rect 339500 3476 339552 3528
rect 370412 3476 370464 3528
rect 373908 3476 373960 3528
rect 435824 3476 435876 3528
rect 442908 3476 442960 3528
rect 567844 3476 567896 3528
rect 10048 3408 10100 3460
rect 154672 3408 154724 3460
rect 165896 3408 165948 3460
rect 234620 3408 234672 3460
rect 234804 3408 234856 3460
rect 268476 3408 268528 3460
rect 270500 3408 270552 3460
rect 32680 3340 32732 3392
rect 35164 3340 35216 3392
rect 68284 3340 68336 3392
rect 177304 3340 177356 3392
rect 183744 3340 183796 3392
rect 200396 3340 200448 3392
rect 201408 3340 201460 3392
rect 38568 3272 38620 3324
rect 71044 3272 71096 3324
rect 75460 3272 75512 3324
rect 180064 3272 180116 3324
rect 45744 3204 45796 3256
rect 75184 3204 75236 3256
rect 82636 3204 82688 3256
rect 181444 3204 181496 3256
rect 209872 3204 209924 3256
rect 244372 3204 244424 3256
rect 253848 3272 253900 3324
rect 254676 3272 254728 3324
rect 257436 3272 257488 3324
rect 257988 3272 258040 3324
rect 258632 3340 258684 3392
rect 259368 3340 259420 3392
rect 261576 3340 261628 3392
rect 262220 3340 262272 3392
rect 263508 3340 263560 3392
rect 276480 3408 276532 3460
rect 277308 3408 277360 3460
rect 278872 3408 278924 3460
rect 284944 3340 284996 3392
rect 289544 3408 289596 3460
rect 297364 3408 297416 3460
rect 297916 3408 297968 3460
rect 301596 3408 301648 3460
rect 311808 3408 311860 3460
rect 314568 3408 314620 3460
rect 315948 3408 316000 3460
rect 322848 3408 322900 3460
rect 326988 3408 327040 3460
rect 343088 3408 343140 3460
rect 344928 3408 344980 3460
rect 378784 3408 378836 3460
rect 291844 3340 291896 3392
rect 294328 3340 294380 3392
rect 297456 3340 297508 3392
rect 322940 3340 322992 3392
rect 334716 3340 334768 3392
rect 340144 3340 340196 3392
rect 259828 3272 259880 3324
rect 280804 3272 280856 3324
rect 284760 3272 284812 3324
rect 290464 3272 290516 3324
rect 323584 3272 323636 3324
rect 328828 3272 328880 3324
rect 330484 3272 330536 3324
rect 340696 3272 340748 3324
rect 349068 3340 349120 3392
rect 350264 3272 350316 3324
rect 254584 3204 254636 3256
rect 320824 3204 320876 3256
rect 324044 3204 324096 3256
rect 50528 3136 50580 3188
rect 77944 3136 77996 3188
rect 89720 3136 89772 3188
rect 93124 3136 93176 3188
rect 57612 3068 57664 3120
rect 84844 3068 84896 3120
rect 86132 3068 86184 3120
rect 184204 3136 184256 3188
rect 217048 3136 217100 3188
rect 224132 3136 224184 3188
rect 262864 3136 262916 3188
rect 299112 3136 299164 3188
rect 301504 3136 301556 3188
rect 341524 3136 341576 3188
rect 353760 3340 353812 3392
rect 359464 3340 359516 3392
rect 371608 3340 371660 3392
rect 358084 3272 358136 3324
rect 368020 3272 368072 3324
rect 380164 3272 380216 3324
rect 389456 3272 389508 3324
rect 380256 3204 380308 3256
rect 443000 3408 443052 3460
rect 445668 3408 445720 3460
rect 575020 3408 575072 3460
rect 391204 3340 391256 3392
rect 403716 3340 403768 3392
rect 403808 3340 403860 3392
rect 482284 3340 482336 3392
rect 523684 3340 523736 3392
rect 550088 3340 550140 3392
rect 392584 3272 392636 3324
rect 424324 3272 424376 3324
rect 503628 3272 503680 3324
rect 520924 3272 520976 3324
rect 542912 3272 542964 3324
rect 467932 3204 467984 3256
rect 518164 3204 518216 3256
rect 535736 3204 535788 3256
rect 384304 3136 384356 3188
rect 393044 3136 393096 3188
rect 93308 3068 93360 3120
rect 185584 3068 185636 3120
rect 221740 3068 221792 3120
rect 266452 3068 266504 3120
rect 267004 3068 267056 3120
rect 267648 3068 267700 3120
rect 377404 3068 377456 3120
rect 382372 3068 382424 3120
rect 388536 3068 388588 3120
rect 460848 3136 460900 3188
rect 514024 3136 514076 3188
rect 528652 3136 528704 3188
rect 46940 3000 46992 3052
rect 95884 3000 95936 3052
rect 96896 3000 96948 3052
rect 98644 3000 98696 3052
rect 103980 3000 104032 3052
rect 104808 3000 104860 3052
rect 111156 3000 111208 3052
rect 111708 3000 111760 3052
rect 71872 2932 71924 2984
rect 86224 2932 86276 2984
rect 100484 2932 100536 2984
rect 186964 3000 187016 3052
rect 193220 3000 193272 3052
rect 198004 3000 198056 3052
rect 206284 3000 206336 3052
rect 226984 3000 227036 3052
rect 230112 3000 230164 3052
rect 267832 3000 267884 3052
rect 275284 3000 275336 3052
rect 275928 3000 275980 3052
rect 287152 3000 287204 3052
rect 288256 3000 288308 3052
rect 293132 3000 293184 3052
rect 298836 3000 298888 3052
rect 338764 3000 338816 3052
rect 341892 3000 341944 3052
rect 388444 3000 388496 3052
rect 396632 3000 396684 3052
rect 64788 2864 64840 2916
rect 106924 2864 106976 2916
rect 79048 2796 79100 2848
rect 88984 2796 89036 2848
rect 107568 2796 107620 2848
rect 188620 2932 188672 2984
rect 226524 2932 226576 2984
rect 264980 2932 265032 2984
rect 283656 2932 283708 2984
rect 284208 2932 284260 2984
rect 384396 2932 384448 2984
rect 114744 2864 114796 2916
rect 115848 2864 115900 2916
rect 121828 2864 121880 2916
rect 122748 2864 122800 2916
rect 125416 2864 125468 2916
rect 118240 2796 118292 2848
rect 188344 2864 188396 2916
rect 227720 2864 227772 2916
rect 232504 2864 232556 2916
rect 269212 2864 269264 2916
rect 296720 2864 296772 2916
rect 302424 2864 302476 2916
rect 450176 3068 450228 3120
rect 411904 3000 411956 3052
rect 425152 3000 425204 3052
rect 435364 3000 435416 3052
rect 496544 3000 496596 3052
rect 502984 3000 503036 3052
rect 507216 3000 507268 3052
rect 421472 2932 421524 2984
rect 481088 2932 481140 2984
rect 420184 2864 420236 2916
rect 477500 2864 477552 2916
rect 191104 2796 191156 2848
rect 218152 2796 218204 2848
rect 257344 2796 257396 2848
rect 291108 2796 291160 2848
rect 431224 2796 431276 2848
rect 489368 2796 489420 2848
rect 374276 2660 374328 2712
rect 374092 1504 374144 1556
rect 375196 1504 375248 1556
rect 238392 552 238444 604
rect 238576 552 238628 604
rect 256240 552 256292 604
rect 256608 552 256660 604
rect 281264 552 281316 604
rect 281448 552 281500 604
rect 290740 595 290792 604
rect 290740 561 290749 595
rect 290749 561 290783 595
rect 290783 561 290792 595
rect 290740 552 290792 561
rect 325792 552 325844 604
rect 326436 552 326488 604
rect 350816 552 350868 604
rect 351368 552 351420 604
rect 361856 552 361908 604
rect 362132 552 362184 604
rect 368480 552 368532 604
rect 369216 552 369268 604
rect 372620 552 372672 604
rect 372804 552 372856 604
rect 374000 595 374052 604
rect 374000 561 374009 595
rect 374009 561 374043 595
rect 374043 561 374052 595
rect 374000 552 374052 561
rect 379704 552 379756 604
rect 379980 552 380032 604
rect 382464 552 382516 604
rect 383568 552 383620 604
rect 439044 552 439096 604
rect 439412 552 439464 604
rect 445760 552 445812 604
rect 446588 552 446640 604
rect 470600 552 470652 604
rect 471520 552 471572 604
rect 473360 552 473412 604
rect 473912 552 473964 604
rect 477592 552 477644 604
rect 478696 552 478748 604
rect 499580 552 499632 604
rect 500132 552 500184 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700602 73016 703520
rect 89180 700670 89208 703520
rect 105464 700738 105492 703520
rect 137848 700942 137876 703520
rect 154132 701010 154160 703520
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 105452 700732 105504 700738
rect 105452 700674 105504 700680
rect 89168 700664 89220 700670
rect 89168 700606 89220 700612
rect 72976 700596 73028 700602
rect 72976 700538 73028 700544
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 170324 700262 170352 703520
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 202800 700058 202828 703520
rect 202788 700052 202840 700058
rect 202788 699994 202840 700000
rect 218992 699990 219020 703520
rect 218980 699984 219032 699990
rect 218980 699926 219032 699932
rect 235184 699718 235212 703520
rect 267660 699786 267688 703520
rect 278688 700868 278740 700874
rect 278688 700810 278740 700816
rect 270408 700528 270460 700534
rect 270408 700470 270460 700476
rect 267648 699780 267700 699786
rect 267648 699722 267700 699728
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 567254 3464 567287
rect 3424 567248 3476 567254
rect 3424 567190 3476 567196
rect 3422 553072 3478 553081
rect 3422 553007 3478 553016
rect 3436 552158 3464 553007
rect 3424 552152 3476 552158
rect 3424 552094 3476 552100
rect 156420 552084 156472 552090
rect 156420 552026 156472 552032
rect 4802 549264 4858 549273
rect 4802 549199 4858 549208
rect 2964 549024 3016 549030
rect 2964 548966 3016 548972
rect 2976 538665 3004 548966
rect 4712 548956 4764 548962
rect 4712 548898 4764 548904
rect 3056 548820 3108 548826
rect 3056 548762 3108 548768
rect 2962 538656 3018 538665
rect 2962 538591 3018 538600
rect 2964 509992 3016 509998
rect 2962 509960 2964 509969
rect 3016 509960 3018 509969
rect 2962 509895 3018 509904
rect 2780 495576 2832 495582
rect 2778 495544 2780 495553
rect 2832 495544 2834 495553
rect 2778 495479 2834 495488
rect 2780 481160 2832 481166
rect 2778 481128 2780 481137
rect 2832 481128 2834 481137
rect 2778 481063 2834 481072
rect 3068 452441 3096 548762
rect 3148 548684 3200 548690
rect 3148 548626 3200 548632
rect 3054 452432 3110 452441
rect 3054 452367 3110 452376
rect 2780 438592 2832 438598
rect 2780 438534 2832 438540
rect 2792 438025 2820 438534
rect 2778 438016 2834 438025
rect 2778 437951 2834 437960
rect 2780 424856 2832 424862
rect 2780 424798 2832 424804
rect 2792 423745 2820 424798
rect 2778 423736 2834 423745
rect 2778 423671 2834 423680
rect 3160 395049 3188 548626
rect 3240 548480 3292 548486
rect 3240 548422 3292 548428
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 2964 380656 3016 380662
rect 2962 380624 2964 380633
rect 3016 380624 3018 380633
rect 2962 380559 3018 380568
rect 2780 366988 2832 366994
rect 2780 366930 2832 366936
rect 2792 366217 2820 366930
rect 2778 366208 2834 366217
rect 2778 366143 2834 366152
rect 3252 337521 3280 548422
rect 4068 548344 4120 548350
rect 4068 548286 4120 548292
rect 3976 548072 4028 548078
rect 3698 548040 3754 548049
rect 3976 548014 4028 548020
rect 3698 547975 3754 547984
rect 3608 543856 3660 543862
rect 3608 543798 3660 543804
rect 3424 543788 3476 543794
rect 3424 543730 3476 543736
rect 3330 543008 3386 543017
rect 3330 542943 3386 542952
rect 3238 337512 3294 337521
rect 3238 337447 3294 337456
rect 3148 324148 3200 324154
rect 3148 324090 3200 324096
rect 3160 323105 3188 324090
rect 3146 323096 3202 323105
rect 3146 323031 3202 323040
rect 3344 308825 3372 542943
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3148 280152 3200 280158
rect 3146 280120 3148 280129
rect 3200 280120 3202 280129
rect 3146 280055 3202 280064
rect 2780 266212 2832 266218
rect 2780 266154 2832 266160
rect 2792 265713 2820 266154
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 3056 237380 3108 237386
rect 3056 237322 3108 237328
rect 3068 237017 3096 237322
rect 3054 237008 3110 237017
rect 3054 236943 3110 236952
rect 3332 223576 3384 223582
rect 3332 223518 3384 223524
rect 3344 222601 3372 223518
rect 3330 222592 3386 222601
rect 3330 222527 3386 222536
rect 2780 193928 2832 193934
rect 2778 193896 2780 193905
rect 2832 193896 2834 193905
rect 2778 193831 2834 193840
rect 2780 179512 2832 179518
rect 2778 179480 2780 179489
rect 2832 179480 2834 179489
rect 2778 179415 2834 179424
rect 3332 151768 3384 151774
rect 3332 151710 3384 151716
rect 3344 150793 3372 151710
rect 3330 150784 3386 150793
rect 3330 150719 3386 150728
rect 2962 122768 3018 122777
rect 2962 122703 3018 122712
rect 2976 122097 3004 122703
rect 2962 122088 3018 122097
rect 2962 122023 3018 122032
rect 3330 80064 3386 80073
rect 3330 79999 3386 80008
rect 3344 78985 3372 79999
rect 3330 78976 3386 78985
rect 3330 78911 3386 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3436 21457 3464 543730
rect 3516 542836 3568 542842
rect 3516 542778 3568 542784
rect 3528 35873 3556 542778
rect 3620 50153 3648 543798
rect 3712 93265 3740 547975
rect 3884 544060 3936 544066
rect 3884 544002 3936 544008
rect 3792 543924 3844 543930
rect 3792 543866 3844 543872
rect 3804 107681 3832 543866
rect 3896 136377 3924 544002
rect 3988 251297 4016 548014
rect 4080 294409 4108 548286
rect 4724 495582 4752 548898
rect 4712 495576 4764 495582
rect 4712 495518 4764 495524
rect 4066 294400 4122 294409
rect 4066 294335 4122 294344
rect 3974 251288 4030 251297
rect 3974 251223 4030 251232
rect 3882 136368 3938 136377
rect 3882 136303 3938 136312
rect 3790 107672 3846 107681
rect 3790 107607 3846 107616
rect 3698 93256 3754 93265
rect 3698 93191 3754 93200
rect 3606 50144 3662 50153
rect 3606 50079 3662 50088
rect 3514 35864 3570 35873
rect 3514 35799 3570 35808
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 4816 8226 4844 549199
rect 5264 548888 5316 548894
rect 5264 548830 5316 548836
rect 5172 548616 5224 548622
rect 5172 548558 5224 548564
rect 5080 548276 5132 548282
rect 5080 548218 5132 548224
rect 4896 547936 4948 547942
rect 4896 547878 4948 547884
rect 4908 179518 4936 547878
rect 4988 544264 5040 544270
rect 4988 544206 5040 544212
rect 5000 193934 5028 544206
rect 5092 266218 5120 548218
rect 5184 366994 5212 548558
rect 5276 424862 5304 548830
rect 5356 548752 5408 548758
rect 5356 548694 5408 548700
rect 5368 438598 5396 548694
rect 6368 548548 6420 548554
rect 6368 548490 6420 548496
rect 6276 548412 6328 548418
rect 6276 548354 6328 548360
rect 6184 548208 6236 548214
rect 6184 548150 6236 548156
rect 5448 545284 5500 545290
rect 5448 545226 5500 545232
rect 5460 481166 5488 545226
rect 5448 481160 5500 481166
rect 5448 481102 5500 481108
rect 5356 438592 5408 438598
rect 5356 438534 5408 438540
rect 5264 424856 5316 424862
rect 5264 424798 5316 424804
rect 5172 366988 5224 366994
rect 5172 366930 5224 366936
rect 6196 280158 6224 548150
rect 6288 324154 6316 548354
rect 6380 380662 6408 548490
rect 21362 548312 21418 548321
rect 21362 548247 21418 548256
rect 10324 548140 10376 548146
rect 10324 548082 10376 548088
rect 6460 544672 6512 544678
rect 6460 544614 6512 544620
rect 6472 509998 6500 544614
rect 6460 509992 6512 509998
rect 6460 509934 6512 509940
rect 6368 380656 6420 380662
rect 6368 380598 6420 380604
rect 6276 324148 6328 324154
rect 6276 324090 6328 324096
rect 6184 280152 6236 280158
rect 6184 280094 6236 280100
rect 5080 266212 5132 266218
rect 5080 266154 5132 266160
rect 10336 237386 10364 548082
rect 19984 548004 20036 548010
rect 19984 547946 20036 547952
rect 17224 242208 17276 242214
rect 13082 242176 13138 242185
rect 17224 242150 17276 242156
rect 13082 242111 13138 242120
rect 10324 237380 10376 237386
rect 10324 237322 10376 237328
rect 4988 193928 5040 193934
rect 4988 193870 5040 193876
rect 4896 179512 4948 179518
rect 4896 179454 4948 179460
rect 2780 8220 2832 8226
rect 2780 8162 2832 8168
rect 4804 8220 4856 8226
rect 4804 8162 4856 8168
rect 2792 7177 2820 8162
rect 2778 7168 2834 7177
rect 2778 7103 2834 7112
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 572 4888 624 4894
rect 572 4830 624 4836
rect 584 480 612 4830
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1688 480 1716 4762
rect 2884 480 2912 4898
rect 4080 480 4108 6122
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 6472 480 6500 3538
rect 7668 480 7696 4966
rect 8864 480 8892 6190
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10060 480 10088 3402
rect 11256 480 11284 3470
rect 12452 480 12480 4791
rect 13096 3602 13124 242111
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13648 480 13676 6258
rect 17236 4010 17264 242150
rect 19996 151774 20024 547946
rect 19984 151768 20036 151774
rect 19984 151710 20036 151716
rect 21376 64870 21404 548247
rect 156432 546244 156460 552026
rect 235920 550186 235948 699654
rect 263508 696992 263560 696998
rect 263508 696934 263560 696940
rect 260748 673532 260800 673538
rect 260748 673474 260800 673480
rect 255228 650072 255280 650078
rect 255228 650014 255280 650020
rect 252468 626612 252520 626618
rect 252468 626554 252520 626560
rect 246948 603152 247000 603158
rect 246948 603094 247000 603100
rect 245568 579692 245620 579698
rect 245568 579634 245620 579640
rect 240048 556232 240100 556238
rect 240048 556174 240100 556180
rect 235908 550180 235960 550186
rect 235908 550122 235960 550128
rect 226248 549228 226300 549234
rect 226248 549170 226300 549176
rect 223672 549160 223724 549166
rect 210698 549128 210754 549137
rect 223672 549102 223724 549108
rect 210698 549063 210754 549072
rect 218428 549092 218480 549098
rect 197818 548992 197874 549001
rect 197818 548927 197874 548936
rect 189998 548720 190054 548729
rect 189998 548655 190054 548664
rect 166722 548448 166778 548457
rect 166722 548383 166778 548392
rect 158994 548176 159050 548185
rect 158994 548111 159050 548120
rect 159008 546244 159036 548111
rect 166736 546244 166764 548383
rect 190012 546244 190040 548655
rect 197832 546244 197860 548927
rect 210712 546244 210740 549063
rect 218428 549034 218480 549040
rect 218440 546244 218468 549034
rect 223684 546244 223712 549102
rect 226260 546244 226288 549170
rect 240060 546394 240088 556174
rect 245580 546394 245608 579634
rect 239784 546366 240088 546394
rect 244936 546366 245608 546394
rect 239784 546258 239812 546366
rect 244936 546258 244964 546366
rect 239154 546230 239812 546258
rect 244398 546230 244964 546258
rect 246960 546244 246988 603094
rect 249708 592068 249760 592074
rect 249708 592010 249760 592016
rect 249720 546258 249748 592010
rect 252480 546258 252508 626554
rect 255240 546394 255268 650014
rect 257988 638988 258040 638994
rect 257988 638930 258040 638936
rect 258000 546394 258028 638930
rect 260760 546394 260788 673474
rect 263520 546394 263548 696934
rect 266268 685908 266320 685914
rect 266268 685850 266320 685856
rect 266280 546394 266308 685850
rect 267648 549908 267700 549914
rect 267648 549850 267700 549856
rect 255056 546366 255268 546394
rect 257632 546366 258028 546394
rect 260300 546366 260788 546394
rect 262876 546366 263548 546394
rect 265452 546366 266308 546394
rect 255056 546258 255084 546366
rect 257632 546258 257660 546366
rect 249550 546230 249748 546258
rect 252126 546230 252508 546258
rect 254702 546230 255084 546258
rect 257278 546230 257660 546258
rect 260300 546122 260328 546366
rect 262876 546122 262904 546366
rect 265452 546122 265480 546366
rect 267660 546244 267688 549850
rect 270420 546258 270448 700470
rect 273168 700460 273220 700466
rect 273168 700402 273220 700408
rect 273180 546258 273208 700402
rect 275376 549976 275428 549982
rect 275376 549918 275428 549924
rect 270250 546230 270448 546258
rect 272826 546230 273208 546258
rect 275388 546244 275416 549918
rect 278700 546122 278728 700810
rect 281448 700800 281500 700806
rect 281448 700742 281500 700748
rect 281460 546394 281488 700742
rect 283852 699718 283880 703520
rect 288348 700188 288400 700194
rect 288348 700130 288400 700136
rect 286968 700120 287020 700126
rect 286968 700062 287020 700068
rect 283840 699712 283892 699718
rect 283840 699654 283892 699660
rect 283104 550044 283156 550050
rect 283104 549986 283156 549992
rect 281184 546366 281488 546394
rect 281184 546258 281212 546366
rect 280554 546230 281212 546258
rect 283116 546244 283144 549986
rect 286980 546394 287008 700062
rect 286336 546366 287008 546394
rect 286336 546258 286364 546366
rect 288360 546258 288388 700130
rect 296628 699916 296680 699922
rect 296628 699858 296680 699864
rect 293868 699848 293920 699854
rect 293868 699790 293920 699796
rect 290924 550112 290976 550118
rect 290924 550054 290976 550060
rect 285706 546230 286364 546258
rect 288282 546230 288388 546258
rect 290936 546244 290964 550054
rect 293880 546258 293908 699790
rect 293526 546230 293908 546258
rect 296640 546122 296668 699858
rect 300136 688634 300164 703520
rect 318800 701004 318852 701010
rect 318800 700946 318852 700952
rect 316040 700936 316092 700942
rect 316040 700878 316092 700884
rect 313280 700256 313332 700262
rect 313280 700198 313332 700204
rect 307760 700052 307812 700058
rect 307760 699994 307812 700000
rect 300860 699780 300912 699786
rect 300860 699722 300912 699728
rect 299664 688628 299716 688634
rect 299664 688570 299716 688576
rect 300124 688628 300176 688634
rect 300124 688570 300176 688576
rect 299676 685930 299704 688570
rect 299584 685902 299704 685930
rect 299584 684486 299612 685902
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 299940 666596 299992 666602
rect 299940 666538 299992 666544
rect 299952 659682 299980 666538
rect 299768 659654 299980 659682
rect 299768 647290 299796 659654
rect 299664 647284 299716 647290
rect 299664 647226 299716 647232
rect 299756 647284 299808 647290
rect 299756 647226 299808 647232
rect 299676 640422 299704 647226
rect 299664 640416 299716 640422
rect 299664 640358 299716 640364
rect 299756 640416 299808 640422
rect 299756 640358 299808 640364
rect 299768 630698 299796 640358
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299756 630692 299808 630698
rect 299756 630634 299808 630640
rect 299584 630578 299612 630634
rect 299584 630550 299704 630578
rect 299676 621058 299704 630550
rect 299676 621030 299796 621058
rect 299768 611386 299796 621030
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 299584 611266 299612 611322
rect 299584 611238 299704 611266
rect 299676 608598 299704 611238
rect 299664 608592 299716 608598
rect 299664 608534 299716 608540
rect 299848 601724 299900 601730
rect 299848 601666 299900 601672
rect 299860 598942 299888 601666
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 299940 589348 299992 589354
rect 299940 589290 299992 589296
rect 299952 582486 299980 589290
rect 299940 582480 299992 582486
rect 299940 582422 299992 582428
rect 299848 582344 299900 582350
rect 299848 582286 299900 582292
rect 299860 572642 299888 582286
rect 299676 572614 299888 572642
rect 299676 569922 299704 572614
rect 299584 569894 299704 569922
rect 299584 563174 299612 569894
rect 299572 563168 299624 563174
rect 299572 563110 299624 563116
rect 299572 563032 299624 563038
rect 299572 562974 299624 562980
rect 299584 560561 299612 562974
rect 299570 560552 299626 560561
rect 299570 560487 299626 560496
rect 299570 560416 299626 560425
rect 299570 560351 299626 560360
rect 299584 560250 299612 560351
rect 299572 560244 299624 560250
rect 299572 560186 299624 560192
rect 299676 550662 299704 550693
rect 299664 550656 299716 550662
rect 299584 550604 299664 550610
rect 299584 550598 299716 550604
rect 299584 550582 299704 550598
rect 299584 549302 299612 550582
rect 298652 549296 298704 549302
rect 298652 549238 298704 549244
rect 299572 549296 299624 549302
rect 299572 549238 299624 549244
rect 298664 546244 298692 549238
rect 300872 546258 300900 699722
rect 303620 699712 303672 699718
rect 303620 699654 303672 699660
rect 303632 546258 303660 699654
rect 306380 550180 306432 550186
rect 306380 550122 306432 550128
rect 300872 546230 301254 546258
rect 303632 546230 303830 546258
rect 306392 546244 306420 550122
rect 307772 546394 307800 699994
rect 310520 699984 310572 699990
rect 310520 699926 310572 699932
rect 310532 546394 310560 699926
rect 313292 546394 313320 700198
rect 316052 546394 316080 700878
rect 307772 546366 308536 546394
rect 310532 546366 311112 546394
rect 313292 546366 313872 546394
rect 316052 546366 316264 546394
rect 308508 546258 308536 546366
rect 311084 546258 311112 546366
rect 313844 546258 313872 546366
rect 316236 546258 316264 546366
rect 318812 546258 318840 700946
rect 321560 700732 321612 700738
rect 321560 700674 321612 700680
rect 321572 546258 321600 700674
rect 327080 700664 327132 700670
rect 327080 700606 327132 700612
rect 324320 700596 324372 700602
rect 324320 700538 324372 700544
rect 324332 546258 324360 700538
rect 308508 546230 308982 546258
rect 311084 546230 311558 546258
rect 313844 546230 314226 546258
rect 316236 546230 316802 546258
rect 318812 546230 319378 546258
rect 321572 546230 321954 546258
rect 324332 546230 324530 546258
rect 327092 546244 327120 700606
rect 328460 700392 328512 700398
rect 328460 700334 328512 700340
rect 331310 700360 331366 700369
rect 328472 546394 328500 700334
rect 331310 700295 331366 700304
rect 331324 546394 331352 700295
rect 332520 699854 332548 703520
rect 333980 700324 334032 700330
rect 333980 700266 334032 700272
rect 332508 699848 332560 699854
rect 332508 699790 332560 699796
rect 333992 546394 334020 700266
rect 348804 699922 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365116 703474
rect 348792 699916 348844 699922
rect 348792 699858 348844 699864
rect 365088 686089 365116 703446
rect 397472 700126 397500 703520
rect 413664 700194 413692 703520
rect 413652 700188 413704 700194
rect 413652 700130 413704 700136
rect 397460 700120 397512 700126
rect 397460 700062 397512 700068
rect 429856 688634 429884 703520
rect 462332 700874 462360 703520
rect 462320 700868 462372 700874
rect 462320 700810 462372 700816
rect 478524 700806 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 365074 686080 365130 686089
rect 365074 686015 365130 686024
rect 364522 685944 364578 685953
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700534 527220 703520
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 543476 700466 543504 703520
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 364522 685879 364578 685888
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 336740 681760 336792 681766
rect 336740 681702 336792 681708
rect 328472 546366 329328 546394
rect 331324 546366 331904 546394
rect 333992 546366 334480 546394
rect 329300 546258 329328 546366
rect 331876 546258 331904 546366
rect 334452 546258 334480 546366
rect 329300 546230 329682 546258
rect 331876 546230 332258 546258
rect 334452 546230 334834 546258
rect 259854 546094 260328 546122
rect 262430 546094 262904 546122
rect 265006 546094 265480 546122
rect 277978 546094 278728 546122
rect 296102 546094 296668 546122
rect 336752 546122 336780 681702
rect 364536 678994 364564 685879
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 364352 678966 364564 678994
rect 494072 678966 494284 678994
rect 364352 676190 364380 678966
rect 494072 676190 494100 678966
rect 364340 676184 364392 676190
rect 364340 676126 364392 676132
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 342260 667956 342312 667962
rect 342260 667898 342312 667904
rect 339500 652792 339552 652798
rect 339500 652734 339552 652740
rect 339512 546394 339540 652734
rect 339512 546366 339632 546394
rect 339604 546258 339632 546366
rect 342272 546258 342300 667898
rect 364432 666596 364484 666602
rect 364432 666538 364484 666544
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 364444 659682 364472 666538
rect 429672 659682 429700 666538
rect 364444 659654 364564 659682
rect 364536 654158 364564 659654
rect 429488 659654 429700 659682
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 364352 644450 364380 654094
rect 429488 647290 429516 659654
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 364352 644422 364564 644450
rect 364536 634846 364564 644422
rect 429396 640422 429424 647226
rect 494072 644450 494100 654094
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 364340 634840 364392 634846
rect 364340 634782 364392 634788
rect 364524 634840 364576 634846
rect 364524 634782 364576 634788
rect 364352 625138 364380 634782
rect 429488 630698 429516 640358
rect 494256 634846 494284 644422
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 364352 625110 364564 625138
rect 345020 623824 345072 623830
rect 345020 623766 345072 623772
rect 345032 546258 345060 623766
rect 364536 615534 364564 625110
rect 429396 621058 429424 630550
rect 494072 625138 494100 634782
rect 559208 630698 559236 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 429396 621030 429516 621058
rect 364340 615528 364392 615534
rect 364340 615470 364392 615476
rect 364524 615528 364576 615534
rect 364524 615470 364576 615476
rect 349160 610020 349212 610026
rect 349160 609962 349212 609968
rect 347780 594856 347832 594862
rect 347780 594798 347832 594804
rect 339604 546230 340078 546258
rect 342272 546230 342654 546258
rect 345032 546230 345230 546258
rect 347792 546244 347820 594798
rect 349172 546394 349200 609962
rect 364352 605826 364380 615470
rect 429488 611386 429516 621030
rect 494256 615534 494284 625110
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 429396 608598 429424 611238
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 494072 605826 494100 615470
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 364352 605798 364564 605826
rect 494072 605798 494284 605826
rect 364536 596222 364564 605798
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 598942 429608 601666
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 494256 596222 494284 605798
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 364340 596216 364392 596222
rect 364524 596216 364576 596222
rect 364392 596164 364472 596170
rect 364340 596158 364472 596164
rect 364524 596158 364576 596164
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 364352 596142 364472 596158
rect 494072 596142 494192 596158
rect 364444 596034 364472 596142
rect 494164 596034 494192 596142
rect 364444 596006 364564 596034
rect 494164 596006 494284 596034
rect 364536 591954 364564 596006
rect 494256 591954 494284 596006
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 364444 591926 364564 591954
rect 494164 591926 494284 591954
rect 364444 589286 364472 591926
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 364156 589280 364208 589286
rect 364156 589222 364208 589228
rect 364432 589280 364484 589286
rect 364432 589222 364484 589228
rect 364168 579737 364196 589222
rect 429672 582486 429700 589290
rect 494164 589286 494192 591926
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 493876 589280 493928 589286
rect 493876 589222 493928 589228
rect 494152 589280 494204 589286
rect 494152 589222 494204 589228
rect 429660 582480 429712 582486
rect 429660 582422 429712 582428
rect 429568 582344 429620 582350
rect 429568 582286 429620 582292
rect 364154 579728 364210 579737
rect 364154 579663 364210 579672
rect 364338 579728 364394 579737
rect 364338 579663 364394 579672
rect 364352 572642 364380 579663
rect 429580 572642 429608 582286
rect 493888 579737 493916 589222
rect 559392 582486 559420 589290
rect 559380 582480 559432 582486
rect 559380 582422 559432 582428
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 493874 579728 493930 579737
rect 493874 579663 493930 579672
rect 494058 579728 494114 579737
rect 494058 579663 494114 579672
rect 364352 572614 364472 572642
rect 351920 567248 351972 567254
rect 351920 567190 351972 567196
rect 351932 546394 351960 567190
rect 364444 563122 364472 572614
rect 429396 572614 429608 572642
rect 494072 572642 494100 579663
rect 559300 572642 559328 582286
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 494072 572614 494192 572642
rect 429396 569922 429424 572614
rect 429304 569894 429424 569922
rect 429304 563174 429332 569894
rect 429292 563168 429344 563174
rect 364444 563094 364564 563122
rect 429292 563110 429344 563116
rect 494164 563122 494192 572614
rect 559116 572614 559328 572642
rect 559116 569922 559144 572614
rect 559024 569894 559144 569922
rect 559024 563174 559052 569894
rect 559012 563168 559064 563174
rect 494164 563094 494284 563122
rect 559012 563110 559064 563116
rect 364536 557546 364564 563094
rect 429292 563032 429344 563038
rect 429292 562974 429344 562980
rect 429304 560266 429332 562974
rect 364352 557518 364564 557546
rect 429212 560238 429332 560266
rect 357440 552152 357492 552158
rect 357440 552094 357492 552100
rect 355508 549024 355560 549030
rect 355508 548966 355560 548972
rect 349172 546366 349752 546394
rect 351932 546366 352328 546394
rect 349724 546258 349752 546366
rect 352300 546258 352328 546366
rect 349724 546230 350382 546258
rect 352300 546230 352958 546258
rect 355520 546244 355548 548966
rect 357452 546258 357480 552094
rect 364352 550118 364380 557518
rect 429212 553450 429240 560238
rect 494256 557546 494284 563094
rect 559012 563032 559064 563038
rect 559012 562974 559064 562980
rect 559024 560250 559052 562974
rect 559012 560244 559064 560250
rect 559012 560186 559064 560192
rect 494072 557518 494284 557546
rect 429200 553444 429252 553450
rect 429200 553386 429252 553392
rect 429200 550656 429252 550662
rect 429200 550598 429252 550604
rect 364340 550112 364392 550118
rect 364340 550054 364392 550060
rect 429212 550050 429240 550598
rect 429200 550044 429252 550050
rect 429200 549986 429252 549992
rect 494072 549982 494100 557518
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 577504 552084 577556 552090
rect 577504 552026 577556 552032
rect 559104 550656 559156 550662
rect 559104 550598 559156 550604
rect 494060 549976 494112 549982
rect 494060 549918 494112 549924
rect 559116 549914 559144 550598
rect 559104 549908 559156 549914
rect 559104 549850 559156 549856
rect 440882 549264 440938 549273
rect 440882 549199 440938 549208
rect 449532 549228 449584 549234
rect 365904 548956 365956 548962
rect 365904 548898 365956 548904
rect 357452 546230 358110 546258
rect 365916 546244 365944 548898
rect 371056 548888 371108 548894
rect 371056 548830 371108 548836
rect 407302 548856 407358 548865
rect 368480 548820 368532 548826
rect 368480 548762 368532 548768
rect 368492 546244 368520 548762
rect 371068 546244 371096 548830
rect 407302 548791 407358 548800
rect 373632 548752 373684 548758
rect 373632 548694 373684 548700
rect 373644 546244 373672 548694
rect 376208 548684 376260 548690
rect 376208 548626 376260 548632
rect 376220 546244 376248 548626
rect 378784 548616 378836 548622
rect 378784 548558 378836 548564
rect 378796 546244 378824 548558
rect 381360 548548 381412 548554
rect 381360 548490 381412 548496
rect 381372 546244 381400 548490
rect 384028 548480 384080 548486
rect 384028 548422 384080 548428
rect 384040 546244 384068 548422
rect 389180 548412 389232 548418
rect 389180 548354 389232 548360
rect 389192 546244 389220 548354
rect 391756 548344 391808 548350
rect 391756 548286 391808 548292
rect 391768 546244 391796 548286
rect 394332 548276 394384 548282
rect 394332 548218 394384 548224
rect 394344 546244 394372 548218
rect 396908 548208 396960 548214
rect 396908 548150 396960 548156
rect 396920 546244 396948 548150
rect 404636 548140 404688 548146
rect 404636 548082 404688 548088
rect 399484 548072 399536 548078
rect 399484 548014 399536 548020
rect 399496 546244 399524 548014
rect 404648 546244 404676 548082
rect 407316 546244 407344 548791
rect 415030 548584 415086 548593
rect 415030 548519 415086 548528
rect 409880 547936 409932 547942
rect 409880 547878 409932 547884
rect 409892 546244 409920 547878
rect 415044 546244 415072 548519
rect 435730 548312 435786 548321
rect 435730 548247 435786 548256
rect 425334 548040 425390 548049
rect 420184 548004 420236 548010
rect 425334 547975 425390 547984
rect 420184 547946 420236 547952
rect 420196 546244 420224 547946
rect 425348 546244 425376 547975
rect 435744 546244 435772 548247
rect 440896 546244 440924 549199
rect 449532 549170 449584 549176
rect 449348 549092 449400 549098
rect 449348 549034 449400 549040
rect 336752 546094 337502 546122
rect 401704 545562 402086 545578
rect 149704 545556 149756 545562
rect 149704 545498 149756 545504
rect 401692 545556 402086 545562
rect 401744 545550 402086 545556
rect 401692 545498 401744 545504
rect 71044 242888 71096 242894
rect 71044 242830 71096 242836
rect 42064 242820 42116 242826
rect 42064 242762 42116 242768
rect 35164 242480 35216 242486
rect 35164 242422 35216 242428
rect 31024 242412 31076 242418
rect 31024 242354 31076 242360
rect 24124 242344 24176 242350
rect 24124 242286 24176 242292
rect 21364 64864 21416 64870
rect 21364 64806 21416 64812
rect 23112 7608 23164 7614
rect 23112 7550 23164 7556
rect 18328 6384 18380 6390
rect 18328 6326 18380 6332
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 14844 480 14872 3946
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16040 480 16068 3674
rect 17328 2530 17356 5034
rect 17236 2502 17356 2530
rect 17236 480 17264 2502
rect 18340 480 18368 6326
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19536 480 19564 3538
rect 20732 480 20760 3606
rect 21928 480 21956 5102
rect 23124 480 23152 7550
rect 24136 3738 24164 242286
rect 28264 242276 28316 242282
rect 28264 242218 28316 242224
rect 27894 8936 27950 8945
rect 27894 8871 27950 8880
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 24308 3936 24360 3942
rect 24308 3878 24360 3884
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24320 480 24348 3878
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 25516 480 25544 3742
rect 26712 480 26740 5170
rect 27908 480 27936 8871
rect 28276 3942 28304 242218
rect 30288 5296 30340 5302
rect 30288 5238 30340 5244
rect 28264 3936 28316 3942
rect 28264 3878 28316 3884
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 29104 480 29132 3674
rect 30300 480 30328 5238
rect 31036 3806 31064 242354
rect 31484 8968 31536 8974
rect 31484 8910 31536 8916
rect 31024 3800 31076 3806
rect 31024 3742 31076 3748
rect 31496 480 31524 8910
rect 33876 5364 33928 5370
rect 33876 5306 33928 5312
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 32692 480 32720 3334
rect 33888 480 33916 5306
rect 34980 3800 35032 3806
rect 34980 3742 35032 3748
rect 34992 480 35020 3742
rect 35176 3398 35204 242422
rect 40960 6452 41012 6458
rect 40960 6394 41012 6400
rect 37370 6216 37426 6225
rect 37370 6151 37426 6160
rect 36176 3868 36228 3874
rect 36176 3810 36228 3816
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36188 480 36216 3810
rect 37384 480 37412 6151
rect 39764 4140 39816 4146
rect 39764 4082 39816 4088
rect 38568 3324 38620 3330
rect 38568 3266 38620 3272
rect 38580 480 38608 3266
rect 39776 480 39804 4082
rect 40972 480 41000 6394
rect 42076 4146 42104 242762
rect 70674 7576 70730 7585
rect 70674 7511 70730 7520
rect 67180 6860 67232 6866
rect 67180 6802 67232 6808
rect 63592 6792 63644 6798
rect 63592 6734 63644 6740
rect 60004 6724 60056 6730
rect 60004 6666 60056 6672
rect 56416 6656 56468 6662
rect 56416 6598 56468 6604
rect 52828 6588 52880 6594
rect 52828 6530 52880 6536
rect 49332 6520 49384 6526
rect 49332 6462 49384 6468
rect 44546 6352 44602 6361
rect 44546 6287 44602 6296
rect 42064 4140 42116 4146
rect 42064 4082 42116 4088
rect 43352 4004 43404 4010
rect 43352 3946 43404 3952
rect 42156 3936 42208 3942
rect 42156 3878 42208 3884
rect 42168 480 42196 3878
rect 43364 480 43392 3946
rect 44560 480 44588 6287
rect 48136 5432 48188 5438
rect 48136 5374 48188 5380
rect 45744 3256 45796 3262
rect 45744 3198 45796 3204
rect 45756 480 45784 3198
rect 46940 3052 46992 3058
rect 46940 2994 46992 3000
rect 46952 480 46980 2994
rect 48148 480 48176 5374
rect 49344 480 49372 6462
rect 51632 5500 51684 5506
rect 51632 5442 51684 5448
rect 50528 3188 50580 3194
rect 50528 3130 50580 3136
rect 50540 480 50568 3130
rect 51644 480 51672 5442
rect 52840 480 52868 6530
rect 55220 4752 55272 4758
rect 55220 4694 55272 4700
rect 54024 4072 54076 4078
rect 54024 4014 54076 4020
rect 54036 480 54064 4014
rect 55232 480 55260 4694
rect 56428 480 56456 6598
rect 58808 4684 58860 4690
rect 58808 4626 58860 4632
rect 57612 3120 57664 3126
rect 57612 3062 57664 3068
rect 57624 480 57652 3062
rect 58820 480 58848 4626
rect 60016 480 60044 6666
rect 62396 4548 62448 4554
rect 62396 4490 62448 4496
rect 61200 4140 61252 4146
rect 61200 4082 61252 4088
rect 61212 480 61240 4082
rect 62408 480 62436 4490
rect 63604 480 63632 6734
rect 65984 4616 66036 4622
rect 65984 4558 66036 4564
rect 64788 2916 64840 2922
rect 64788 2858 64840 2864
rect 64800 480 64828 2858
rect 65996 480 66024 4558
rect 67192 480 67220 6802
rect 69480 4480 69532 4486
rect 69480 4422 69532 4428
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 68296 480 68324 3334
rect 69492 480 69520 4422
rect 70688 480 70716 7511
rect 71056 3330 71084 242830
rect 103428 242820 103480 242826
rect 103428 242762 103480 242768
rect 86224 242752 86276 242758
rect 86224 242694 86276 242700
rect 77944 242072 77996 242078
rect 77944 242014 77996 242020
rect 75184 242004 75236 242010
rect 75184 241946 75236 241952
rect 74264 9036 74316 9042
rect 74264 8978 74316 8984
rect 73068 4412 73120 4418
rect 73068 4354 73120 4360
rect 71044 3324 71096 3330
rect 71044 3266 71096 3272
rect 71872 2984 71924 2990
rect 71872 2926 71924 2932
rect 71884 480 71912 2926
rect 73080 480 73108 4354
rect 74276 480 74304 8978
rect 75196 3262 75224 241946
rect 77852 9104 77904 9110
rect 77852 9046 77904 9052
rect 76656 4344 76708 4350
rect 76656 4286 76708 4292
rect 75460 3324 75512 3330
rect 75460 3266 75512 3272
rect 75184 3256 75236 3262
rect 75184 3198 75236 3204
rect 75472 480 75500 3266
rect 76668 480 76696 4286
rect 77864 480 77892 9046
rect 77956 3194 77984 242014
rect 84844 241868 84896 241874
rect 84844 241810 84896 241816
rect 81440 9172 81492 9178
rect 81440 9114 81492 9120
rect 80244 4276 80296 4282
rect 80244 4218 80296 4224
rect 77944 3188 77996 3194
rect 77944 3130 77996 3136
rect 79048 2848 79100 2854
rect 79048 2790 79100 2796
rect 79060 480 79088 2790
rect 80256 480 80284 4218
rect 81452 480 81480 9114
rect 83832 4208 83884 4214
rect 83832 4150 83884 4156
rect 82636 3256 82688 3262
rect 82636 3198 82688 3204
rect 82648 480 82676 3198
rect 83844 480 83872 4150
rect 84856 3126 84884 241810
rect 84936 9240 84988 9246
rect 84936 9182 84988 9188
rect 84844 3120 84896 3126
rect 84844 3062 84896 3068
rect 84948 480 84976 9182
rect 86132 3120 86184 3126
rect 86132 3062 86184 3068
rect 86144 480 86172 3062
rect 86236 2990 86264 242694
rect 88984 242684 89036 242690
rect 88984 242626 89036 242632
rect 88524 9308 88576 9314
rect 88524 9250 88576 9256
rect 87328 7676 87380 7682
rect 87328 7618 87380 7624
rect 86224 2984 86276 2990
rect 86224 2926 86276 2932
rect 87340 480 87368 7618
rect 88536 480 88564 9250
rect 88996 2854 89024 242626
rect 93124 242616 93176 242622
rect 93124 242558 93176 242564
rect 92112 9376 92164 9382
rect 92112 9318 92164 9324
rect 90916 7744 90968 7750
rect 90916 7686 90968 7692
rect 89720 3188 89772 3194
rect 89720 3130 89772 3136
rect 88984 2848 89036 2854
rect 88984 2790 89036 2796
rect 89732 480 89760 3130
rect 90928 480 90956 7686
rect 92124 480 92152 9318
rect 93136 3194 93164 242558
rect 103440 242146 103468 242762
rect 113180 242548 113232 242554
rect 113180 242490 113232 242496
rect 122748 242548 122800 242554
rect 122748 242490 122800 242496
rect 98644 242140 98696 242146
rect 98644 242082 98696 242088
rect 103428 242140 103480 242146
rect 103428 242082 103480 242088
rect 104808 242140 104860 242146
rect 104808 242082 104860 242088
rect 95884 241664 95936 241670
rect 95884 241606 95936 241612
rect 95700 9444 95752 9450
rect 95700 9386 95752 9392
rect 94504 7812 94556 7818
rect 94504 7754 94556 7760
rect 93858 5400 93914 5409
rect 93858 5335 93860 5344
rect 93912 5335 93914 5344
rect 93860 5306 93912 5312
rect 93124 3188 93176 3194
rect 93124 3130 93176 3136
rect 93308 3120 93360 3126
rect 93308 3062 93360 3068
rect 93320 480 93348 3062
rect 94516 480 94544 7754
rect 95712 480 95740 9386
rect 95896 3058 95924 241606
rect 98092 7880 98144 7886
rect 98092 7822 98144 7828
rect 95884 3052 95936 3058
rect 95884 2994 95936 3000
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 96908 480 96936 2994
rect 98104 480 98132 7822
rect 98656 3058 98684 242082
rect 102784 9512 102836 9518
rect 102784 9454 102836 9460
rect 101588 7948 101640 7954
rect 101588 7890 101640 7896
rect 99288 5636 99340 5642
rect 99288 5578 99340 5584
rect 98644 3052 98696 3058
rect 98644 2994 98696 3000
rect 99300 480 99328 5578
rect 100484 2984 100536 2990
rect 100484 2926 100536 2932
rect 100496 480 100524 2926
rect 101600 480 101628 7890
rect 102796 480 102824 9454
rect 103426 5400 103482 5409
rect 103426 5335 103428 5344
rect 103480 5335 103482 5344
rect 103428 5306 103480 5312
rect 104820 3058 104848 242082
rect 111708 241936 111760 241942
rect 111708 241878 111760 241884
rect 106924 241596 106976 241602
rect 106924 241538 106976 241544
rect 106372 9580 106424 9586
rect 106372 9522 106424 9528
rect 105176 8016 105228 8022
rect 105176 7958 105228 7964
rect 103980 3052 104032 3058
rect 103980 2994 104032 3000
rect 104808 3052 104860 3058
rect 104808 2994 104860 3000
rect 103992 480 104020 2994
rect 105188 480 105216 7958
rect 106384 480 106412 9522
rect 106936 2922 106964 241538
rect 109960 9648 110012 9654
rect 109960 9590 110012 9596
rect 108764 8084 108816 8090
rect 108764 8026 108816 8032
rect 106924 2916 106976 2922
rect 106924 2858 106976 2864
rect 107568 2848 107620 2854
rect 107568 2790 107620 2796
rect 107580 480 107608 2790
rect 108776 480 108804 8026
rect 109972 480 110000 9590
rect 111720 3058 111748 241878
rect 113192 241534 113220 242490
rect 122760 241890 122788 242490
rect 122668 241862 122788 241890
rect 115848 241800 115900 241806
rect 115848 241742 115900 241748
rect 113180 241528 113232 241534
rect 113180 241470 113232 241476
rect 112352 8152 112404 8158
rect 112352 8094 112404 8100
rect 111156 3052 111208 3058
rect 111156 2994 111208 3000
rect 111708 3052 111760 3058
rect 111708 2994 111760 3000
rect 111168 480 111196 2994
rect 112364 480 112392 8094
rect 113548 5568 113600 5574
rect 113548 5510 113600 5516
rect 113178 5400 113234 5409
rect 113178 5335 113180 5344
rect 113232 5335 113234 5344
rect 113180 5306 113232 5312
rect 113560 480 113588 5510
rect 115860 2922 115888 241742
rect 122668 241534 122696 241862
rect 122748 241732 122800 241738
rect 122748 241674 122800 241680
rect 122656 241528 122708 241534
rect 122656 241470 122708 241476
rect 117136 8900 117188 8906
rect 117136 8842 117188 8848
rect 115940 8220 115992 8226
rect 115940 8162 115992 8168
rect 114744 2916 114796 2922
rect 114744 2858 114796 2864
rect 115848 2916 115900 2922
rect 115848 2858 115900 2864
rect 114756 480 114784 2858
rect 115952 480 115980 8162
rect 117148 480 117176 8842
rect 120632 8832 120684 8838
rect 120632 8774 120684 8780
rect 119436 8288 119488 8294
rect 119436 8230 119488 8236
rect 118240 2848 118292 2854
rect 118240 2790 118292 2796
rect 118252 480 118280 2790
rect 119448 480 119476 8230
rect 120644 480 120672 8774
rect 122654 5400 122710 5409
rect 122654 5335 122656 5344
rect 122708 5335 122710 5344
rect 122656 5306 122708 5312
rect 122760 2922 122788 241674
rect 149060 239352 149112 239358
rect 149060 239294 149112 239300
rect 124220 8764 124272 8770
rect 124220 8706 124272 8712
rect 123024 7540 123076 7546
rect 123024 7482 123076 7488
rect 121828 2916 121880 2922
rect 121828 2858 121880 2864
rect 122748 2916 122800 2922
rect 122748 2858 122800 2864
rect 121840 480 121868 2858
rect 123036 480 123064 7482
rect 124232 480 124260 8706
rect 131396 8696 131448 8702
rect 131396 8638 131448 8644
rect 127808 7472 127860 7478
rect 127808 7414 127860 7420
rect 126612 7404 126664 7410
rect 126612 7346 126664 7352
rect 125416 2916 125468 2922
rect 125416 2858 125468 2864
rect 125428 480 125456 2858
rect 126624 480 126652 7346
rect 127820 480 127848 7414
rect 130200 7336 130252 7342
rect 130200 7278 130252 7284
rect 129004 6112 129056 6118
rect 129004 6054 129056 6060
rect 129016 480 129044 6054
rect 130212 480 130240 7278
rect 131408 480 131436 8638
rect 134892 8628 134944 8634
rect 134892 8570 134944 8576
rect 133788 7268 133840 7274
rect 133788 7210 133840 7216
rect 132592 6044 132644 6050
rect 132592 5986 132644 5992
rect 132498 5400 132554 5409
rect 132498 5335 132500 5344
rect 132552 5335 132554 5344
rect 132500 5306 132552 5312
rect 132604 480 132632 5986
rect 133800 480 133828 7210
rect 134904 480 134932 8570
rect 138480 8560 138532 8566
rect 138480 8502 138532 8508
rect 137284 7200 137336 7206
rect 137284 7142 137336 7148
rect 136088 5976 136140 5982
rect 136088 5918 136140 5924
rect 136100 480 136128 5918
rect 137296 480 137324 7142
rect 138492 480 138520 8502
rect 142068 8492 142120 8498
rect 142068 8434 142120 8440
rect 140872 7132 140924 7138
rect 140872 7074 140924 7080
rect 139676 5908 139728 5914
rect 139676 5850 139728 5856
rect 139688 480 139716 5850
rect 140884 480 140912 7074
rect 141974 5400 142030 5409
rect 141974 5335 141976 5344
rect 142028 5335 142030 5344
rect 141976 5306 142028 5312
rect 142080 480 142108 8434
rect 145656 8424 145708 8430
rect 145656 8366 145708 8372
rect 144460 7064 144512 7070
rect 144460 7006 144512 7012
rect 143264 5840 143316 5846
rect 143264 5782 143316 5788
rect 142160 5024 142212 5030
rect 142158 4992 142160 5001
rect 142212 4992 142214 5001
rect 142158 4927 142214 4936
rect 143276 480 143304 5782
rect 144472 480 144500 7006
rect 145668 480 145696 8366
rect 148048 6996 148100 7002
rect 148048 6938 148100 6944
rect 146852 5772 146904 5778
rect 146852 5714 146904 5720
rect 146864 480 146892 5714
rect 148060 480 148088 6938
rect 149072 4894 149100 239294
rect 149716 223582 149744 545498
rect 184756 545488 184808 545494
rect 177146 545426 177528 545442
rect 449256 545488 449308 545494
rect 184808 545436 184874 545442
rect 184756 545430 184874 545436
rect 449256 545430 449308 545436
rect 177146 545420 177540 545426
rect 177146 545414 177488 545420
rect 184768 545414 184874 545430
rect 449164 545420 449216 545426
rect 177488 545362 177540 545368
rect 449164 545362 449216 545368
rect 242072 545352 242124 545358
rect 241730 545300 242072 545306
rect 422482 545320 422538 545329
rect 241730 545294 242124 545300
rect 241730 545278 242112 545294
rect 363064 545290 363354 545306
rect 363052 545284 363354 545290
rect 363104 545278 363354 545284
rect 422538 545278 422786 545306
rect 422482 545255 422538 545264
rect 363052 545226 363104 545232
rect 192852 545216 192904 545222
rect 187450 545154 187648 545170
rect 192602 545164 192852 545170
rect 192602 545158 192904 545164
rect 430486 545184 430542 545193
rect 187450 545148 187660 545154
rect 187450 545142 187608 545148
rect 192602 545142 192892 545158
rect 430542 545142 430606 545170
rect 430486 545119 430542 545128
rect 187608 545090 187660 545096
rect 236920 544944 236972 544950
rect 228850 544882 229048 544898
rect 236578 544892 236920 544898
rect 236578 544886 236972 544892
rect 449072 544944 449124 544950
rect 449072 544886 449124 544892
rect 228850 544876 229060 544882
rect 228850 544870 229008 544876
rect 236578 544870 236960 544886
rect 229008 544818 229060 544824
rect 216128 544808 216180 544814
rect 161598 544746 161888 544762
rect 164068 544746 164174 544762
rect 161598 544740 161900 544746
rect 161598 544734 161848 544740
rect 161848 544682 161900 544688
rect 164056 544740 164174 544746
rect 164108 544734 164174 544740
rect 169326 544746 169616 544762
rect 171902 544746 172192 544762
rect 174570 544746 174952 544762
rect 179722 544746 180104 544762
rect 182298 544746 182680 544762
rect 195178 544746 195560 544762
rect 200422 544746 200712 544762
rect 215878 544756 216128 544762
rect 215878 544750 216180 544756
rect 169326 544740 169628 544746
rect 169326 544734 169576 544740
rect 164056 544682 164108 544688
rect 171902 544740 172204 544746
rect 171902 544734 172152 544740
rect 169576 544682 169628 544688
rect 174570 544740 174964 544746
rect 174570 544734 174912 544740
rect 172152 544682 172204 544688
rect 179722 544740 180116 544746
rect 179722 544734 180064 544740
rect 174912 544682 174964 544688
rect 182298 544740 182692 544746
rect 182298 544734 182640 544740
rect 180064 544682 180116 544688
rect 195178 544740 195572 544746
rect 195178 544734 195520 544740
rect 182640 544682 182692 544688
rect 200422 544740 200724 544746
rect 200422 544734 200672 544740
rect 195520 544682 195572 544688
rect 215878 544734 216168 544750
rect 234002 544746 234384 544762
rect 234002 544740 234396 544746
rect 234002 544734 234344 544740
rect 200672 544682 200724 544688
rect 234344 544682 234396 544688
rect 360476 544672 360528 544678
rect 151542 544640 151598 544649
rect 151294 544598 151542 544626
rect 154026 544640 154082 544649
rect 153870 544598 154026 544626
rect 151542 544575 151598 544584
rect 203154 544640 203210 544649
rect 202998 544598 203154 544626
rect 154026 544575 154082 544584
rect 203154 544575 203210 544584
rect 205454 544640 205510 544649
rect 208030 544640 208086 544649
rect 205510 544598 205574 544626
rect 205454 544575 205510 544584
rect 213458 544640 213514 544649
rect 208086 544598 208150 544626
rect 213302 544598 213458 544626
rect 208030 544575 208086 544584
rect 221278 544640 221334 544649
rect 221122 544598 221278 544626
rect 213458 544575 213514 544584
rect 231582 544640 231638 544649
rect 231426 544598 231582 544626
rect 221278 544575 221334 544584
rect 412180 544672 412232 544678
rect 386510 544640 386566 544649
rect 360528 544620 360778 544626
rect 360476 544614 360778 544620
rect 360488 544598 360778 544614
rect 231582 544575 231638 544584
rect 386566 544598 386630 544626
rect 417332 544672 417384 544678
rect 412232 544620 412482 544626
rect 412180 544614 412482 544620
rect 427820 544672 427872 544678
rect 417384 544620 417634 544626
rect 417332 544614 417634 544620
rect 432788 544672 432840 544678
rect 427872 544620 427938 544626
rect 427820 544614 427938 544620
rect 438216 544672 438268 544678
rect 432840 544620 433182 544626
rect 432788 544614 433182 544620
rect 443092 544672 443144 544678
rect 438268 544620 438334 544626
rect 438216 544614 438334 544620
rect 443144 544620 443486 544626
rect 443092 544614 443486 544620
rect 412192 544598 412482 544614
rect 417344 544598 417634 544614
rect 427832 544598 427938 544614
rect 432800 544598 433182 544614
rect 438228 544598 438334 544614
rect 443104 544598 443486 544614
rect 386510 544575 386566 544584
rect 449084 534070 449112 544886
rect 449072 534064 449124 534070
rect 449072 534006 449124 534012
rect 163240 244174 163714 244202
rect 178512 244174 178986 244202
rect 179708 244174 180182 244202
rect 185228 244174 185702 244202
rect 190748 244174 191130 244202
rect 192588 244174 192970 244202
rect 194980 244174 195454 244202
rect 196268 244174 196650 244202
rect 206020 244174 206494 244202
rect 207216 244174 207690 244202
rect 211540 244174 211922 244202
rect 223684 244174 224158 244202
rect 226812 244174 227194 244202
rect 229204 244174 229678 244202
rect 229848 244174 230322 244202
rect 234724 244174 235198 244202
rect 236564 244174 237038 244202
rect 237760 244174 238234 244202
rect 245764 244174 246146 244202
rect 283576 244174 284050 244202
rect 303816 244174 304198 244202
rect 345782 244174 346256 244202
rect 422786 244174 423260 244202
rect 149992 244038 150282 244066
rect 150452 244038 150834 244066
rect 151188 244038 151478 244066
rect 151924 244038 152030 244066
rect 152200 244038 152674 244066
rect 149992 239358 150020 244038
rect 149980 239352 150032 239358
rect 149980 239294 150032 239300
rect 149704 223576 149756 223582
rect 149704 223518 149756 223524
rect 150452 6236 150480 244038
rect 151188 239358 151216 244038
rect 150716 239352 150768 239358
rect 150716 239294 150768 239300
rect 151176 239352 151228 239358
rect 151176 239294 151228 239300
rect 150728 227066 150756 239294
rect 151726 237144 151782 237153
rect 151726 237079 151782 237088
rect 150728 227038 150940 227066
rect 150912 209846 150940 227038
rect 151740 221105 151768 237079
rect 151726 221096 151782 221105
rect 151726 221031 151782 221040
rect 150808 209840 150860 209846
rect 150808 209782 150860 209788
rect 150900 209840 150952 209846
rect 150900 209782 150952 209788
rect 150820 205698 150848 209782
rect 151634 206272 151690 206281
rect 151634 206207 151690 206216
rect 150808 205692 150860 205698
rect 150808 205634 150860 205640
rect 150808 205556 150860 205562
rect 150808 205498 150860 205504
rect 150820 201482 150848 205498
rect 150808 201476 150860 201482
rect 150808 201418 150860 201424
rect 151648 193225 151676 206207
rect 151634 193216 151690 193225
rect 151634 193151 151690 193160
rect 151818 193216 151874 193225
rect 151818 193151 151874 193160
rect 151832 183598 151860 193151
rect 150808 183592 150860 183598
rect 150808 183534 150860 183540
rect 151820 183592 151872 183598
rect 151820 183534 151872 183540
rect 150820 182170 150848 183534
rect 150808 182164 150860 182170
rect 150808 182106 150860 182112
rect 151450 177304 151506 177313
rect 151450 177239 151506 177248
rect 150716 173732 150768 173738
rect 150716 173674 150768 173680
rect 150728 164393 150756 173674
rect 151464 165481 151492 177239
rect 151450 165472 151506 165481
rect 151450 165407 151506 165416
rect 150714 164384 150770 164393
rect 150714 164319 150770 164328
rect 150806 164248 150862 164257
rect 150806 164183 150862 164192
rect 150820 156618 150848 164183
rect 150728 156590 150848 156618
rect 150728 147098 150756 156590
rect 150728 147070 150848 147098
rect 150820 142202 150848 147070
rect 150728 142174 150848 142202
rect 150728 140758 150756 142174
rect 150716 140752 150768 140758
rect 150716 140694 150768 140700
rect 150808 131164 150860 131170
rect 150808 131106 150860 131112
rect 150820 121394 150848 131106
rect 150728 121366 150848 121394
rect 150728 116346 150756 121366
rect 150716 116340 150768 116346
rect 150716 116282 150768 116288
rect 151542 112976 151598 112985
rect 151542 112911 151598 112920
rect 151556 104281 151584 112911
rect 151542 104272 151598 104281
rect 151542 104207 151598 104216
rect 150808 103556 150860 103562
rect 150808 103498 150860 103504
rect 150820 103442 150848 103498
rect 150820 103414 151032 103442
rect 151004 92721 151032 103414
rect 151082 92848 151138 92857
rect 151082 92783 151138 92792
rect 150990 92712 151046 92721
rect 150990 92647 151046 92656
rect 150714 92576 150770 92585
rect 150714 92511 150770 92520
rect 150728 92478 150756 92511
rect 150716 92472 150768 92478
rect 150716 92414 150768 92420
rect 150992 92472 151044 92478
rect 150992 92414 151044 92420
rect 151004 78010 151032 92414
rect 151096 91361 151124 92783
rect 151082 91352 151138 91361
rect 151082 91287 151138 91296
rect 151358 81424 151414 81433
rect 151358 81359 151414 81368
rect 150820 77982 151032 78010
rect 150820 70394 150848 77982
rect 151372 71913 151400 81359
rect 151358 71904 151414 71913
rect 151358 71839 151414 71848
rect 150728 70366 150848 70394
rect 150728 70310 150756 70366
rect 150716 70304 150768 70310
rect 150716 70246 150768 70252
rect 150716 64864 150768 64870
rect 150716 64806 150768 64812
rect 150728 60738 150756 64806
rect 150728 60710 150848 60738
rect 150820 51218 150848 60710
rect 150728 51190 150848 51218
rect 150728 51105 150756 51190
rect 150530 51096 150586 51105
rect 150530 51031 150586 51040
rect 150714 51096 150770 51105
rect 150714 51031 150770 51040
rect 150544 45694 150572 51031
rect 150532 45688 150584 45694
rect 150532 45630 150584 45636
rect 150716 45688 150768 45694
rect 150716 45630 150768 45636
rect 150728 33153 150756 45630
rect 150530 33144 150586 33153
rect 150530 33079 150586 33088
rect 150714 33144 150770 33153
rect 150714 33079 150770 33088
rect 150544 28354 150572 33079
rect 150532 28348 150584 28354
rect 150532 28290 150584 28296
rect 150716 28348 150768 28354
rect 150716 28290 150768 28296
rect 150728 23474 150756 28290
rect 150728 23446 150848 23474
rect 150820 16538 150848 23446
rect 150820 16510 150940 16538
rect 150912 6934 150940 16510
rect 150808 6928 150860 6934
rect 150808 6870 150860 6876
rect 150900 6928 150952 6934
rect 150900 6870 150952 6876
rect 150452 6208 150572 6236
rect 150440 5704 150492 5710
rect 150440 5646 150492 5652
rect 149060 4888 149112 4894
rect 149060 4830 149112 4836
rect 149244 4888 149296 4894
rect 149244 4830 149296 4836
rect 149256 480 149284 4830
rect 150452 480 150480 5646
rect 150544 4826 150572 6208
rect 150820 4962 150848 6870
rect 151924 6186 151952 244038
rect 152200 239306 152228 244038
rect 153304 242185 153332 244052
rect 153488 244038 153870 244066
rect 154040 244038 154514 244066
rect 154684 244038 155158 244066
rect 155328 244038 155710 244066
rect 155972 244038 156354 244066
rect 156524 244038 156998 244066
rect 153290 242176 153346 242185
rect 153290 242111 153346 242120
rect 153488 239306 153516 244038
rect 152016 239278 152228 239306
rect 153212 239278 153516 239306
rect 152016 234546 152044 239278
rect 152016 234518 152136 234546
rect 152002 201376 152058 201385
rect 152002 201311 152058 201320
rect 152016 196625 152044 201311
rect 152002 196616 152058 196625
rect 152002 196551 152058 196560
rect 152108 196058 152136 234518
rect 152738 215248 152794 215257
rect 152738 215183 152794 215192
rect 152752 208321 152780 215183
rect 152738 208312 152794 208321
rect 152738 208247 152794 208256
rect 152016 196030 152136 196058
rect 152016 193225 152044 196030
rect 152002 193216 152058 193225
rect 152002 193151 152058 193160
rect 152004 183592 152056 183598
rect 152004 183534 152056 183540
rect 152016 182170 152044 183534
rect 152004 182164 152056 182170
rect 152004 182106 152056 182112
rect 152188 182164 152240 182170
rect 152188 182106 152240 182112
rect 152200 164286 152228 182106
rect 152004 164280 152056 164286
rect 152004 164222 152056 164228
rect 152188 164280 152240 164286
rect 152188 164222 152240 164228
rect 152016 142118 152044 164222
rect 152004 142112 152056 142118
rect 152004 142054 152056 142060
rect 152188 142112 152240 142118
rect 152188 142054 152240 142060
rect 152200 140758 152228 142054
rect 152188 140752 152240 140758
rect 152188 140694 152240 140700
rect 152188 131164 152240 131170
rect 152188 131106 152240 131112
rect 152200 124386 152228 131106
rect 152108 124358 152228 124386
rect 152108 122874 152136 124358
rect 152004 122868 152056 122874
rect 152004 122810 152056 122816
rect 152096 122868 152148 122874
rect 152096 122810 152148 122816
rect 152016 121446 152044 122810
rect 152004 121440 152056 121446
rect 152004 121382 152056 121388
rect 152004 111852 152056 111858
rect 152004 111794 152056 111800
rect 152016 102134 152044 111794
rect 152004 102128 152056 102134
rect 152004 102070 152056 102076
rect 152004 92540 152056 92546
rect 152004 92482 152056 92488
rect 152016 82822 152044 92482
rect 152004 82816 152056 82822
rect 152004 82758 152056 82764
rect 152004 73228 152056 73234
rect 152004 73170 152056 73176
rect 152016 26314 152044 73170
rect 152004 26308 152056 26314
rect 152004 26250 152056 26256
rect 152096 26308 152148 26314
rect 152096 26250 152148 26256
rect 152108 15201 152136 26250
rect 152094 15192 152150 15201
rect 152094 15127 152150 15136
rect 152278 15192 152334 15201
rect 152278 15127 152334 15136
rect 151912 6180 151964 6186
rect 151912 6122 151964 6128
rect 152292 5681 152320 15127
rect 152002 5672 152058 5681
rect 152002 5607 152058 5616
rect 152278 5672 152334 5681
rect 152278 5607 152334 5616
rect 150898 4992 150954 5001
rect 150808 4956 150860 4962
rect 150898 4927 150900 4936
rect 150808 4898 150860 4904
rect 150952 4927 150954 4936
rect 150900 4898 150952 4904
rect 150532 4820 150584 4826
rect 150532 4762 150584 4768
rect 151544 4820 151596 4826
rect 151544 4762 151596 4768
rect 151556 480 151584 4762
rect 152016 3369 152044 5607
rect 152740 5364 152792 5370
rect 152740 5306 152792 5312
rect 152002 3360 152058 3369
rect 152002 3295 152058 3304
rect 152752 480 152780 5306
rect 153212 4962 153240 239278
rect 154040 236994 154068 244038
rect 153396 236966 154068 236994
rect 153396 220833 153424 236966
rect 153382 220824 153438 220833
rect 153382 220759 153438 220768
rect 153566 220824 153622 220833
rect 153566 220759 153622 220768
rect 153580 212242 153608 220759
rect 153396 212214 153608 212242
rect 153396 207754 153424 212214
rect 153304 207726 153424 207754
rect 153304 195922 153332 207726
rect 153304 195894 153424 195922
rect 153396 176746 153424 195894
rect 153304 176718 153424 176746
rect 153304 176610 153332 176718
rect 153304 176582 153424 176610
rect 153396 157434 153424 176582
rect 153304 157406 153424 157434
rect 153304 157298 153332 157406
rect 153304 157270 153424 157298
rect 153396 137986 153424 157270
rect 153396 137958 153608 137986
rect 153580 133929 153608 137958
rect 153382 133920 153438 133929
rect 153382 133855 153384 133864
rect 153436 133855 153438 133864
rect 153566 133920 153622 133929
rect 153566 133855 153622 133864
rect 153384 133826 153436 133832
rect 153384 124228 153436 124234
rect 153384 124170 153436 124176
rect 153396 118810 153424 124170
rect 153396 118782 153516 118810
rect 153488 114646 153516 118782
rect 153476 114640 153528 114646
rect 153476 114582 153528 114588
rect 153292 114572 153344 114578
rect 153292 114514 153344 114520
rect 153304 114442 153332 114514
rect 153292 114436 153344 114442
rect 153292 114378 153344 114384
rect 153384 104916 153436 104922
rect 153384 104858 153436 104864
rect 153396 99482 153424 104858
rect 153384 99476 153436 99482
rect 153384 99418 153436 99424
rect 153384 99340 153436 99346
rect 153384 99282 153436 99288
rect 153396 6254 153424 99282
rect 153384 6248 153436 6254
rect 153384 6190 153436 6196
rect 153936 6180 153988 6186
rect 153936 6122 153988 6128
rect 153200 4956 153252 4962
rect 153200 4898 153252 4904
rect 153948 480 153976 6122
rect 154684 3466 154712 244038
rect 155328 239306 155356 244038
rect 154868 239278 155356 239306
rect 154868 225010 154896 239278
rect 154856 225004 154908 225010
rect 154856 224946 154908 224952
rect 154868 222222 154896 222253
rect 154856 222216 154908 222222
rect 154776 222164 154856 222170
rect 154776 222158 154908 222164
rect 154776 222142 154896 222158
rect 154776 212566 154804 222142
rect 154764 212560 154816 212566
rect 154764 212502 154816 212508
rect 154856 212560 154908 212566
rect 154856 212502 154908 212508
rect 154868 196058 154896 212502
rect 154776 196030 154896 196058
rect 154776 183569 154804 196030
rect 154762 183560 154818 183569
rect 154762 183495 154818 183504
rect 154946 183560 155002 183569
rect 154946 183495 155002 183504
rect 154960 174010 154988 183495
rect 154856 174004 154908 174010
rect 154856 173946 154908 173952
rect 154948 174004 155000 174010
rect 154948 173946 155000 173952
rect 154868 173913 154896 173946
rect 154854 173904 154910 173913
rect 154854 173839 154910 173848
rect 155038 173904 155094 173913
rect 155038 173839 155094 173848
rect 155052 164257 155080 173839
rect 154854 164248 154910 164257
rect 154854 164183 154910 164192
rect 155038 164248 155094 164257
rect 155038 164183 155094 164192
rect 154868 154578 154896 164183
rect 154776 154550 154896 154578
rect 154776 106214 154804 154550
rect 154764 106208 154816 106214
rect 154764 106150 154816 106156
rect 154764 96756 154816 96762
rect 154764 96698 154816 96704
rect 154776 96626 154804 96698
rect 154764 96620 154816 96626
rect 154764 96562 154816 96568
rect 154948 96620 155000 96626
rect 154948 96562 155000 96568
rect 154960 87009 154988 96562
rect 154762 87000 154818 87009
rect 154762 86935 154818 86944
rect 154946 87000 155002 87009
rect 154946 86935 155002 86944
rect 154776 77246 154804 86935
rect 154764 77240 154816 77246
rect 154764 77182 154816 77188
rect 154764 67652 154816 67658
rect 154764 67594 154816 67600
rect 154776 57934 154804 67594
rect 154764 57928 154816 57934
rect 154764 57870 154816 57876
rect 154764 48408 154816 48414
rect 154764 48350 154816 48356
rect 154776 48278 154804 48350
rect 154764 48272 154816 48278
rect 154764 48214 154816 48220
rect 155040 43716 155092 43722
rect 155040 43658 155092 43664
rect 155052 29050 155080 43658
rect 154868 29022 155080 29050
rect 154868 17950 154896 29022
rect 154856 17944 154908 17950
rect 154856 17886 154908 17892
rect 154856 12436 154908 12442
rect 154856 12378 154908 12384
rect 154868 3534 154896 12378
rect 155224 4956 155276 4962
rect 155224 4898 155276 4904
rect 154856 3528 154908 3534
rect 154856 3470 154908 3476
rect 154672 3460 154724 3466
rect 154672 3402 154724 3408
rect 155236 2530 155264 4898
rect 155972 4865 156000 244038
rect 156524 239306 156552 244038
rect 157536 242214 157564 244052
rect 158180 242350 158208 244052
rect 158746 244038 158852 244066
rect 158168 242344 158220 242350
rect 158168 242286 158220 242292
rect 157524 242208 157576 242214
rect 157524 242150 157576 242156
rect 156156 239278 156552 239306
rect 158720 239352 158772 239358
rect 158720 239294 158772 239300
rect 156156 225010 156184 239278
rect 156144 225004 156196 225010
rect 156144 224946 156196 224952
rect 156144 222216 156196 222222
rect 156144 222158 156196 222164
rect 156156 217410 156184 222158
rect 156064 217382 156184 217410
rect 156064 195922 156092 217382
rect 156064 195894 156184 195922
rect 156156 176662 156184 195894
rect 156144 176656 156196 176662
rect 156144 176598 156196 176604
rect 156144 176520 156196 176526
rect 156144 176462 156196 176468
rect 156156 164218 156184 176462
rect 156144 164212 156196 164218
rect 156144 164154 156196 164160
rect 156144 154624 156196 154630
rect 156144 154566 156196 154572
rect 156156 136218 156184 154566
rect 156156 136190 156368 136218
rect 156340 133929 156368 136190
rect 156142 133920 156198 133929
rect 156142 133855 156144 133864
rect 156196 133855 156198 133864
rect 156326 133920 156382 133929
rect 156326 133855 156382 133864
rect 156144 133826 156196 133832
rect 156144 124228 156196 124234
rect 156144 124170 156196 124176
rect 156156 118794 156184 124170
rect 156144 118788 156196 118794
rect 156144 118730 156196 118736
rect 156144 118652 156196 118658
rect 156144 118594 156196 118600
rect 156156 99482 156184 118594
rect 156144 99476 156196 99482
rect 156144 99418 156196 99424
rect 156144 99340 156196 99346
rect 156144 99282 156196 99288
rect 156156 6322 156184 99282
rect 156328 8356 156380 8362
rect 156328 8298 156380 8304
rect 156144 6316 156196 6322
rect 156144 6258 156196 6264
rect 155958 4856 156014 4865
rect 155958 4791 156014 4800
rect 155144 2502 155264 2530
rect 155144 480 155172 2502
rect 156340 480 156368 8298
rect 157524 6248 157576 6254
rect 157524 6190 157576 6196
rect 157536 480 157564 6190
rect 158732 3602 158760 239294
rect 158824 5098 158852 244038
rect 158916 244038 159390 244066
rect 159744 244038 160034 244066
rect 160204 244038 160586 244066
rect 160756 244038 161230 244066
rect 161584 244038 161874 244066
rect 158916 6390 158944 244038
rect 159744 239358 159772 244038
rect 159732 239352 159784 239358
rect 160204 239340 160232 244038
rect 159732 239294 159784 239300
rect 160112 239312 160232 239340
rect 158904 6384 158956 6390
rect 158904 6326 158956 6332
rect 159916 6316 159968 6322
rect 159916 6258 159968 6264
rect 158812 5092 158864 5098
rect 158812 5034 158864 5040
rect 158996 5024 159048 5030
rect 158996 4966 159048 4972
rect 158720 3596 158772 3602
rect 158720 3538 158772 3544
rect 159008 2530 159036 4966
rect 158732 2502 159036 2530
rect 158732 480 158760 2502
rect 159928 480 159956 6258
rect 160112 3670 160140 239312
rect 160756 239170 160784 244038
rect 160836 241528 160888 241534
rect 160836 241470 160888 241476
rect 160204 239142 160784 239170
rect 160204 5098 160232 239142
rect 160848 236586 160876 241470
rect 160756 236558 160876 236586
rect 160756 5574 160784 236558
rect 161584 7614 161612 244038
rect 162412 242282 162440 244052
rect 163056 242418 163084 244052
rect 163044 242412 163096 242418
rect 163044 242354 163096 242360
rect 162400 242276 162452 242282
rect 162400 242218 162452 242224
rect 163240 231878 163268 244174
rect 164266 244038 164464 244066
rect 163504 242276 163556 242282
rect 163504 242218 163556 242224
rect 163044 231872 163096 231878
rect 163044 231814 163096 231820
rect 163228 231872 163280 231878
rect 163228 231814 163280 231820
rect 163056 205698 163084 231814
rect 162860 205692 162912 205698
rect 162860 205634 162912 205640
rect 163044 205692 163096 205698
rect 163044 205634 163096 205640
rect 162872 205578 162900 205634
rect 162872 205550 162992 205578
rect 162964 196058 162992 205550
rect 162964 196030 163084 196058
rect 163056 186386 163084 196030
rect 162860 186380 162912 186386
rect 162860 186322 162912 186328
rect 163044 186380 163096 186386
rect 163044 186322 163096 186328
rect 162872 186266 162900 186322
rect 162872 186238 162992 186266
rect 162964 176730 162992 186238
rect 162952 176724 163004 176730
rect 162952 176666 163004 176672
rect 163044 176588 163096 176594
rect 163044 176530 163096 176536
rect 163056 167074 163084 176530
rect 162860 167068 162912 167074
rect 162860 167010 162912 167016
rect 163044 167068 163096 167074
rect 163044 167010 163096 167016
rect 162872 166954 162900 167010
rect 162872 166926 162992 166954
rect 162964 157418 162992 166926
rect 162952 157412 163004 157418
rect 162952 157354 163004 157360
rect 163044 157276 163096 157282
rect 163044 157218 163096 157224
rect 163056 147694 163084 157218
rect 162860 147688 162912 147694
rect 163044 147688 163096 147694
rect 162912 147636 162992 147642
rect 162860 147630 162992 147636
rect 163044 147630 163096 147636
rect 162872 147614 162992 147630
rect 162964 143546 162992 147614
rect 162952 143540 163004 143546
rect 162952 143482 163004 143488
rect 162952 137964 163004 137970
rect 162952 137906 163004 137912
rect 162964 133906 162992 137906
rect 162964 133878 163084 133906
rect 163056 128382 163084 133878
rect 162860 128376 162912 128382
rect 163044 128376 163096 128382
rect 162912 128324 162992 128330
rect 162860 128318 162992 128324
rect 163044 128318 163096 128324
rect 162872 128302 162992 128318
rect 162964 124166 162992 128302
rect 162952 124160 163004 124166
rect 162952 124102 163004 124108
rect 163044 114572 163096 114578
rect 163044 114514 163096 114520
rect 163056 109070 163084 114514
rect 162860 109064 162912 109070
rect 163044 109064 163096 109070
rect 162912 109012 162992 109018
rect 162860 109006 162992 109012
rect 163044 109006 163096 109012
rect 162872 108990 162992 109006
rect 162964 99414 162992 108990
rect 162952 99408 163004 99414
rect 162952 99350 163004 99356
rect 163044 99340 163096 99346
rect 163044 99282 163096 99288
rect 163056 96626 163084 99282
rect 162860 96620 162912 96626
rect 162860 96562 162912 96568
rect 163044 96620 163096 96626
rect 163044 96562 163096 96568
rect 162872 87145 162900 96562
rect 162858 87136 162914 87145
rect 162858 87071 162914 87080
rect 162950 87000 163006 87009
rect 162950 86935 163006 86944
rect 162964 85542 162992 86935
rect 162952 85536 163004 85542
rect 162952 85478 163004 85484
rect 163228 75948 163280 75954
rect 163228 75890 163280 75896
rect 163240 67726 163268 75890
rect 162952 67720 163004 67726
rect 162952 67662 163004 67668
rect 163228 67720 163280 67726
rect 163228 67662 163280 67668
rect 162964 66230 162992 67662
rect 162952 66224 163004 66230
rect 162952 66166 163004 66172
rect 162860 56636 162912 56642
rect 162860 56578 162912 56584
rect 162872 48362 162900 56578
rect 162872 48334 162992 48362
rect 162964 42106 162992 48334
rect 162964 42078 163268 42106
rect 163240 38570 163268 42078
rect 163148 38542 163268 38570
rect 163148 33674 163176 38542
rect 163056 33646 163176 33674
rect 163056 12458 163084 33646
rect 162872 12430 163084 12458
rect 161572 7608 161624 7614
rect 161572 7550 161624 7556
rect 162308 7608 162360 7614
rect 162308 7550 162360 7556
rect 161112 6384 161164 6390
rect 161112 6326 161164 6332
rect 160744 5568 160796 5574
rect 160744 5510 160796 5516
rect 160192 5092 160244 5098
rect 160192 5034 160244 5040
rect 160100 3664 160152 3670
rect 160100 3606 160152 3612
rect 161124 480 161152 6326
rect 162320 480 162348 7550
rect 162872 5166 162900 12430
rect 163516 5642 163544 242218
rect 164332 239352 164384 239358
rect 164332 239294 164384 239300
rect 164240 234796 164292 234802
rect 164240 234738 164292 234744
rect 163504 5636 163556 5642
rect 163504 5578 163556 5584
rect 162860 5160 162912 5166
rect 162860 5102 162912 5108
rect 163504 5092 163556 5098
rect 163504 5034 163556 5040
rect 163516 480 163544 5034
rect 164252 3738 164280 234738
rect 164344 5166 164372 239294
rect 164436 8945 164464 244038
rect 164528 244038 164910 244066
rect 165264 244038 165554 244066
rect 165724 244038 166106 244066
rect 164528 234802 164556 244038
rect 165264 239358 165292 244038
rect 165252 239352 165304 239358
rect 165252 239294 165304 239300
rect 164516 234796 164568 234802
rect 164516 234738 164568 234744
rect 165724 8974 165752 244038
rect 166736 242486 166764 244052
rect 167104 244038 167302 244066
rect 167656 244038 167946 244066
rect 168392 244038 168590 244066
rect 168852 244038 169142 244066
rect 166724 242480 166776 242486
rect 166724 242422 166776 242428
rect 167000 239352 167052 239358
rect 167000 239294 167052 239300
rect 165712 8968 165764 8974
rect 164422 8936 164478 8945
rect 165712 8910 165764 8916
rect 164422 8871 164478 8880
rect 164700 5636 164752 5642
rect 164700 5578 164752 5584
rect 164332 5160 164384 5166
rect 164332 5102 164384 5108
rect 164240 3732 164292 3738
rect 164240 3674 164292 3680
rect 164712 480 164740 5578
rect 167012 3806 167040 239294
rect 167104 5370 167132 244038
rect 167656 239358 167684 244038
rect 167644 239352 167696 239358
rect 167644 239294 167696 239300
rect 168196 5568 168248 5574
rect 168196 5510 168248 5516
rect 167092 5364 167144 5370
rect 167092 5306 167144 5312
rect 167184 5160 167236 5166
rect 167184 5102 167236 5108
rect 167000 3800 167052 3806
rect 167000 3742 167052 3748
rect 165896 3460 165948 3466
rect 165896 3402 165948 3408
rect 165908 480 165936 3402
rect 167196 1442 167224 5102
rect 167104 1414 167224 1442
rect 167104 480 167132 1414
rect 168208 480 168236 5510
rect 168392 3874 168420 244038
rect 168852 239306 168880 244038
rect 169772 242894 169800 244052
rect 169760 242888 169812 242894
rect 169760 242830 169812 242836
rect 170416 242554 170444 244052
rect 170692 244038 170982 244066
rect 171244 244038 171626 244066
rect 171888 244038 172270 244066
rect 172624 244038 172822 244066
rect 170404 242548 170456 242554
rect 170404 242490 170456 242496
rect 170692 239306 170720 244038
rect 168668 239278 168880 239306
rect 169956 239278 170720 239306
rect 171140 239352 171192 239358
rect 171140 239294 171192 239300
rect 168668 225078 168696 239278
rect 169956 227050 169984 239278
rect 169944 227044 169996 227050
rect 169944 226986 169996 226992
rect 168656 225072 168708 225078
rect 168656 225014 168708 225020
rect 168564 224936 168616 224942
rect 168564 224878 168616 224884
rect 168576 222154 168604 224878
rect 170048 222222 170076 222253
rect 170036 222216 170088 222222
rect 170088 222164 170168 222170
rect 170036 222158 170168 222164
rect 168564 222148 168616 222154
rect 170048 222142 170168 222158
rect 168564 222090 168616 222096
rect 168656 222012 168708 222018
rect 168656 221954 168708 221960
rect 168668 205578 168696 221954
rect 170140 212566 170168 222142
rect 170036 212560 170088 212566
rect 170036 212502 170088 212508
rect 170128 212560 170180 212566
rect 170128 212502 170180 212508
rect 170048 205578 170076 212502
rect 168576 205550 168696 205578
rect 169956 205550 170076 205578
rect 168576 202881 168604 205550
rect 169956 202881 169984 205550
rect 168562 202872 168618 202881
rect 168562 202807 168618 202816
rect 168838 202872 168894 202881
rect 168838 202807 168894 202816
rect 169758 202872 169814 202881
rect 169758 202807 169814 202816
rect 169942 202872 169998 202881
rect 169942 202807 169998 202816
rect 168852 193254 168880 202807
rect 169772 193254 169800 202807
rect 168656 193248 168708 193254
rect 168656 193190 168708 193196
rect 168840 193248 168892 193254
rect 168840 193190 168892 193196
rect 169760 193248 169812 193254
rect 169760 193190 169812 193196
rect 170036 193248 170088 193254
rect 170036 193190 170088 193196
rect 168668 186266 168696 193190
rect 170048 186266 170076 193190
rect 168576 186238 168696 186266
rect 169956 186238 170076 186266
rect 168576 183569 168604 186238
rect 169956 183569 169984 186238
rect 168562 183560 168618 183569
rect 168562 183495 168618 183504
rect 168838 183560 168894 183569
rect 168838 183495 168894 183504
rect 169758 183560 169814 183569
rect 169758 183495 169814 183504
rect 169942 183560 169998 183569
rect 169942 183495 169998 183504
rect 168852 173942 168880 183495
rect 169772 173942 169800 183495
rect 168656 173936 168708 173942
rect 168656 173878 168708 173884
rect 168840 173936 168892 173942
rect 168840 173878 168892 173884
rect 169760 173936 169812 173942
rect 169760 173878 169812 173884
rect 170036 173936 170088 173942
rect 170036 173878 170088 173884
rect 168668 166954 168696 173878
rect 170048 166954 170076 173878
rect 168576 166926 168696 166954
rect 169956 166926 170076 166954
rect 168576 159338 168604 166926
rect 169956 164218 169984 166926
rect 169944 164212 169996 164218
rect 169944 164154 169996 164160
rect 170036 164212 170088 164218
rect 170036 164154 170088 164160
rect 168576 159310 168788 159338
rect 168760 154578 168788 159310
rect 168668 154550 168788 154578
rect 168668 148322 168696 154550
rect 168484 148294 168696 148322
rect 168484 143585 168512 148294
rect 170048 147642 170076 164154
rect 169956 147614 170076 147642
rect 169956 144888 169984 147614
rect 169772 144860 169984 144888
rect 168470 143576 168526 143585
rect 168470 143511 168526 143520
rect 168838 143576 168894 143585
rect 168838 143511 168894 143520
rect 168852 134858 168880 143511
rect 169772 135289 169800 144860
rect 169758 135280 169814 135289
rect 169758 135215 169814 135224
rect 170034 135280 170090 135289
rect 170034 135215 170090 135224
rect 168760 134830 168880 134858
rect 168760 134026 168788 134830
rect 168748 134020 168800 134026
rect 168748 133962 168800 133968
rect 168840 134020 168892 134026
rect 168840 133962 168892 133968
rect 168852 133890 168880 133962
rect 168840 133884 168892 133890
rect 168840 133826 168892 133832
rect 170048 128330 170076 135215
rect 169956 128302 170076 128330
rect 169956 125576 169984 128302
rect 169772 125548 169984 125576
rect 168840 124228 168892 124234
rect 168840 124170 168892 124176
rect 168852 115870 168880 124170
rect 169772 115977 169800 125548
rect 169758 115968 169814 115977
rect 169758 115903 169814 115912
rect 170034 115968 170090 115977
rect 170034 115903 170090 115912
rect 168840 115864 168892 115870
rect 168840 115806 168892 115812
rect 168748 115796 168800 115802
rect 168748 115738 168800 115744
rect 168760 114594 168788 115738
rect 168760 114566 168880 114594
rect 168852 114510 168880 114566
rect 168840 114504 168892 114510
rect 168840 114446 168892 114452
rect 170048 109018 170076 115903
rect 169956 108990 170076 109018
rect 168840 106276 168892 106282
rect 169956 106264 169984 108990
rect 168840 106218 168892 106224
rect 169772 106236 169984 106264
rect 168852 104854 168880 106218
rect 168840 104848 168892 104854
rect 168840 104790 168892 104796
rect 169772 96665 169800 106236
rect 169758 96656 169814 96665
rect 169758 96591 169814 96600
rect 170034 96656 170090 96665
rect 170034 96591 170090 96600
rect 168840 95260 168892 95266
rect 168840 95202 168892 95208
rect 168852 91798 168880 95202
rect 168472 91792 168524 91798
rect 168472 91734 168524 91740
rect 168840 91792 168892 91798
rect 168840 91734 168892 91740
rect 168484 77382 168512 91734
rect 170048 89706 170076 96591
rect 169864 89678 170076 89706
rect 169864 86970 169892 89678
rect 169852 86964 169904 86970
rect 169852 86906 169904 86912
rect 168472 77376 168524 77382
rect 168472 77318 168524 77324
rect 168656 77376 168708 77382
rect 168656 77318 168708 77324
rect 168668 67833 168696 77318
rect 169760 77308 169812 77314
rect 169760 77250 169812 77256
rect 169772 70258 169800 77250
rect 169772 70230 169892 70258
rect 168654 67824 168710 67833
rect 168654 67759 168710 67768
rect 168562 67654 168618 67663
rect 168562 67589 168618 67598
rect 168576 66230 168604 67589
rect 168564 66224 168616 66230
rect 168564 66166 168616 66172
rect 169864 60722 169892 70230
rect 169852 60716 169904 60722
rect 169852 60658 169904 60664
rect 170036 60716 170088 60722
rect 170036 60658 170088 60664
rect 168472 56636 168524 56642
rect 168472 56578 168524 56584
rect 168484 50946 168512 56578
rect 168484 50918 168604 50946
rect 168576 46918 168604 50918
rect 170048 48328 170076 60658
rect 169864 48300 170076 48328
rect 169864 46918 169892 48300
rect 168564 46912 168616 46918
rect 168564 46854 168616 46860
rect 169852 46912 169904 46918
rect 169852 46854 169904 46860
rect 168656 37324 168708 37330
rect 168656 37266 168708 37272
rect 169944 37324 169996 37330
rect 169944 37266 169996 37272
rect 168668 31822 168696 37266
rect 169956 31822 169984 37266
rect 168656 31816 168708 31822
rect 168656 31758 168708 31764
rect 169944 31816 169996 31822
rect 169944 31758 169996 31764
rect 168748 31680 168800 31686
rect 168748 31622 168800 31628
rect 169944 31680 169996 31686
rect 169944 31622 169996 31628
rect 168760 27606 168788 31622
rect 168564 27600 168616 27606
rect 168564 27542 168616 27548
rect 168748 27600 168800 27606
rect 168748 27542 168800 27548
rect 169956 27554 169984 31622
rect 168576 12510 168604 27542
rect 169956 27526 170168 27554
rect 168564 12504 168616 12510
rect 168564 12446 168616 12452
rect 168472 12436 168524 12442
rect 168472 12378 168524 12384
rect 168484 6225 168512 12378
rect 170140 9722 170168 27526
rect 169852 9716 169904 9722
rect 169852 9658 169904 9664
rect 170128 9716 170180 9722
rect 170128 9658 170180 9664
rect 169864 6458 169892 9658
rect 169852 6452 169904 6458
rect 169852 6394 169904 6400
rect 168470 6216 168526 6225
rect 168470 6151 168526 6160
rect 170588 5228 170640 5234
rect 170588 5170 170640 5176
rect 168380 3868 168432 3874
rect 168380 3810 168432 3816
rect 169392 3528 169444 3534
rect 169392 3470 169444 3476
rect 169404 480 169432 3470
rect 170600 480 170628 5170
rect 171152 4010 171180 239294
rect 171140 4004 171192 4010
rect 171140 3946 171192 3952
rect 171244 3942 171272 244038
rect 171888 239358 171916 244038
rect 171876 239352 171928 239358
rect 171876 239294 171928 239300
rect 171784 6452 171836 6458
rect 171784 6394 171836 6400
rect 171232 3936 171284 3942
rect 171232 3878 171284 3884
rect 171796 480 171824 6394
rect 172624 6361 172652 244038
rect 173452 242010 173480 244052
rect 173440 242004 173492 242010
rect 173440 241946 173492 241952
rect 174096 241670 174124 244052
rect 174372 244038 174662 244066
rect 175306 244038 175412 244066
rect 174084 241664 174136 241670
rect 174084 241606 174136 241612
rect 174372 231878 174400 244038
rect 174544 241664 174596 241670
rect 174544 241606 174596 241612
rect 174084 231872 174136 231878
rect 174084 231814 174136 231820
rect 174360 231872 174412 231878
rect 174360 231814 174412 231820
rect 174096 205698 174124 231814
rect 173900 205692 173952 205698
rect 173900 205634 173952 205640
rect 174084 205692 174136 205698
rect 174084 205634 174136 205640
rect 173912 205578 173940 205634
rect 173912 205550 174032 205578
rect 174004 196058 174032 205550
rect 174004 196030 174124 196058
rect 174096 186386 174124 196030
rect 173900 186380 173952 186386
rect 173900 186322 173952 186328
rect 174084 186380 174136 186386
rect 174084 186322 174136 186328
rect 173912 186266 173940 186322
rect 173912 186238 174032 186266
rect 174004 183569 174032 186238
rect 173990 183560 174046 183569
rect 173990 183495 174046 183504
rect 174266 183560 174322 183569
rect 174266 183495 174322 183504
rect 174280 173942 174308 183495
rect 174084 173936 174136 173942
rect 174084 173878 174136 173884
rect 174268 173936 174320 173942
rect 174268 173878 174320 173884
rect 174096 167074 174124 173878
rect 173900 167068 173952 167074
rect 173900 167010 173952 167016
rect 174084 167068 174136 167074
rect 174084 167010 174136 167016
rect 173912 166954 173940 167010
rect 173912 166926 174032 166954
rect 174004 164218 174032 166926
rect 173992 164212 174044 164218
rect 173992 164154 174044 164160
rect 173992 157344 174044 157350
rect 173992 157286 174044 157292
rect 174004 154578 174032 157286
rect 174004 154550 174124 154578
rect 174096 147694 174124 154550
rect 173900 147688 173952 147694
rect 174084 147688 174136 147694
rect 173952 147636 174032 147642
rect 173900 147630 174032 147636
rect 174084 147630 174136 147636
rect 173912 147614 174032 147630
rect 174004 144906 174032 147614
rect 173992 144900 174044 144906
rect 173992 144842 174044 144848
rect 173992 137964 174044 137970
rect 173992 137906 174044 137912
rect 174004 135266 174032 137906
rect 174004 135238 174124 135266
rect 174096 128382 174124 135238
rect 173900 128376 173952 128382
rect 174084 128376 174136 128382
rect 173952 128324 174032 128330
rect 173900 128318 174032 128324
rect 174084 128318 174136 128324
rect 173912 128302 174032 128318
rect 174004 125594 174032 128302
rect 173992 125588 174044 125594
rect 173992 125530 174044 125536
rect 173992 118652 174044 118658
rect 173992 118594 174044 118600
rect 174004 115954 174032 118594
rect 174004 115926 174124 115954
rect 174096 109070 174124 115926
rect 173900 109064 173952 109070
rect 174084 109064 174136 109070
rect 173952 109012 174032 109018
rect 173900 109006 174032 109012
rect 174084 109006 174136 109012
rect 173912 108990 174032 109006
rect 174004 106282 174032 108990
rect 173992 106276 174044 106282
rect 173992 106218 174044 106224
rect 173992 99340 174044 99346
rect 173992 99282 174044 99288
rect 174004 96642 174032 99282
rect 174004 96614 174124 96642
rect 174096 89758 174124 96614
rect 173900 89752 173952 89758
rect 174084 89752 174136 89758
rect 173952 89700 174032 89706
rect 173900 89694 174032 89700
rect 174084 89694 174136 89700
rect 173912 89678 174032 89694
rect 174004 86970 174032 89678
rect 173992 86964 174044 86970
rect 173992 86906 174044 86912
rect 174084 77308 174136 77314
rect 174084 77250 174136 77256
rect 174096 67658 174124 77250
rect 173992 67652 174044 67658
rect 173992 67594 174044 67600
rect 174084 67652 174136 67658
rect 174084 67594 174136 67600
rect 174004 60738 174032 67594
rect 174004 60710 174124 60738
rect 174096 57934 174124 60710
rect 174084 57928 174136 57934
rect 174084 57870 174136 57876
rect 173992 48340 174044 48346
rect 173992 48282 174044 48288
rect 174004 41426 174032 48282
rect 174004 41398 174124 41426
rect 174096 33862 174124 41398
rect 174084 33856 174136 33862
rect 174084 33798 174136 33804
rect 173992 29028 174044 29034
rect 173992 28970 174044 28976
rect 174004 27606 174032 28970
rect 173992 27600 174044 27606
rect 173992 27542 174044 27548
rect 173992 22092 174044 22098
rect 173992 22034 174044 22040
rect 173900 16720 173952 16726
rect 173898 16688 173900 16697
rect 173952 16688 173954 16697
rect 173898 16623 173954 16632
rect 172610 6352 172666 6361
rect 172610 6287 172666 6296
rect 174004 5438 174032 22034
rect 173992 5432 174044 5438
rect 173992 5374 174044 5380
rect 174176 5432 174228 5438
rect 174176 5374 174228 5380
rect 172980 3664 173032 3670
rect 172980 3606 173032 3612
rect 172992 480 173020 3606
rect 174188 480 174216 5374
rect 174556 4078 174584 241606
rect 175384 6610 175412 244038
rect 175844 242078 175872 244052
rect 176028 244038 176502 244066
rect 176764 244038 177146 244066
rect 175832 242072 175884 242078
rect 175832 242014 175884 242020
rect 176028 239306 176056 244038
rect 176108 242480 176160 242486
rect 176108 242422 176160 242428
rect 175292 6582 175412 6610
rect 175476 239278 176056 239306
rect 175292 6526 175320 6582
rect 175280 6520 175332 6526
rect 175280 6462 175332 6468
rect 175372 6520 175424 6526
rect 175372 6462 175424 6468
rect 174544 4072 174596 4078
rect 174544 4014 174596 4020
rect 175384 480 175412 6462
rect 175476 5506 175504 239278
rect 176120 238490 176148 242422
rect 175936 238462 176148 238490
rect 175464 5500 175516 5506
rect 175464 5442 175516 5448
rect 175936 4146 175964 238462
rect 176382 40352 176438 40361
rect 176566 40352 176622 40361
rect 176438 40310 176566 40338
rect 176382 40287 176438 40296
rect 176566 40287 176622 40296
rect 176764 6594 176792 244038
rect 177304 242004 177356 242010
rect 177304 241946 177356 241952
rect 176752 6588 176804 6594
rect 176752 6530 176804 6536
rect 175924 4140 175976 4146
rect 175924 4082 175976 4088
rect 176568 3800 176620 3806
rect 176568 3742 176620 3748
rect 176580 480 176608 3742
rect 177316 3398 177344 241946
rect 177684 241670 177712 244052
rect 178052 244038 178342 244066
rect 177672 241664 177724 241670
rect 177672 241606 177724 241612
rect 177948 62824 178000 62830
rect 177948 62766 178000 62772
rect 177960 58041 177988 62766
rect 177946 58032 178002 58041
rect 177946 57967 178002 57976
rect 178052 4758 178080 244038
rect 178512 239306 178540 244174
rect 179524 241874 179552 244052
rect 179512 241868 179564 241874
rect 179512 241810 179564 241816
rect 179708 241505 179736 244174
rect 180826 244038 180932 244066
rect 180064 242548 180116 242554
rect 180064 242490 180116 242496
rect 179694 241496 179750 241505
rect 179694 241431 179750 241440
rect 179878 241496 179934 241505
rect 179878 241431 179934 241440
rect 178236 239278 178540 239306
rect 178236 215286 178264 239278
rect 179892 231878 179920 241431
rect 179604 231872 179656 231878
rect 179602 231840 179604 231849
rect 179880 231872 179932 231878
rect 179656 231840 179658 231849
rect 179602 231775 179658 231784
rect 179786 231840 179842 231849
rect 179880 231814 179932 231820
rect 179786 231775 179842 231784
rect 179800 222222 179828 231775
rect 179604 222216 179656 222222
rect 179604 222158 179656 222164
rect 179788 222216 179840 222222
rect 179788 222158 179840 222164
rect 179616 215422 179644 222158
rect 179604 215416 179656 215422
rect 179604 215358 179656 215364
rect 178224 215280 178276 215286
rect 178224 215222 178276 215228
rect 178224 212560 178276 212566
rect 178224 212502 178276 212508
rect 179512 212560 179564 212566
rect 179512 212502 179564 212508
rect 178236 202881 178264 212502
rect 179524 205714 179552 212502
rect 179432 205686 179552 205714
rect 179432 205578 179460 205686
rect 179432 205550 179552 205578
rect 178222 202872 178278 202881
rect 178222 202807 178278 202816
rect 178406 202872 178462 202881
rect 178406 202807 178462 202816
rect 178420 193254 178448 202807
rect 178224 193248 178276 193254
rect 178224 193190 178276 193196
rect 178408 193248 178460 193254
rect 178408 193190 178460 193196
rect 178236 183569 178264 193190
rect 179524 186402 179552 205550
rect 179432 186374 179552 186402
rect 179432 186266 179460 186374
rect 179432 186238 179552 186266
rect 178222 183560 178278 183569
rect 178222 183495 178278 183504
rect 178406 183560 178462 183569
rect 178406 183495 178462 183504
rect 178420 173942 178448 183495
rect 178224 173936 178276 173942
rect 178224 173878 178276 173884
rect 178408 173936 178460 173942
rect 178408 173878 178460 173884
rect 178236 164218 178264 173878
rect 179524 167090 179552 186238
rect 179432 167062 179552 167090
rect 179432 166954 179460 167062
rect 179432 166926 179552 166954
rect 178224 164212 178276 164218
rect 178224 164154 178276 164160
rect 178408 164212 178460 164218
rect 178408 164154 178460 164160
rect 178420 154601 178448 164154
rect 178222 154592 178278 154601
rect 178222 154527 178278 154536
rect 178406 154592 178462 154601
rect 178406 154527 178462 154536
rect 178236 144906 178264 154527
rect 179524 147778 179552 166926
rect 179432 147750 179552 147778
rect 179432 147642 179460 147750
rect 179432 147614 179552 147642
rect 178224 144900 178276 144906
rect 178224 144842 178276 144848
rect 178408 144900 178460 144906
rect 178408 144842 178460 144848
rect 178420 135289 178448 144842
rect 178222 135280 178278 135289
rect 178222 135215 178278 135224
rect 178406 135280 178462 135289
rect 178406 135215 178462 135224
rect 178236 125594 178264 135215
rect 179524 128466 179552 147614
rect 179432 128438 179552 128466
rect 179432 128330 179460 128438
rect 179432 128302 179552 128330
rect 178224 125588 178276 125594
rect 178224 125530 178276 125536
rect 178224 116000 178276 116006
rect 178224 115942 178276 115948
rect 178236 106282 178264 115942
rect 179524 109154 179552 128302
rect 179432 109126 179552 109154
rect 179432 109018 179460 109126
rect 179432 108990 179552 109018
rect 178224 106276 178276 106282
rect 178224 106218 178276 106224
rect 178224 96688 178276 96694
rect 178224 96630 178276 96636
rect 178236 86970 178264 96630
rect 179524 89842 179552 108990
rect 179432 89814 179552 89842
rect 179432 89706 179460 89814
rect 179432 89678 179552 89706
rect 178224 86964 178276 86970
rect 178224 86906 178276 86912
rect 178224 77308 178276 77314
rect 178224 77250 178276 77256
rect 178236 62830 178264 77250
rect 179524 70394 179552 89678
rect 179432 70366 179552 70394
rect 179432 70258 179460 70366
rect 179432 70230 179552 70258
rect 178224 62824 178276 62830
rect 178224 62766 178276 62772
rect 178130 58032 178186 58041
rect 178186 57990 178264 58018
rect 178130 57967 178186 57976
rect 178236 57934 178264 57990
rect 178224 57928 178276 57934
rect 178224 57870 178276 57876
rect 179524 51202 179552 70230
rect 179512 51196 179564 51202
rect 179512 51138 179564 51144
rect 179512 51060 179564 51066
rect 179512 51002 179564 51008
rect 178316 48340 178368 48346
rect 178316 48282 178368 48288
rect 178328 41426 178356 48282
rect 178144 41410 178356 41426
rect 179524 41426 179552 51002
rect 178132 41404 178368 41410
rect 178184 41398 178316 41404
rect 178132 41346 178184 41352
rect 179524 41398 179644 41426
rect 178316 41346 178368 41352
rect 178328 31278 178356 41346
rect 178316 31272 178368 31278
rect 178316 31214 178368 31220
rect 178316 31136 178368 31142
rect 178316 31078 178368 31084
rect 178328 22250 178356 31078
rect 179616 29102 179644 41398
rect 179604 29096 179656 29102
rect 179604 29038 179656 29044
rect 179512 29028 179564 29034
rect 179512 28970 179564 28976
rect 179524 27606 179552 28970
rect 179512 27600 179564 27606
rect 179512 27542 179564 27548
rect 178236 22222 178356 22250
rect 178236 22114 178264 22222
rect 178144 22086 178264 22114
rect 178144 21978 178172 22086
rect 178144 21950 178264 21978
rect 178236 6662 178264 21950
rect 179512 18012 179564 18018
rect 179512 17954 179564 17960
rect 178224 6656 178276 6662
rect 178224 6598 178276 6604
rect 178960 6588 179012 6594
rect 178960 6530 179012 6536
rect 178682 5400 178738 5409
rect 178682 5335 178738 5344
rect 178696 5302 178724 5335
rect 178684 5296 178736 5302
rect 178684 5238 178736 5244
rect 178040 4752 178092 4758
rect 178040 4694 178092 4700
rect 177764 3936 177816 3942
rect 177764 3878 177816 3884
rect 177304 3392 177356 3398
rect 177304 3334 177356 3340
rect 177776 480 177804 3878
rect 178972 480 179000 6530
rect 179524 4690 179552 17954
rect 179512 4684 179564 4690
rect 179512 4626 179564 4632
rect 180076 3330 180104 242490
rect 180904 6730 180932 244038
rect 181364 242486 181392 244052
rect 181548 244038 182022 244066
rect 182284 244038 182666 244066
rect 181352 242480 181404 242486
rect 181352 242422 181404 242428
rect 181548 239306 181576 244038
rect 181628 242208 181680 242214
rect 181628 242150 181680 242156
rect 180996 239278 181576 239306
rect 180892 6724 180944 6730
rect 180892 6666 180944 6672
rect 180996 4554 181024 239278
rect 181640 238354 181668 242150
rect 181456 238326 181668 238354
rect 180984 4548 181036 4554
rect 180984 4490 181036 4496
rect 180156 3868 180208 3874
rect 180156 3810 180208 3816
rect 180064 3324 180116 3330
rect 180064 3266 180116 3272
rect 180168 480 180196 3810
rect 181456 3262 181484 238326
rect 182284 6798 182312 244038
rect 183204 241602 183232 244052
rect 183572 244038 183862 244066
rect 184124 244038 184414 244066
rect 183376 242820 183428 242826
rect 183376 242762 183428 242768
rect 183388 242706 183416 242762
rect 183388 242690 183508 242706
rect 183388 242684 183520 242690
rect 183388 242678 183468 242684
rect 183468 242626 183520 242632
rect 183192 241596 183244 241602
rect 183192 241538 183244 241544
rect 183468 16720 183520 16726
rect 183466 16688 183468 16697
rect 183520 16688 183522 16697
rect 183466 16623 183522 16632
rect 182272 6792 182324 6798
rect 182272 6734 182324 6740
rect 183468 5500 183520 5506
rect 183468 5442 183520 5448
rect 181536 5432 181588 5438
rect 183480 5409 183508 5442
rect 181536 5374 181588 5380
rect 183466 5400 183522 5409
rect 181444 3256 181496 3262
rect 181444 3198 181496 3204
rect 181548 2802 181576 5374
rect 183466 5335 183522 5344
rect 183572 4622 183600 244038
rect 184124 239306 184152 244038
rect 184204 242480 184256 242486
rect 184204 242422 184256 242428
rect 183756 239278 184152 239306
rect 183756 176610 183784 239278
rect 183664 176582 183784 176610
rect 183664 176338 183692 176582
rect 183664 176310 183784 176338
rect 183756 157434 183784 176310
rect 183664 157406 183784 157434
rect 183664 157298 183692 157406
rect 183664 157270 183784 157298
rect 183756 138122 183784 157270
rect 183664 138094 183784 138122
rect 183664 137714 183692 138094
rect 183664 137686 183784 137714
rect 183756 118810 183784 137686
rect 183664 118782 183784 118810
rect 183664 118674 183692 118782
rect 183664 118646 183784 118674
rect 183756 60738 183784 118646
rect 183664 60710 183784 60738
rect 183664 60602 183692 60710
rect 183664 60574 183784 60602
rect 183756 22114 183784 60574
rect 183664 22086 183784 22114
rect 183664 21978 183692 22086
rect 183664 21950 183784 21978
rect 183756 6866 183784 21950
rect 183744 6860 183796 6866
rect 183744 6802 183796 6808
rect 183560 4616 183612 4622
rect 183560 4558 183612 4564
rect 182548 3936 182600 3942
rect 182548 3878 182600 3884
rect 181364 2774 181576 2802
rect 181364 480 181392 2774
rect 182560 480 182588 3878
rect 183744 3392 183796 3398
rect 183744 3334 183796 3340
rect 183756 480 183784 3334
rect 184216 3194 184244 242422
rect 185044 242010 185072 244052
rect 185032 242004 185084 242010
rect 185032 241946 185084 241952
rect 185228 241505 185256 244174
rect 185872 244038 186254 244066
rect 185584 242344 185636 242350
rect 185584 242286 185636 242292
rect 185214 241496 185270 241505
rect 185214 241431 185270 241440
rect 185398 241496 185454 241505
rect 185398 241431 185454 241440
rect 185032 231940 185084 231946
rect 185032 231882 185084 231888
rect 185044 7585 185072 231882
rect 185412 231878 185440 241431
rect 185124 231872 185176 231878
rect 185122 231840 185124 231849
rect 185400 231872 185452 231878
rect 185176 231840 185178 231849
rect 185122 231775 185178 231784
rect 185306 231840 185362 231849
rect 185400 231814 185452 231820
rect 185306 231775 185362 231784
rect 185320 222222 185348 231775
rect 185124 222216 185176 222222
rect 185124 222158 185176 222164
rect 185308 222216 185360 222222
rect 185308 222158 185360 222164
rect 185136 212566 185164 222158
rect 185124 212560 185176 212566
rect 185124 212502 185176 212508
rect 185216 212560 185268 212566
rect 185216 212502 185268 212508
rect 185228 176610 185256 212502
rect 185136 176582 185256 176610
rect 185136 176338 185164 176582
rect 185136 176310 185256 176338
rect 185228 157434 185256 176310
rect 185136 157406 185256 157434
rect 185136 157298 185164 157406
rect 185136 157270 185256 157298
rect 185228 138122 185256 157270
rect 185136 138094 185256 138122
rect 185136 137714 185164 138094
rect 185136 137686 185256 137714
rect 185228 118810 185256 137686
rect 185136 118782 185256 118810
rect 185136 118674 185164 118782
rect 185136 118646 185256 118674
rect 185228 60738 185256 118646
rect 185136 60710 185256 60738
rect 185136 60602 185164 60710
rect 185136 60574 185256 60602
rect 185228 22114 185256 60574
rect 185136 22086 185256 22114
rect 185136 21978 185164 22086
rect 185136 21950 185256 21978
rect 185030 7576 185086 7585
rect 185030 7511 185086 7520
rect 184848 4684 184900 4690
rect 184848 4626 184900 4632
rect 184204 3188 184256 3194
rect 184204 3130 184256 3136
rect 184860 480 184888 4626
rect 185228 4486 185256 21950
rect 185216 4480 185268 4486
rect 185216 4422 185268 4428
rect 185596 3126 185624 242286
rect 185872 231946 185900 244038
rect 186884 243030 186912 244052
rect 187068 244038 187542 244066
rect 187804 244038 188094 244066
rect 186872 243024 186924 243030
rect 186872 242966 186924 242972
rect 187068 239306 187096 244038
rect 187148 242412 187200 242418
rect 187148 242354 187200 242360
rect 186424 239278 187096 239306
rect 185860 231940 185912 231946
rect 185860 231882 185912 231888
rect 186424 4418 186452 239278
rect 187160 238490 187188 242354
rect 186976 238462 187188 238490
rect 186412 4412 186464 4418
rect 186412 4354 186464 4360
rect 186044 4004 186096 4010
rect 186044 3946 186096 3952
rect 185584 3120 185636 3126
rect 185584 3062 185636 3068
rect 186056 480 186084 3946
rect 186976 3058 187004 238462
rect 187804 9042 187832 244038
rect 188344 242684 188396 242690
rect 188344 242626 188396 242632
rect 187792 9036 187844 9042
rect 187792 8978 187844 8984
rect 187240 5500 187292 5506
rect 187240 5442 187292 5448
rect 186964 3052 187016 3058
rect 186964 2994 187016 3000
rect 187252 480 187280 5442
rect 188356 2922 188384 242626
rect 188724 242554 188752 244052
rect 189092 244038 189382 244066
rect 189644 244038 189934 244066
rect 188712 242548 188764 242554
rect 188712 242490 188764 242496
rect 188436 241868 188488 241874
rect 188436 241810 188488 241816
rect 188448 4842 188476 241810
rect 188986 95296 189042 95305
rect 188986 95231 189042 95240
rect 189000 95198 189028 95231
rect 188988 95192 189040 95198
rect 188988 95134 189040 95140
rect 189092 87038 189120 244038
rect 189644 239306 189672 244038
rect 190564 242894 190592 244052
rect 190552 242888 190604 242894
rect 190552 242830 190604 242836
rect 189276 239278 189672 239306
rect 190552 239352 190604 239358
rect 190552 239294 190604 239300
rect 189276 157434 189304 239278
rect 190458 212528 190514 212537
rect 190458 212463 190514 212472
rect 190472 202910 190500 212463
rect 190460 202904 190512 202910
rect 190458 202872 190460 202881
rect 190512 202872 190514 202881
rect 190458 202807 190514 202816
rect 190472 193254 190500 202807
rect 190460 193248 190512 193254
rect 190460 193190 190512 193196
rect 190460 162852 190512 162858
rect 190460 162794 190512 162800
rect 189184 157406 189304 157434
rect 189184 157298 189212 157406
rect 189184 157270 189304 157298
rect 189276 145081 189304 157270
rect 190472 153241 190500 162794
rect 190458 153232 190514 153241
rect 190458 153167 190514 153176
rect 189262 145072 189318 145081
rect 189262 145007 189318 145016
rect 189262 144936 189318 144945
rect 189262 144871 189318 144880
rect 189276 143546 189304 144871
rect 189264 143540 189316 143546
rect 189264 143482 189316 143488
rect 190368 143540 190420 143546
rect 190368 143482 190420 143488
rect 189264 133952 189316 133958
rect 190380 133929 190408 143482
rect 189264 133894 189316 133900
rect 190366 133920 190422 133929
rect 189276 125769 189304 133894
rect 190366 133855 190422 133864
rect 190460 133884 190512 133890
rect 190460 133826 190512 133832
rect 189262 125760 189318 125769
rect 189262 125695 189318 125704
rect 189262 125624 189318 125633
rect 189262 125559 189318 125568
rect 189276 124166 189304 125559
rect 190472 124273 190500 133826
rect 190458 124264 190514 124273
rect 190458 124199 190514 124208
rect 189264 124160 189316 124166
rect 189264 124102 189316 124108
rect 189264 114572 189316 114578
rect 189264 114514 189316 114520
rect 189276 104922 189304 114514
rect 189172 104916 189224 104922
rect 189172 104858 189224 104864
rect 189264 104916 189316 104922
rect 189264 104858 189316 104864
rect 189184 104825 189212 104858
rect 189170 104816 189226 104825
rect 189170 104751 189226 104760
rect 189080 87032 189132 87038
rect 189080 86974 189132 86980
rect 189080 86896 189132 86902
rect 189080 86838 189132 86844
rect 188448 4814 188660 4842
rect 188436 4752 188488 4758
rect 188436 4694 188488 4700
rect 188344 2916 188396 2922
rect 188344 2858 188396 2864
rect 188448 480 188476 4694
rect 188632 2990 188660 4814
rect 189092 4350 189120 86838
rect 189172 85604 189224 85610
rect 189172 85546 189224 85552
rect 189184 85513 189212 85546
rect 189170 85504 189226 85513
rect 189170 85439 189226 85448
rect 189262 85368 189318 85377
rect 189262 85303 189318 85312
rect 189276 66212 189304 85303
rect 189184 66184 189304 66212
rect 189184 64870 189212 66184
rect 189172 64864 189224 64870
rect 189172 64806 189224 64812
rect 189356 46980 189408 46986
rect 189356 46922 189408 46928
rect 189368 38690 189396 46922
rect 189264 38684 189316 38690
rect 189264 38626 189316 38632
rect 189356 38684 189408 38690
rect 189356 38626 189408 38632
rect 189276 27849 189304 38626
rect 189262 27840 189318 27849
rect 189262 27775 189318 27784
rect 189170 27704 189226 27713
rect 189170 27639 189226 27648
rect 189184 26246 189212 27639
rect 189172 26240 189224 26246
rect 189172 26182 189224 26188
rect 189172 16652 189224 16658
rect 189172 16594 189224 16600
rect 189184 9110 189212 16594
rect 190460 13524 190512 13530
rect 190460 13466 190512 13472
rect 189172 9104 189224 9110
rect 189172 9046 189224 9052
rect 189080 4344 189132 4350
rect 189080 4286 189132 4292
rect 190472 4282 190500 13466
rect 190564 9178 190592 239294
rect 190748 231878 190776 244174
rect 191392 244038 191774 244066
rect 191104 241664 191156 241670
rect 191104 241606 191156 241612
rect 190644 231872 190696 231878
rect 190644 231814 190696 231820
rect 190736 231872 190788 231878
rect 190736 231814 190788 231820
rect 190656 224890 190684 231814
rect 190656 224862 190776 224890
rect 190748 222193 190776 224862
rect 190734 222184 190790 222193
rect 190734 222119 190790 222128
rect 190918 222184 190974 222193
rect 190918 222119 190974 222128
rect 190932 212566 190960 222119
rect 190736 212560 190788 212566
rect 190734 212528 190736 212537
rect 190920 212560 190972 212566
rect 190788 212528 190790 212537
rect 190920 212502 190972 212508
rect 190734 212463 190790 212472
rect 190644 202904 190696 202910
rect 190642 202872 190644 202881
rect 190696 202872 190698 202881
rect 190642 202807 190698 202816
rect 190736 193248 190788 193254
rect 190734 193216 190736 193225
rect 190788 193216 190790 193225
rect 190734 193151 190790 193160
rect 190918 193216 190974 193225
rect 190918 193151 190974 193160
rect 190932 186130 190960 193151
rect 190748 186102 190960 186130
rect 190748 183530 190776 186102
rect 190736 183524 190788 183530
rect 190736 183466 190788 183472
rect 190736 173936 190788 173942
rect 190736 173878 190788 173884
rect 190748 169130 190776 173878
rect 190656 169102 190776 169130
rect 190656 162858 190684 169102
rect 190644 162852 190696 162858
rect 190644 162794 190696 162800
rect 190734 153232 190790 153241
rect 190734 153167 190790 153176
rect 190748 144922 190776 153167
rect 190656 144906 190776 144922
rect 190644 144900 190776 144906
rect 190696 144894 190776 144900
rect 190644 144842 190696 144848
rect 190736 144832 190788 144838
rect 190736 144774 190788 144780
rect 190748 143546 190776 144774
rect 190736 143540 190788 143546
rect 190736 143482 190788 143488
rect 190642 133920 190698 133929
rect 190642 133855 190644 133864
rect 190696 133855 190698 133864
rect 190644 133826 190696 133832
rect 190642 124264 190698 124273
rect 190642 124199 190698 124208
rect 190656 124166 190684 124199
rect 190644 124160 190696 124166
rect 190644 124102 190696 124108
rect 190920 124092 190972 124098
rect 190920 124034 190972 124040
rect 190932 115818 190960 124034
rect 190840 115790 190960 115818
rect 190840 106321 190868 115790
rect 190642 106312 190698 106321
rect 190642 106247 190644 106256
rect 190696 106247 190698 106256
rect 190826 106312 190882 106321
rect 190826 106247 190882 106256
rect 190644 106218 190696 106224
rect 190644 101380 190696 101386
rect 190644 101322 190696 101328
rect 190656 91798 190684 101322
rect 190644 91792 190696 91798
rect 190644 91734 190696 91740
rect 190828 91792 190880 91798
rect 190828 91734 190880 91740
rect 190840 87009 190868 91734
rect 190642 87000 190698 87009
rect 190642 86935 190644 86944
rect 190696 86935 190698 86944
rect 190826 87000 190882 87009
rect 190826 86935 190882 86944
rect 190644 86906 190696 86912
rect 190644 80708 190696 80714
rect 190644 80650 190696 80656
rect 190656 70514 190684 80650
rect 190644 70508 190696 70514
rect 190644 70450 190696 70456
rect 190644 66292 190696 66298
rect 190644 66234 190696 66240
rect 190656 64666 190684 66234
rect 190644 64660 190696 64666
rect 190644 64602 190696 64608
rect 190736 56636 190788 56642
rect 190736 56578 190788 56584
rect 190748 48346 190776 56578
rect 190644 48340 190696 48346
rect 190644 48282 190696 48288
rect 190736 48340 190788 48346
rect 190736 48282 190788 48288
rect 190656 38690 190684 48282
rect 190644 38684 190696 38690
rect 190644 38626 190696 38632
rect 190736 38684 190788 38690
rect 190736 38626 190788 38632
rect 190748 37262 190776 38626
rect 190736 37256 190788 37262
rect 190736 37198 190788 37204
rect 190644 27736 190696 27742
rect 190644 27678 190696 27684
rect 190656 22166 190684 27678
rect 190644 22160 190696 22166
rect 190644 22102 190696 22108
rect 190736 22024 190788 22030
rect 190736 21966 190788 21972
rect 190748 13530 190776 21966
rect 190736 13524 190788 13530
rect 190736 13466 190788 13472
rect 190552 9172 190604 9178
rect 190552 9114 190604 9120
rect 190828 4548 190880 4554
rect 190828 4490 190880 4496
rect 190460 4276 190512 4282
rect 190460 4218 190512 4224
rect 189632 4072 189684 4078
rect 189632 4014 189684 4020
rect 188620 2984 188672 2990
rect 188620 2926 188672 2932
rect 189644 480 189672 4014
rect 190840 480 190868 4490
rect 191116 2854 191144 241606
rect 191392 239358 191420 244038
rect 192404 242214 192432 244052
rect 192392 242208 192444 242214
rect 192392 242150 192444 242156
rect 191380 239352 191432 239358
rect 192588 239306 192616 244174
rect 191380 239294 191432 239300
rect 192036 239278 192616 239306
rect 193324 244038 193614 244066
rect 192036 231826 192064 239278
rect 191944 231798 192064 231826
rect 191944 225010 191972 231798
rect 191932 225004 191984 225010
rect 191932 224946 191984 224952
rect 191932 222216 191984 222222
rect 191746 222184 191802 222193
rect 191746 222119 191802 222128
rect 191930 222184 191932 222193
rect 191984 222184 191986 222193
rect 191930 222119 191986 222128
rect 191760 212566 191788 222119
rect 191748 212560 191800 212566
rect 191748 212502 191800 212508
rect 192024 212560 192076 212566
rect 192024 212502 192076 212508
rect 192036 205766 192064 212502
rect 192024 205760 192076 205766
rect 192024 205702 192076 205708
rect 192024 205624 192076 205630
rect 192024 205566 192076 205572
rect 192036 203017 192064 205566
rect 192022 203008 192078 203017
rect 192022 202943 192078 202952
rect 191838 202872 191894 202881
rect 191838 202807 191894 202816
rect 191852 193254 191880 202807
rect 191840 193248 191892 193254
rect 192024 193248 192076 193254
rect 191840 193190 191892 193196
rect 192022 193216 192024 193225
rect 192076 193216 192078 193225
rect 192022 193151 192078 193160
rect 192206 193216 192262 193225
rect 192206 193151 192262 193160
rect 192220 186130 192248 193151
rect 192036 186102 192248 186130
rect 192036 183462 192064 186102
rect 192024 183456 192076 183462
rect 192024 183398 192076 183404
rect 192024 173936 192076 173942
rect 192024 173878 192076 173884
rect 192036 162897 192064 173878
rect 192022 162888 192078 162897
rect 192022 162823 192078 162832
rect 192114 162752 192170 162761
rect 192114 162687 192170 162696
rect 192128 144945 192156 162687
rect 191930 144936 191986 144945
rect 191840 144900 191892 144906
rect 191930 144871 191932 144880
rect 191840 144842 191892 144848
rect 191984 144871 191986 144880
rect 192114 144936 192170 144945
rect 192114 144871 192170 144880
rect 191932 144842 191984 144848
rect 191852 135289 191880 144842
rect 191838 135280 191894 135289
rect 191838 135215 191894 135224
rect 192022 135280 192078 135289
rect 192022 135215 192078 135224
rect 192036 132462 192064 135215
rect 192024 132456 192076 132462
rect 192024 132398 192076 132404
rect 192024 124160 192076 124166
rect 192024 124102 192076 124108
rect 192036 113286 192064 124102
rect 192024 113280 192076 113286
rect 192024 113222 192076 113228
rect 191932 111852 191984 111858
rect 191932 111794 191984 111800
rect 191944 111761 191972 111794
rect 191746 111752 191802 111761
rect 191746 111687 191802 111696
rect 191930 111752 191986 111761
rect 191930 111687 191986 111696
rect 191760 102202 191788 111687
rect 191748 102196 191800 102202
rect 191748 102138 191800 102144
rect 192208 102196 192260 102202
rect 192208 102138 192260 102144
rect 192220 99226 192248 102138
rect 192128 99198 192248 99226
rect 192128 92546 192156 99198
rect 192024 92540 192076 92546
rect 192024 92482 192076 92488
rect 192116 92540 192168 92546
rect 192116 92482 192168 92488
rect 192036 91610 192064 92482
rect 191944 91582 192064 91610
rect 191944 86970 191972 91582
rect 191932 86964 191984 86970
rect 191932 86906 191984 86912
rect 192024 75948 192076 75954
rect 192024 75890 192076 75896
rect 192036 70514 192064 75890
rect 192024 70508 192076 70514
rect 192024 70450 192076 70456
rect 191932 70372 191984 70378
rect 191932 70314 191984 70320
rect 191944 66230 191972 70314
rect 191932 66224 191984 66230
rect 191932 66166 191984 66172
rect 192116 66224 192168 66230
rect 192116 66166 192168 66172
rect 192128 55350 192156 66166
rect 192116 55344 192168 55350
rect 192116 55286 192168 55292
rect 192024 53848 192076 53854
rect 192024 53790 192076 53796
rect 192036 45914 192064 53790
rect 191944 45886 192064 45914
rect 191944 44169 191972 45886
rect 191930 44160 191986 44169
rect 191930 44095 191986 44104
rect 192114 44160 192170 44169
rect 192114 44095 192170 44104
rect 192128 35714 192156 44095
rect 191944 35686 192156 35714
rect 191944 27674 191972 35686
rect 191932 27668 191984 27674
rect 191932 27610 191984 27616
rect 191932 26308 191984 26314
rect 191932 26250 191984 26256
rect 191944 26217 191972 26250
rect 191746 26208 191802 26217
rect 191746 26143 191802 26152
rect 191930 26208 191986 26217
rect 191930 26143 191986 26152
rect 191760 21418 191788 26143
rect 191748 21412 191800 21418
rect 191748 21354 191800 21360
rect 191932 9716 191984 9722
rect 191932 9658 191984 9664
rect 191944 9602 191972 9658
rect 191852 9574 191972 9602
rect 191852 4214 191880 9574
rect 193324 9246 193352 244038
rect 194244 242486 194272 244052
rect 194612 244038 194810 244066
rect 194232 242480 194284 242486
rect 194232 242422 194284 242428
rect 194508 216640 194560 216646
rect 194508 216582 194560 216588
rect 194520 198801 194548 216582
rect 194506 198792 194562 198801
rect 194506 198727 194562 198736
rect 194506 44160 194562 44169
rect 194506 44095 194562 44104
rect 194520 34542 194548 44095
rect 194508 34536 194560 34542
rect 194508 34478 194560 34484
rect 193312 9240 193364 9246
rect 193312 9182 193364 9188
rect 194612 7682 194640 244038
rect 194980 235958 195008 244174
rect 196084 242622 196112 244052
rect 196072 242616 196124 242622
rect 196072 242558 196124 242564
rect 196072 239352 196124 239358
rect 196072 239294 196124 239300
rect 194968 235952 195020 235958
rect 194968 235894 195020 235900
rect 194968 226364 195020 226370
rect 194968 226306 195020 226312
rect 194980 216646 195008 226306
rect 194968 216640 195020 216646
rect 194968 216582 195020 216588
rect 195980 201612 196032 201618
rect 195980 201554 196032 201560
rect 195992 198801 196020 201554
rect 195978 198792 196034 198801
rect 195978 198727 196034 198736
rect 194782 198520 194838 198529
rect 194782 198455 194838 198464
rect 194796 179382 194824 198455
rect 194784 179376 194836 179382
rect 194784 179318 194836 179324
rect 194784 169788 194836 169794
rect 194784 169730 194836 169736
rect 194796 168366 194824 169730
rect 194784 168360 194836 168366
rect 194784 168302 194836 168308
rect 194876 158772 194928 158778
rect 194876 158714 194928 158720
rect 194888 157162 194916 158714
rect 194796 157134 194916 157162
rect 194796 150414 194824 157134
rect 194784 150408 194836 150414
rect 194784 150350 194836 150356
rect 194692 140820 194744 140826
rect 194692 140762 194744 140768
rect 194704 113218 194732 140762
rect 194692 113212 194744 113218
rect 194692 113154 194744 113160
rect 194784 113212 194836 113218
rect 194784 113154 194836 113160
rect 194796 109154 194824 113154
rect 194796 109126 194916 109154
rect 194888 108474 194916 109126
rect 194796 108446 194916 108474
rect 194796 85610 194824 108446
rect 194692 85604 194744 85610
rect 194692 85546 194744 85552
rect 194784 85604 194836 85610
rect 194784 85546 194836 85552
rect 194704 85490 194732 85546
rect 194704 85462 194824 85490
rect 194796 84182 194824 85462
rect 194784 84176 194836 84182
rect 194784 84118 194836 84124
rect 194784 74588 194836 74594
rect 194784 74530 194836 74536
rect 194796 70514 194824 74530
rect 194784 70508 194836 70514
rect 194784 70450 194836 70456
rect 194692 70372 194744 70378
rect 194692 70314 194744 70320
rect 194704 55282 194732 70314
rect 194692 55276 194744 55282
rect 194692 55218 194744 55224
rect 194692 53848 194744 53854
rect 194692 53790 194744 53796
rect 194704 45830 194732 53790
rect 194692 45824 194744 45830
rect 194692 45766 194744 45772
rect 194784 45620 194836 45626
rect 194784 45562 194836 45568
rect 194796 44169 194824 45562
rect 194782 44160 194838 44169
rect 194782 44095 194838 44104
rect 194692 34536 194744 34542
rect 194692 34478 194744 34484
rect 194704 26246 194732 34478
rect 194692 26240 194744 26246
rect 194692 26182 194744 26188
rect 194692 16652 194744 16658
rect 194692 16594 194744 16600
rect 194704 9602 194732 16594
rect 194704 9574 194824 9602
rect 194796 9314 194824 9574
rect 196084 9382 196112 239294
rect 196268 231878 196296 244174
rect 196912 244038 197294 244066
rect 196912 239358 196940 244038
rect 197924 242350 197952 244052
rect 198108 244038 198490 244066
rect 198844 244038 199134 244066
rect 197912 242344 197964 242350
rect 197912 242286 197964 242292
rect 197268 242208 197320 242214
rect 197268 242150 197320 242156
rect 196900 239352 196952 239358
rect 196900 239294 196952 239300
rect 196164 231872 196216 231878
rect 196164 231814 196216 231820
rect 196256 231872 196308 231878
rect 196256 231814 196308 231820
rect 196176 222222 196204 231814
rect 196164 222216 196216 222222
rect 196164 222158 196216 222164
rect 196348 222216 196400 222222
rect 196348 222158 196400 222164
rect 196360 211274 196388 222158
rect 196256 211268 196308 211274
rect 196256 211210 196308 211216
rect 196348 211268 196400 211274
rect 196348 211210 196400 211216
rect 196268 201618 196296 211210
rect 196256 201612 196308 201618
rect 196256 201554 196308 201560
rect 196346 198520 196402 198529
rect 196346 198455 196402 198464
rect 196360 189038 196388 198455
rect 196348 189032 196400 189038
rect 196348 188974 196400 188980
rect 196256 179444 196308 179450
rect 196256 179386 196308 179392
rect 196268 162926 196296 179386
rect 196256 162920 196308 162926
rect 196256 162862 196308 162868
rect 196256 162784 196308 162790
rect 196256 162726 196308 162732
rect 196268 142254 196296 162726
rect 196256 142248 196308 142254
rect 196256 142190 196308 142196
rect 196164 142112 196216 142118
rect 196164 142054 196216 142060
rect 196176 140729 196204 142054
rect 196162 140720 196218 140729
rect 196162 140655 196218 140664
rect 196254 140584 196310 140593
rect 196254 140519 196310 140528
rect 196268 122874 196296 140519
rect 196164 122868 196216 122874
rect 196164 122810 196216 122816
rect 196256 122868 196308 122874
rect 196256 122810 196308 122816
rect 196176 113218 196204 122810
rect 196164 113212 196216 113218
rect 196164 113154 196216 113160
rect 196256 113212 196308 113218
rect 196256 113154 196308 113160
rect 196268 90386 196296 113154
rect 196268 90358 196388 90386
rect 196360 82498 196388 90358
rect 196268 82470 196388 82498
rect 196268 75886 196296 82470
rect 196256 75880 196308 75886
rect 196256 75822 196308 75828
rect 196348 75880 196400 75886
rect 196348 75822 196400 75828
rect 196360 61282 196388 75822
rect 196268 61254 196388 61282
rect 196268 51134 196296 61254
rect 196256 51128 196308 51134
rect 196256 51070 196308 51076
rect 196164 51060 196216 51066
rect 196164 51002 196216 51008
rect 196176 45558 196204 51002
rect 196164 45552 196216 45558
rect 196164 45494 196216 45500
rect 196348 45552 196400 45558
rect 196348 45494 196400 45500
rect 196360 22114 196388 45494
rect 196176 22098 196388 22114
rect 196164 22092 196400 22098
rect 196216 22086 196348 22092
rect 196164 22034 196216 22040
rect 196348 22034 196400 22040
rect 196360 12050 196388 22034
rect 196360 12022 196480 12050
rect 196452 11778 196480 12022
rect 196360 11750 196480 11778
rect 196072 9376 196124 9382
rect 196072 9318 196124 9324
rect 194784 9308 194836 9314
rect 194784 9250 194836 9256
rect 196360 7750 196388 11750
rect 196348 7744 196400 7750
rect 196348 7686 196400 7692
rect 194600 7676 194652 7682
rect 194600 7618 194652 7624
rect 194416 4684 194468 4690
rect 194416 4626 194468 4632
rect 192024 4616 192076 4622
rect 192024 4558 192076 4564
rect 191840 4208 191892 4214
rect 191840 4150 191892 4156
rect 191104 2848 191156 2854
rect 191104 2790 191156 2796
rect 192036 480 192064 4558
rect 193220 3052 193272 3058
rect 193220 2994 193272 3000
rect 193232 480 193260 2994
rect 194428 480 194456 4626
rect 195612 4480 195664 4486
rect 195612 4422 195664 4428
rect 195624 480 195652 4422
rect 197280 4146 197308 242150
rect 198108 239306 198136 244038
rect 198280 242480 198332 242486
rect 198280 242422 198332 242428
rect 198188 242344 198240 242350
rect 198188 242286 198240 242292
rect 197464 239278 198136 239306
rect 197464 7818 197492 239278
rect 198200 238490 198228 242286
rect 198292 241466 198320 242422
rect 198280 241460 198332 241466
rect 198280 241402 198332 241408
rect 198016 238462 198228 238490
rect 197452 7812 197504 7818
rect 197452 7754 197504 7760
rect 196808 4140 196860 4146
rect 196808 4082 196860 4088
rect 197268 4140 197320 4146
rect 197268 4082 197320 4088
rect 196820 480 196848 4082
rect 198016 3058 198044 238462
rect 198280 231872 198332 231878
rect 198280 231814 198332 231820
rect 198292 225010 198320 231814
rect 198280 225004 198332 225010
rect 198280 224946 198332 224952
rect 198372 224868 198424 224874
rect 198372 224810 198424 224816
rect 198384 211177 198412 224810
rect 198186 211168 198242 211177
rect 198186 211103 198188 211112
rect 198240 211103 198242 211112
rect 198370 211168 198426 211177
rect 198370 211103 198372 211112
rect 198188 211074 198240 211080
rect 198424 211103 198426 211112
rect 198372 211074 198424 211080
rect 198384 201618 198412 211074
rect 198372 201612 198424 201618
rect 198372 201554 198424 201560
rect 198372 201476 198424 201482
rect 198372 201418 198424 201424
rect 198384 189106 198412 201418
rect 198280 189100 198332 189106
rect 198280 189042 198332 189048
rect 198372 189100 198424 189106
rect 198372 189042 198424 189048
rect 198292 162858 198320 189042
rect 198280 162852 198332 162858
rect 198280 162794 198332 162800
rect 198372 162852 198424 162858
rect 198372 162794 198424 162800
rect 198384 158710 198412 162794
rect 198372 158704 198424 158710
rect 198372 158646 198424 158652
rect 198280 149116 198332 149122
rect 198280 149058 198332 149064
rect 198292 138106 198320 149058
rect 198280 138100 198332 138106
rect 198280 138042 198332 138048
rect 198280 137964 198332 137970
rect 198280 137906 198332 137912
rect 198292 113234 198320 137906
rect 198200 113206 198320 113234
rect 198200 109154 198228 113206
rect 198200 109126 198412 109154
rect 198384 108882 198412 109126
rect 198292 108854 198412 108882
rect 198292 98734 198320 108854
rect 198280 98728 198332 98734
rect 198280 98670 198332 98676
rect 198280 98592 198332 98598
rect 198280 98534 198332 98540
rect 198292 76022 198320 98534
rect 198280 76016 198332 76022
rect 198280 75958 198332 75964
rect 198188 75948 198240 75954
rect 198188 75890 198240 75896
rect 198200 74526 198228 75890
rect 198188 74520 198240 74526
rect 198188 74462 198240 74468
rect 198280 74520 198332 74526
rect 198280 74462 198332 74468
rect 198292 64954 198320 74462
rect 198200 64926 198320 64954
rect 198200 63510 198228 64926
rect 198188 63504 198240 63510
rect 198188 63446 198240 63452
rect 198188 53848 198240 53854
rect 198188 53790 198240 53796
rect 198200 50402 198228 53790
rect 198200 50374 198320 50402
rect 198292 40746 198320 50374
rect 198200 40718 198320 40746
rect 198200 27674 198228 40718
rect 198188 27668 198240 27674
rect 198188 27610 198240 27616
rect 198280 27668 198332 27674
rect 198280 27610 198332 27616
rect 198292 22166 198320 27610
rect 198280 22160 198332 22166
rect 198280 22102 198332 22108
rect 198188 22092 198240 22098
rect 198188 22034 198240 22040
rect 198200 14634 198228 22034
rect 198200 14606 198320 14634
rect 198292 14362 198320 14606
rect 198200 14334 198320 14362
rect 198096 4412 198148 4418
rect 198096 4354 198148 4360
rect 198004 3052 198056 3058
rect 198004 2994 198056 3000
rect 198108 2258 198136 4354
rect 198200 4078 198228 14334
rect 198844 9450 198872 244038
rect 199672 242894 199700 244052
rect 200224 244038 200330 244066
rect 199660 242888 199712 242894
rect 199660 242830 199712 242836
rect 199384 242752 199436 242758
rect 199384 242694 199436 242700
rect 198832 9444 198884 9450
rect 198832 9386 198884 9392
rect 199200 4140 199252 4146
rect 199200 4082 199252 4088
rect 198188 4072 198240 4078
rect 198188 4014 198240 4020
rect 198016 2230 198136 2258
rect 198016 480 198044 2230
rect 199212 480 199240 4082
rect 199396 4010 199424 242694
rect 200224 7886 200252 244038
rect 200960 242282 200988 244052
rect 201512 242418 201540 244052
rect 201696 244038 202170 244066
rect 202432 244038 202814 244066
rect 201500 242412 201552 242418
rect 201500 242354 201552 242360
rect 200948 242276 201000 242282
rect 200948 242218 201000 242224
rect 201408 242276 201460 242282
rect 201408 242218 201460 242224
rect 200764 242004 200816 242010
rect 200764 241946 200816 241952
rect 200212 7880 200264 7886
rect 200212 7822 200264 7828
rect 200776 4350 200804 241946
rect 200764 4344 200816 4350
rect 200764 4286 200816 4292
rect 199384 4004 199436 4010
rect 199384 3946 199436 3952
rect 201420 3398 201448 242218
rect 201592 239352 201644 239358
rect 201592 239294 201644 239300
rect 201498 40216 201554 40225
rect 201498 40151 201500 40160
rect 201552 40151 201554 40160
rect 201500 40122 201552 40128
rect 201604 9518 201632 239294
rect 201592 9512 201644 9518
rect 201592 9454 201644 9460
rect 201696 7954 201724 244038
rect 202144 242072 202196 242078
rect 202144 242014 202196 242020
rect 201684 7948 201736 7954
rect 201684 7890 201736 7896
rect 201500 4344 201552 4350
rect 201500 4286 201552 4292
rect 200396 3392 200448 3398
rect 200396 3334 200448 3340
rect 201408 3392 201460 3398
rect 201408 3334 201460 3340
rect 200408 480 200436 3334
rect 201512 480 201540 4286
rect 202156 3942 202184 242014
rect 202432 239358 202460 244038
rect 203352 242146 203380 244052
rect 203536 244038 204010 244066
rect 204364 244038 204654 244066
rect 204824 244038 205206 244066
rect 205652 244038 205850 244066
rect 203340 242140 203392 242146
rect 203340 242082 203392 242088
rect 202420 239352 202472 239358
rect 203536 239306 203564 244038
rect 203616 242548 203668 242554
rect 203616 242490 203668 242496
rect 202420 239294 202472 239300
rect 202984 239278 203564 239306
rect 202984 8022 203012 239278
rect 203628 238626 203656 242490
rect 204168 242412 204220 242418
rect 204168 242354 204220 242360
rect 203536 238598 203656 238626
rect 202972 8016 203024 8022
rect 202972 7958 203024 7964
rect 203536 4146 203564 238598
rect 203524 4140 203576 4146
rect 203524 4082 203576 4088
rect 202696 4004 202748 4010
rect 202696 3946 202748 3952
rect 202144 3936 202196 3942
rect 202144 3878 202196 3884
rect 202708 480 202736 3946
rect 204180 626 204208 242354
rect 204364 9586 204392 244038
rect 204824 241874 204852 244038
rect 204812 241868 204864 241874
rect 204812 241810 204864 241816
rect 204904 241868 204956 241874
rect 204904 241810 204956 241816
rect 204352 9580 204404 9586
rect 204352 9522 204404 9528
rect 204916 3874 204944 241810
rect 205652 8090 205680 244038
rect 206020 239306 206048 244174
rect 207032 241942 207060 244052
rect 207020 241936 207072 241942
rect 207020 241878 207072 241884
rect 205928 239278 206048 239306
rect 205928 222222 205956 239278
rect 207216 230518 207244 244174
rect 208228 241534 208256 244052
rect 208308 242616 208360 242622
rect 208308 242558 208360 242564
rect 208216 241528 208268 241534
rect 208216 241470 208268 241476
rect 207112 230512 207164 230518
rect 207112 230454 207164 230460
rect 207204 230512 207256 230518
rect 207204 230454 207256 230460
rect 205824 222216 205876 222222
rect 205824 222158 205876 222164
rect 205916 222216 205968 222222
rect 205916 222158 205968 222164
rect 205836 219450 205864 222158
rect 207124 220833 207152 230454
rect 206926 220824 206982 220833
rect 206926 220759 206982 220768
rect 207110 220824 207166 220833
rect 207110 220759 207166 220768
rect 205836 219422 205956 219450
rect 205928 206310 205956 219422
rect 206940 211177 206968 220759
rect 206926 211168 206982 211177
rect 206926 211103 206982 211112
rect 207110 211168 207166 211177
rect 207110 211103 207166 211112
rect 207124 207754 207152 211103
rect 207124 207726 207244 207754
rect 205916 206304 205968 206310
rect 205916 206246 205968 206252
rect 206100 206304 206152 206310
rect 206100 206246 206152 206252
rect 206112 201521 206140 206246
rect 205914 201512 205970 201521
rect 205914 201447 205916 201456
rect 205968 201447 205970 201456
rect 206098 201512 206154 201521
rect 206098 201447 206154 201456
rect 205916 201418 205968 201424
rect 206008 201408 206060 201414
rect 206008 201350 206060 201356
rect 206020 178786 206048 201350
rect 207216 193254 207244 207726
rect 207020 193248 207072 193254
rect 207020 193190 207072 193196
rect 207204 193248 207256 193254
rect 207204 193190 207256 193196
rect 207032 189530 207060 193190
rect 207032 189502 207244 189530
rect 206020 178758 206140 178786
rect 206112 173942 206140 178758
rect 207216 173942 207244 189502
rect 205916 173936 205968 173942
rect 205916 173878 205968 173884
rect 206100 173936 206152 173942
rect 206100 173878 206152 173884
rect 207020 173936 207072 173942
rect 207020 173878 207072 173884
rect 207204 173936 207256 173942
rect 207204 173878 207256 173884
rect 205928 169402 205956 173878
rect 207032 169402 207060 173878
rect 205928 169374 206048 169402
rect 207032 169374 207152 169402
rect 206020 162858 206048 169374
rect 206008 162852 206060 162858
rect 206008 162794 206060 162800
rect 207124 157486 207152 169374
rect 207112 157480 207164 157486
rect 207112 157422 207164 157428
rect 206008 157344 206060 157350
rect 206008 157286 206060 157292
rect 207112 157344 207164 157350
rect 207112 157286 207164 157292
rect 206020 144906 206048 157286
rect 207124 144906 207152 157286
rect 205916 144900 205968 144906
rect 205916 144842 205968 144848
rect 206008 144900 206060 144906
rect 206008 144842 206060 144848
rect 207112 144900 207164 144906
rect 207112 144842 207164 144848
rect 207204 144900 207256 144906
rect 207204 144842 207256 144848
rect 205928 143546 205956 144842
rect 205916 143540 205968 143546
rect 205916 143482 205968 143488
rect 206100 143540 206152 143546
rect 206100 143482 206152 143488
rect 206112 128330 206140 143482
rect 207216 135289 207244 144842
rect 207018 135280 207074 135289
rect 207018 135215 207074 135224
rect 207202 135280 207258 135289
rect 207202 135215 207258 135224
rect 207032 130370 207060 135215
rect 207032 130342 207152 130370
rect 206020 128302 206140 128330
rect 206020 125594 206048 128302
rect 205824 125588 205876 125594
rect 205824 125530 205876 125536
rect 206008 125588 206060 125594
rect 206008 125530 206060 125536
rect 205836 118674 205864 125530
rect 205836 118646 205956 118674
rect 205928 109698 205956 118646
rect 207124 116113 207152 130342
rect 207110 116104 207166 116113
rect 207110 116039 207166 116048
rect 207018 115968 207074 115977
rect 207018 115903 207074 115912
rect 207032 114510 207060 115903
rect 207020 114504 207072 114510
rect 207020 114446 207072 114452
rect 205836 109670 205956 109698
rect 205836 104922 205864 109670
rect 205824 104916 205876 104922
rect 205824 104858 205876 104864
rect 206008 104916 206060 104922
rect 206008 104858 206060 104864
rect 207112 104916 207164 104922
rect 207112 104858 207164 104864
rect 206020 103494 206048 104858
rect 206008 103488 206060 103494
rect 206008 103430 206060 103436
rect 207124 95266 207152 104858
rect 207112 95260 207164 95266
rect 207112 95202 207164 95208
rect 207204 95124 207256 95130
rect 207204 95066 207256 95072
rect 206008 93900 206060 93906
rect 206008 93842 206060 93848
rect 206020 87038 206048 93842
rect 206008 87032 206060 87038
rect 206008 86974 206060 86980
rect 207216 85610 207244 95066
rect 206008 85604 206060 85610
rect 206008 85546 206060 85552
rect 207020 85604 207072 85610
rect 207020 85546 207072 85552
rect 207204 85604 207256 85610
rect 207204 85546 207256 85552
rect 206020 82090 206048 85546
rect 207032 84182 207060 85546
rect 207020 84176 207072 84182
rect 207020 84118 207072 84124
rect 205928 82062 206048 82090
rect 205928 51082 205956 82062
rect 207112 66292 207164 66298
rect 207112 66234 207164 66240
rect 207124 64870 207152 66234
rect 207112 64864 207164 64870
rect 207112 64806 207164 64812
rect 207112 56364 207164 56370
rect 207112 56306 207164 56312
rect 205836 51054 205956 51082
rect 205836 41426 205864 51054
rect 207124 46918 207152 56306
rect 207112 46912 207164 46918
rect 207112 46854 207164 46860
rect 205744 41398 205864 41426
rect 205744 29034 205772 41398
rect 205732 29028 205784 29034
rect 205732 28970 205784 28976
rect 205824 29028 205876 29034
rect 205824 28970 205876 28976
rect 205836 27606 205864 28970
rect 207112 27736 207164 27742
rect 207112 27678 207164 27684
rect 207124 27606 207152 27678
rect 205824 27600 205876 27606
rect 205824 27542 205876 27548
rect 205916 27600 205968 27606
rect 205916 27542 205968 27548
rect 207112 27600 207164 27606
rect 207112 27542 207164 27548
rect 205928 12322 205956 27542
rect 207204 18012 207256 18018
rect 207204 17954 207256 17960
rect 205836 12294 205956 12322
rect 205836 9654 205864 12294
rect 205824 9648 205876 9654
rect 205824 9590 205876 9596
rect 207216 8158 207244 17954
rect 207204 8152 207256 8158
rect 207204 8094 207256 8100
rect 205640 8084 205692 8090
rect 205640 8026 205692 8032
rect 205088 4276 205140 4282
rect 205088 4218 205140 4224
rect 204904 3868 204956 3874
rect 204904 3810 204956 3816
rect 203904 598 204208 626
rect 203904 480 203932 598
rect 205100 480 205128 4218
rect 208320 4146 208348 242558
rect 208872 241806 208900 244052
rect 209148 244038 209530 244066
rect 209884 244038 210082 244066
rect 208860 241800 208912 241806
rect 208860 241742 208912 241748
rect 209148 231878 209176 244038
rect 208492 231872 208544 231878
rect 208492 231814 208544 231820
rect 209136 231872 209188 231878
rect 209136 231814 209188 231820
rect 208504 202910 208532 231814
rect 208492 202904 208544 202910
rect 208492 202846 208544 202852
rect 208584 202904 208636 202910
rect 208584 202846 208636 202852
rect 208596 201482 208624 202846
rect 208400 201476 208452 201482
rect 208400 201418 208452 201424
rect 208584 201476 208636 201482
rect 208584 201418 208636 201424
rect 208412 191865 208440 201418
rect 208398 191856 208454 191865
rect 208398 191791 208454 191800
rect 208582 191856 208638 191865
rect 208582 191791 208638 191800
rect 208596 188442 208624 191791
rect 208504 188414 208624 188442
rect 208504 173942 208532 188414
rect 208492 173936 208544 173942
rect 208492 173878 208544 173884
rect 208584 173936 208636 173942
rect 208584 173878 208636 173884
rect 208596 164234 208624 173878
rect 208504 164206 208624 164234
rect 208504 157486 208532 164206
rect 208492 157480 208544 157486
rect 208492 157422 208544 157428
rect 208492 157344 208544 157350
rect 208492 157286 208544 157292
rect 208504 144906 208532 157286
rect 208492 144900 208544 144906
rect 208492 144842 208544 144848
rect 208676 144900 208728 144906
rect 208676 144842 208728 144848
rect 208688 139890 208716 144842
rect 208596 139862 208716 139890
rect 208596 125610 208624 139862
rect 208504 125594 208624 125610
rect 208492 125588 208624 125594
rect 208544 125582 208624 125588
rect 208676 125588 208728 125594
rect 208492 125530 208544 125536
rect 208676 125530 208728 125536
rect 208688 120562 208716 125530
rect 208584 120556 208636 120562
rect 208584 120498 208636 120504
rect 208676 120556 208728 120562
rect 208676 120498 208728 120504
rect 208596 106350 208624 120498
rect 208584 106344 208636 106350
rect 208584 106286 208636 106292
rect 208400 104916 208452 104922
rect 208400 104858 208452 104864
rect 208412 103494 208440 104858
rect 208400 103488 208452 103494
rect 208400 103430 208452 103436
rect 208768 95124 208820 95130
rect 208768 95066 208820 95072
rect 208780 85649 208808 95066
rect 208582 85640 208638 85649
rect 208582 85575 208638 85584
rect 208766 85640 208822 85649
rect 208766 85575 208822 85584
rect 208596 84182 208624 85575
rect 208584 84176 208636 84182
rect 208584 84118 208636 84124
rect 208492 66360 208544 66366
rect 208492 66302 208544 66308
rect 208504 64870 208532 66302
rect 208492 64864 208544 64870
rect 208492 64806 208544 64812
rect 208492 55276 208544 55282
rect 208492 55218 208544 55224
rect 208504 51762 208532 55218
rect 208504 51734 208624 51762
rect 208596 42090 208624 51734
rect 208584 42084 208636 42090
rect 208584 42026 208636 42032
rect 208584 29028 208636 29034
rect 208584 28970 208636 28976
rect 208596 22114 208624 28970
rect 208504 22086 208624 22114
rect 208504 21978 208532 22086
rect 208504 21950 208624 21978
rect 208596 8226 208624 21950
rect 209884 8906 209912 244038
rect 210712 242894 210740 244052
rect 211172 244038 211370 244066
rect 210700 242888 210752 242894
rect 210700 242830 210752 242836
rect 209872 8900 209924 8906
rect 209872 8842 209924 8848
rect 211172 8294 211200 244038
rect 211540 231878 211568 244174
rect 211896 242888 211948 242894
rect 211896 242830 211948 242836
rect 211804 242684 211856 242690
rect 211804 242626 211856 242632
rect 211252 231872 211304 231878
rect 211252 231814 211304 231820
rect 211528 231872 211580 231878
rect 211528 231814 211580 231820
rect 211264 202910 211292 231814
rect 211252 202904 211304 202910
rect 211252 202846 211304 202852
rect 211344 202904 211396 202910
rect 211344 202846 211396 202852
rect 211356 188442 211384 202846
rect 211264 188414 211384 188442
rect 211264 173942 211292 188414
rect 211252 173936 211304 173942
rect 211252 173878 211304 173884
rect 211344 173936 211396 173942
rect 211344 173878 211396 173884
rect 211356 162874 211384 173878
rect 211264 162846 211384 162874
rect 211264 157418 211292 162846
rect 211252 157412 211304 157418
rect 211252 157354 211304 157360
rect 211252 157276 211304 157282
rect 211252 157218 211304 157224
rect 211264 144906 211292 157218
rect 211252 144900 211304 144906
rect 211252 144842 211304 144848
rect 211436 144900 211488 144906
rect 211436 144842 211488 144848
rect 211448 137714 211476 144842
rect 211356 137686 211476 137714
rect 211356 130370 211384 137686
rect 211264 130342 211384 130370
rect 211264 125594 211292 130342
rect 211252 125588 211304 125594
rect 211252 125530 211304 125536
rect 211344 125520 211396 125526
rect 211344 125462 211396 125468
rect 211356 106350 211384 125462
rect 211344 106344 211396 106350
rect 211344 106286 211396 106292
rect 211344 106140 211396 106146
rect 211344 106082 211396 106088
rect 211356 95198 211384 106082
rect 211344 95192 211396 95198
rect 211344 95134 211396 95140
rect 211344 85604 211396 85610
rect 211344 85546 211396 85552
rect 211356 74610 211384 85546
rect 211264 74582 211384 74610
rect 211264 74526 211292 74582
rect 211252 74520 211304 74526
rect 211252 74462 211304 74468
rect 211344 65000 211396 65006
rect 211344 64942 211396 64948
rect 211356 64870 211384 64942
rect 211344 64864 211396 64870
rect 211344 64806 211396 64812
rect 211528 55276 211580 55282
rect 211528 55218 211580 55224
rect 211540 47326 211568 55218
rect 211528 47320 211580 47326
rect 211528 47262 211580 47268
rect 211252 45620 211304 45626
rect 211252 45562 211304 45568
rect 211264 27606 211292 45562
rect 211252 27600 211304 27606
rect 211252 27542 211304 27548
rect 211344 19372 211396 19378
rect 211344 19314 211396 19320
rect 211356 8838 211384 19314
rect 211344 8832 211396 8838
rect 211344 8774 211396 8780
rect 211160 8288 211212 8294
rect 211160 8230 211212 8236
rect 208584 8220 208636 8226
rect 208584 8162 208636 8168
rect 211816 4146 211844 242626
rect 207480 4140 207532 4146
rect 207480 4082 207532 4088
rect 208308 4140 208360 4146
rect 208308 4082 208360 4088
rect 211068 4140 211120 4146
rect 211068 4082 211120 4088
rect 211804 4140 211856 4146
rect 211804 4082 211856 4088
rect 206284 3052 206336 3058
rect 206284 2994 206336 3000
rect 206296 480 206324 2994
rect 207492 480 207520 4082
rect 208676 3868 208728 3874
rect 208676 3810 208728 3816
rect 208688 480 208716 3810
rect 209872 3256 209924 3262
rect 209872 3198 209924 3204
rect 209884 480 209912 3198
rect 211080 480 211108 4082
rect 211908 3942 211936 242830
rect 212552 241738 212580 244052
rect 212736 244038 213210 244066
rect 213472 244038 213762 244066
rect 212540 241732 212592 241738
rect 212540 241674 212592 241680
rect 212632 239352 212684 239358
rect 212632 239294 212684 239300
rect 212644 8770 212672 239294
rect 212632 8764 212684 8770
rect 212632 8706 212684 8712
rect 212736 7546 212764 244038
rect 213472 239358 213500 244038
rect 213826 242176 213882 242185
rect 213826 242111 213882 242120
rect 213460 239352 213512 239358
rect 213460 239294 213512 239300
rect 212724 7540 212776 7546
rect 212724 7482 212776 7488
rect 212264 4208 212316 4214
rect 212264 4150 212316 4156
rect 211896 3936 211948 3942
rect 211896 3878 211948 3884
rect 212276 480 212304 4150
rect 213840 626 213868 242111
rect 214392 241670 214420 244052
rect 214668 244038 215050 244066
rect 215404 244038 215602 244066
rect 215864 244038 216246 244066
rect 216692 244038 216798 244066
rect 217152 244038 217442 244066
rect 214380 241664 214432 241670
rect 214380 241606 214432 241612
rect 214668 239306 214696 244038
rect 215208 242140 215260 242146
rect 215208 242082 215260 242088
rect 214116 239278 214696 239306
rect 214116 219450 214144 239278
rect 214024 219422 214144 219450
rect 214024 209846 214052 219422
rect 214012 209840 214064 209846
rect 214012 209782 214064 209788
rect 214012 202904 214064 202910
rect 214012 202846 214064 202852
rect 214024 193254 214052 202846
rect 214012 193248 214064 193254
rect 214012 193190 214064 193196
rect 214104 193248 214156 193254
rect 214104 193190 214156 193196
rect 214116 176610 214144 193190
rect 214024 176582 214144 176610
rect 214024 176338 214052 176582
rect 214024 176310 214144 176338
rect 214116 157434 214144 176310
rect 214024 157406 214144 157434
rect 214024 157298 214052 157406
rect 214024 157270 214144 157298
rect 214116 99482 214144 157270
rect 214104 99476 214156 99482
rect 214104 99418 214156 99424
rect 214104 99340 214156 99346
rect 214104 99282 214156 99288
rect 214116 80730 214144 99282
rect 214116 80702 214236 80730
rect 214208 58002 214236 80702
rect 214104 57996 214156 58002
rect 214104 57938 214156 57944
rect 214196 57996 214248 58002
rect 214196 57938 214248 57944
rect 214116 48362 214144 57938
rect 214024 48334 214144 48362
rect 214024 46918 214052 48334
rect 214012 46912 214064 46918
rect 214012 46854 214064 46860
rect 213920 32428 213972 32434
rect 213920 32370 213972 32376
rect 213932 19394 213960 32370
rect 213932 19366 214052 19394
rect 214024 15178 214052 19366
rect 214024 15150 214144 15178
rect 214116 7410 214144 15150
rect 214104 7404 214156 7410
rect 214104 7346 214156 7352
rect 215220 4146 215248 242082
rect 215300 239352 215352 239358
rect 215300 239294 215352 239300
rect 215312 6118 215340 239294
rect 215404 7478 215432 244038
rect 215864 239358 215892 244038
rect 215852 239352 215904 239358
rect 215852 239294 215904 239300
rect 216586 183560 216642 183569
rect 216586 183495 216642 183504
rect 216600 179042 216628 183495
rect 216588 179036 216640 179042
rect 216588 178978 216640 178984
rect 215392 7472 215444 7478
rect 215392 7414 215444 7420
rect 216692 7342 216720 244038
rect 217152 239340 217180 244038
rect 216876 239312 217180 239340
rect 216876 220930 216904 239312
rect 216772 220924 216824 220930
rect 216772 220866 216824 220872
rect 216864 220924 216916 220930
rect 216864 220866 216916 220872
rect 216784 220794 216812 220866
rect 216772 220788 216824 220794
rect 216772 220730 216824 220736
rect 216956 220788 217008 220794
rect 216956 220730 217008 220736
rect 216968 219434 216996 220730
rect 216956 219428 217008 219434
rect 216956 219370 217008 219376
rect 216956 211132 217008 211138
rect 216956 211074 217008 211080
rect 216968 206258 216996 211074
rect 216968 206230 217180 206258
rect 217152 196466 217180 206230
rect 216876 196438 217180 196466
rect 216876 188442 216904 196438
rect 216784 188414 216904 188442
rect 216784 183569 216812 188414
rect 216770 183560 216826 183569
rect 216770 183495 216826 183504
rect 216864 179036 216916 179042
rect 216864 178978 216916 178984
rect 216876 163033 216904 178978
rect 216862 163024 216918 163033
rect 216862 162959 216918 162968
rect 216770 162888 216826 162897
rect 216770 162823 216826 162832
rect 216784 161430 216812 162823
rect 216772 161424 216824 161430
rect 216772 161366 216824 161372
rect 217968 161424 218020 161430
rect 217968 161366 218020 161372
rect 217980 151881 218008 161366
rect 217966 151872 218022 151881
rect 216864 151836 216916 151842
rect 217966 151807 218022 151816
rect 216864 151778 216916 151784
rect 216876 148322 216904 151778
rect 217966 151736 218022 151745
rect 217966 151671 218022 151680
rect 216876 148294 216996 148322
rect 216968 137850 216996 148294
rect 217980 142186 218008 151671
rect 217968 142180 218020 142186
rect 217968 142122 218020 142128
rect 216876 137822 216996 137850
rect 216876 135250 216904 137822
rect 216864 135244 216916 135250
rect 216864 135186 216916 135192
rect 216772 129736 216824 129742
rect 216772 129678 216824 129684
rect 216784 125594 216812 129678
rect 216772 125588 216824 125594
rect 216772 125530 216824 125536
rect 216956 125588 217008 125594
rect 216956 125530 217008 125536
rect 216968 114646 216996 125530
rect 216956 114640 217008 114646
rect 216956 114582 217008 114588
rect 216864 114572 216916 114578
rect 216864 114514 216916 114520
rect 216876 95198 216904 114514
rect 216864 95192 216916 95198
rect 216864 95134 216916 95140
rect 216864 85604 216916 85610
rect 216864 85546 216916 85552
rect 216876 70514 216904 85546
rect 216864 70508 216916 70514
rect 216864 70450 216916 70456
rect 216772 70372 216824 70378
rect 216772 70314 216824 70320
rect 216784 61418 216812 70314
rect 216784 61390 216904 61418
rect 216876 56574 216904 61390
rect 216864 56568 216916 56574
rect 216864 56510 216916 56516
rect 216956 56568 217008 56574
rect 216956 56510 217008 56516
rect 216968 55214 216996 56510
rect 216956 55208 217008 55214
rect 216956 55150 217008 55156
rect 216956 45620 217008 45626
rect 216956 45562 217008 45568
rect 216968 26058 216996 45562
rect 216876 26030 216996 26058
rect 216876 12510 216904 26030
rect 216864 12504 216916 12510
rect 216864 12446 216916 12452
rect 216772 12436 216824 12442
rect 216772 12378 216824 12384
rect 216784 8702 216812 12378
rect 216772 8696 216824 8702
rect 216772 8638 216824 8644
rect 216680 7336 216732 7342
rect 216680 7278 216732 7284
rect 215300 6112 215352 6118
rect 215300 6054 215352 6060
rect 218072 6050 218100 244052
rect 218348 244038 218638 244066
rect 218992 244038 219282 244066
rect 219452 244038 219926 244066
rect 220188 244038 220478 244066
rect 220924 244038 221122 244066
rect 221384 244038 221766 244066
rect 218348 239340 218376 244038
rect 218164 239312 218376 239340
rect 218164 7274 218192 239312
rect 218992 229129 219020 244038
rect 218426 229120 218482 229129
rect 218426 229055 218482 229064
rect 218978 229120 219034 229129
rect 218978 229055 219034 229064
rect 218440 225010 218468 229055
rect 218428 225004 218480 225010
rect 218428 224946 218480 224952
rect 218244 224936 218296 224942
rect 218244 224878 218296 224884
rect 218256 220794 218284 224878
rect 218244 220788 218296 220794
rect 218244 220730 218296 220736
rect 218336 220788 218388 220794
rect 218336 220730 218388 220736
rect 218348 219434 218376 220730
rect 218336 219428 218388 219434
rect 218336 219370 218388 219376
rect 218244 205624 218296 205630
rect 218244 205566 218296 205572
rect 218256 201482 218284 205566
rect 218244 201476 218296 201482
rect 218244 201418 218296 201424
rect 218336 193180 218388 193186
rect 218336 193122 218388 193128
rect 218348 191842 218376 193122
rect 218348 191814 218468 191842
rect 218440 183598 218468 191814
rect 218244 183592 218296 183598
rect 218244 183534 218296 183540
rect 218428 183592 218480 183598
rect 218428 183534 218480 183540
rect 218256 183462 218284 183534
rect 218244 183456 218296 183462
rect 218244 183398 218296 183404
rect 218336 180056 218388 180062
rect 218336 179998 218388 180004
rect 218348 163033 218376 179998
rect 218334 163024 218390 163033
rect 218334 162959 218390 162968
rect 218242 162888 218298 162897
rect 218242 162823 218298 162832
rect 218256 161430 218284 162823
rect 218244 161424 218296 161430
rect 218244 161366 218296 161372
rect 218428 142180 218480 142186
rect 218428 142122 218480 142128
rect 218440 137850 218468 142122
rect 218348 137822 218468 137850
rect 218348 128450 218376 137822
rect 218336 128444 218388 128450
rect 218336 128386 218388 128392
rect 218244 128308 218296 128314
rect 218244 128250 218296 128256
rect 218256 125594 218284 128250
rect 218244 125588 218296 125594
rect 218244 125530 218296 125536
rect 218428 125588 218480 125594
rect 218428 125530 218480 125536
rect 218440 119354 218468 125530
rect 218348 119326 218468 119354
rect 218348 109138 218376 119326
rect 218336 109132 218388 109138
rect 218336 109074 218388 109080
rect 218336 108996 218388 109002
rect 218336 108938 218388 108944
rect 218348 95198 218376 108938
rect 218336 95192 218388 95198
rect 218336 95134 218388 95140
rect 218336 85604 218388 85610
rect 218336 85546 218388 85552
rect 218348 71074 218376 85546
rect 218256 71046 218376 71074
rect 218256 64870 218284 71046
rect 218244 64864 218296 64870
rect 218244 64806 218296 64812
rect 218244 46980 218296 46986
rect 218244 46922 218296 46928
rect 218256 45558 218284 46922
rect 218244 45552 218296 45558
rect 218244 45494 218296 45500
rect 218336 45552 218388 45558
rect 218336 45494 218388 45500
rect 218348 37210 218376 45494
rect 219348 40180 219400 40186
rect 219348 40122 219400 40128
rect 219360 40089 219388 40122
rect 219346 40080 219402 40089
rect 219346 40015 219402 40024
rect 218256 37182 218376 37210
rect 218256 19446 218284 37182
rect 218244 19440 218296 19446
rect 218244 19382 218296 19388
rect 218244 19304 218296 19310
rect 218244 19246 218296 19252
rect 218256 8634 218284 19246
rect 218244 8628 218296 8634
rect 218244 8570 218296 8576
rect 218152 7268 218204 7274
rect 218152 7210 218204 7216
rect 218060 6044 218112 6050
rect 218060 5986 218112 5992
rect 219452 5982 219480 244038
rect 220188 239340 220216 244038
rect 219544 239312 220216 239340
rect 220820 239352 220872 239358
rect 219544 230489 219572 239312
rect 220820 239294 220872 239300
rect 219530 230480 219586 230489
rect 219530 230415 219586 230424
rect 219714 230480 219770 230489
rect 219714 230415 219770 230424
rect 219728 211177 219756 230415
rect 219530 211168 219586 211177
rect 219530 211103 219532 211112
rect 219584 211103 219586 211112
rect 219714 211168 219770 211177
rect 219714 211103 219770 211112
rect 219532 211074 219584 211080
rect 219624 211064 219676 211070
rect 219624 211006 219676 211012
rect 219636 188442 219664 211006
rect 219544 188414 219664 188442
rect 219544 183530 219572 188414
rect 219532 183524 219584 183530
rect 219532 183466 219584 183472
rect 219624 180056 219676 180062
rect 219624 179998 219676 180004
rect 219636 171086 219664 179998
rect 219624 171080 219676 171086
rect 219624 171022 219676 171028
rect 219532 162444 219584 162450
rect 219532 162386 219584 162392
rect 219544 160070 219572 162386
rect 219532 160064 219584 160070
rect 219532 160006 219584 160012
rect 219624 150476 219676 150482
rect 219624 150418 219676 150424
rect 219636 148458 219664 150418
rect 219636 148430 219756 148458
rect 219728 137714 219756 148430
rect 219636 137686 219756 137714
rect 219636 125610 219664 137686
rect 219544 125594 219664 125610
rect 219532 125588 219664 125594
rect 219584 125582 219664 125588
rect 219716 125588 219768 125594
rect 219532 125530 219584 125536
rect 219716 125530 219768 125536
rect 219728 119354 219756 125530
rect 219636 119326 219756 119354
rect 219636 109138 219664 119326
rect 219624 109132 219676 109138
rect 219624 109074 219676 109080
rect 219624 108996 219676 109002
rect 219624 108938 219676 108944
rect 219636 95198 219664 108938
rect 219624 95192 219676 95198
rect 219624 95134 219676 95140
rect 219624 85604 219676 85610
rect 219624 85546 219676 85552
rect 219636 70582 219664 85546
rect 219624 70576 219676 70582
rect 219624 70518 219676 70524
rect 219532 70372 219584 70378
rect 219532 70314 219584 70320
rect 219544 66230 219572 70314
rect 219532 66224 219584 66230
rect 219532 66166 219584 66172
rect 219532 46980 219584 46986
rect 219532 46922 219584 46928
rect 219544 45558 219572 46922
rect 219532 45552 219584 45558
rect 219532 45494 219584 45500
rect 219532 37256 219584 37262
rect 219532 37198 219584 37204
rect 219544 19446 219572 37198
rect 219532 19440 219584 19446
rect 219532 19382 219584 19388
rect 219532 19304 219584 19310
rect 219532 19246 219584 19252
rect 219544 7206 219572 19246
rect 219532 7200 219584 7206
rect 219532 7142 219584 7148
rect 219440 5976 219492 5982
rect 219440 5918 219492 5924
rect 220832 5914 220860 239294
rect 220924 8566 220952 244038
rect 221384 239358 221412 244038
rect 221372 239352 221424 239358
rect 221372 239294 221424 239300
rect 222200 239352 222252 239358
rect 222200 239294 222252 239300
rect 220912 8560 220964 8566
rect 220912 8502 220964 8508
rect 220820 5908 220872 5914
rect 220820 5850 220872 5856
rect 222212 5846 222240 239294
rect 222304 7138 222332 244052
rect 222672 244038 222962 244066
rect 223224 244038 223514 244066
rect 222672 236706 222700 244038
rect 223224 239358 223252 244038
rect 223212 239352 223264 239358
rect 223684 239340 223712 244174
rect 223212 239294 223264 239300
rect 223592 239312 223712 239340
rect 224420 244038 224802 244066
rect 224972 244038 225354 244066
rect 225708 244038 225998 244066
rect 226352 244038 226642 244066
rect 222476 236700 222528 236706
rect 222476 236642 222528 236648
rect 222660 236700 222712 236706
rect 222660 236642 222712 236648
rect 222488 231826 222516 236642
rect 222488 231798 222608 231826
rect 222580 215422 222608 231798
rect 222568 215416 222620 215422
rect 222568 215358 222620 215364
rect 222476 215280 222528 215286
rect 222476 215222 222528 215228
rect 222488 202910 222516 215222
rect 222476 202904 222528 202910
rect 222476 202846 222528 202852
rect 222568 202904 222620 202910
rect 222568 202846 222620 202852
rect 222580 201482 222608 202846
rect 222568 201476 222620 201482
rect 222568 201418 222620 201424
rect 222660 201476 222712 201482
rect 222660 201418 222712 201424
rect 222672 173942 222700 201418
rect 222476 173936 222528 173942
rect 222476 173878 222528 173884
rect 222660 173936 222712 173942
rect 222660 173878 222712 173884
rect 222488 169402 222516 173878
rect 222488 169374 222608 169402
rect 222580 159202 222608 169374
rect 222488 159174 222608 159202
rect 222488 154562 222516 159174
rect 222476 154556 222528 154562
rect 222476 154498 222528 154504
rect 222660 154556 222712 154562
rect 222660 154498 222712 154504
rect 222672 135289 222700 154498
rect 222474 135280 222530 135289
rect 222474 135215 222530 135224
rect 222658 135280 222714 135289
rect 222658 135215 222714 135224
rect 222488 125610 222516 135215
rect 222488 125582 222608 125610
rect 222580 118794 222608 125582
rect 222568 118788 222620 118794
rect 222568 118730 222620 118736
rect 222568 118652 222620 118658
rect 222568 118594 222620 118600
rect 222580 106282 222608 118594
rect 222476 106276 222528 106282
rect 222476 106218 222528 106224
rect 222568 106276 222620 106282
rect 222568 106218 222620 106224
rect 222488 104854 222516 106218
rect 222476 104848 222528 104854
rect 222476 104790 222528 104796
rect 222568 104780 222620 104786
rect 222568 104722 222620 104728
rect 222580 86970 222608 104722
rect 222476 86964 222528 86970
rect 222476 86906 222528 86912
rect 222568 86964 222620 86970
rect 222568 86906 222620 86912
rect 222488 82770 222516 86906
rect 222488 82742 222608 82770
rect 222580 67658 222608 82742
rect 222476 67652 222528 67658
rect 222476 67594 222528 67600
rect 222568 67652 222620 67658
rect 222568 67594 222620 67600
rect 222488 57882 222516 67594
rect 222396 57854 222516 57882
rect 222396 48362 222424 57854
rect 222396 48334 222516 48362
rect 222488 42090 222516 48334
rect 222476 42084 222528 42090
rect 222476 42026 222528 42032
rect 222660 29028 222712 29034
rect 222660 28970 222712 28976
rect 222672 14498 222700 28970
rect 222396 14470 222700 14498
rect 222396 8498 222424 14470
rect 222384 8492 222436 8498
rect 222384 8434 222436 8440
rect 222292 7132 222344 7138
rect 222292 7074 222344 7080
rect 223592 7070 223620 239312
rect 224420 236706 224448 244038
rect 223764 236700 223816 236706
rect 223764 236642 223816 236648
rect 224408 236700 224460 236706
rect 224408 236642 224460 236648
rect 223776 231849 223804 236642
rect 223762 231840 223818 231849
rect 223762 231775 223818 231784
rect 223946 231840 224002 231849
rect 223946 231775 224002 231784
rect 223960 230466 223988 231775
rect 223868 230438 223988 230466
rect 223868 222222 223896 230438
rect 223856 222216 223908 222222
rect 223856 222158 223908 222164
rect 223868 220862 223896 220893
rect 223856 220856 223908 220862
rect 223776 220804 223856 220810
rect 223776 220798 223908 220804
rect 223776 220782 223896 220798
rect 223776 211177 223804 220782
rect 223762 211168 223818 211177
rect 223762 211103 223818 211112
rect 223946 211168 224002 211177
rect 223946 211103 224002 211112
rect 223960 202910 223988 211103
rect 223856 202904 223908 202910
rect 223856 202846 223908 202852
rect 223948 202904 224000 202910
rect 223948 202846 224000 202852
rect 223868 196110 223896 202846
rect 223856 196104 223908 196110
rect 223856 196046 223908 196052
rect 223764 195968 223816 195974
rect 223764 195910 223816 195916
rect 223776 191826 223804 195910
rect 223764 191820 223816 191826
rect 223764 191762 223816 191768
rect 224040 191820 224092 191826
rect 224040 191762 224092 191768
rect 224052 182209 224080 191762
rect 223854 182200 223910 182209
rect 223854 182135 223910 182144
rect 224038 182200 224094 182209
rect 224038 182135 224094 182144
rect 223868 156890 223896 182135
rect 223776 156862 223896 156890
rect 223776 154562 223804 156862
rect 223764 154556 223816 154562
rect 223764 154498 223816 154504
rect 223948 154556 224000 154562
rect 223948 154498 224000 154504
rect 223960 135289 223988 154498
rect 223762 135280 223818 135289
rect 223762 135215 223818 135224
rect 223946 135280 224002 135289
rect 223946 135215 224002 135224
rect 223776 125610 223804 135215
rect 223776 125582 223896 125610
rect 223868 118794 223896 125582
rect 223856 118788 223908 118794
rect 223856 118730 223908 118736
rect 223856 118652 223908 118658
rect 223856 118594 223908 118600
rect 223868 106282 223896 118594
rect 223764 106276 223816 106282
rect 223764 106218 223816 106224
rect 223856 106276 223908 106282
rect 223856 106218 223908 106224
rect 223776 104854 223804 106218
rect 223764 104848 223816 104854
rect 223764 104790 223816 104796
rect 224040 95260 224092 95266
rect 224040 95202 224092 95208
rect 224052 87145 224080 95202
rect 224038 87136 224094 87145
rect 224038 87071 224094 87080
rect 223854 87000 223910 87009
rect 223764 86964 223816 86970
rect 223854 86935 223856 86944
rect 223764 86906 223816 86912
rect 223908 86935 223910 86944
rect 223856 86906 223908 86912
rect 223776 85542 223804 86906
rect 223764 85536 223816 85542
rect 223764 85478 223816 85484
rect 223764 74588 223816 74594
rect 223764 74530 223816 74536
rect 223776 64870 223804 74530
rect 223764 64864 223816 64870
rect 223764 64806 223816 64812
rect 223672 55276 223724 55282
rect 223672 55218 223724 55224
rect 223684 48362 223712 55218
rect 223684 48334 223804 48362
rect 223776 42090 223804 48334
rect 223764 42084 223816 42090
rect 223764 42026 223816 42032
rect 223764 29028 223816 29034
rect 223764 28970 223816 28976
rect 223776 27606 223804 28970
rect 223764 27600 223816 27606
rect 223764 27542 223816 27548
rect 223672 9716 223724 9722
rect 223672 9658 223724 9664
rect 223684 8430 223712 9658
rect 223672 8424 223724 8430
rect 223672 8366 223724 8372
rect 223580 7064 223632 7070
rect 223580 7006 223632 7012
rect 222200 5840 222252 5846
rect 222200 5782 222252 5788
rect 224972 5778 225000 244038
rect 225708 231878 225736 244038
rect 226248 242140 226300 242146
rect 226248 242082 226300 242088
rect 225052 231872 225104 231878
rect 225050 231840 225052 231849
rect 225696 231872 225748 231878
rect 225104 231840 225106 231849
rect 225050 231775 225106 231784
rect 225234 231840 225290 231849
rect 225696 231814 225748 231820
rect 225234 231775 225290 231784
rect 225248 230466 225276 231775
rect 225156 230438 225276 230466
rect 225156 222222 225184 230438
rect 225144 222216 225196 222222
rect 225144 222158 225196 222164
rect 225144 220856 225196 220862
rect 225142 220824 225144 220833
rect 225196 220824 225198 220833
rect 225142 220759 225198 220768
rect 225326 220824 225382 220833
rect 225326 220759 225382 220768
rect 225340 215914 225368 220759
rect 225156 215886 225368 215914
rect 225156 196058 225184 215886
rect 225064 196030 225184 196058
rect 225064 195922 225092 196030
rect 225064 195894 225184 195922
rect 225156 176610 225184 195894
rect 225064 176582 225184 176610
rect 225064 176338 225092 176582
rect 225064 176310 225184 176338
rect 225156 138122 225184 176310
rect 225064 138094 225184 138122
rect 225064 137714 225092 138094
rect 225064 137686 225184 137714
rect 225156 53122 225184 137686
rect 225064 53094 225184 53122
rect 225064 48278 225092 53094
rect 225052 48272 225104 48278
rect 225052 48214 225104 48220
rect 225144 48272 225196 48278
rect 225144 48214 225196 48220
rect 225156 7002 225184 48214
rect 225144 6996 225196 7002
rect 225144 6938 225196 6944
rect 224960 5772 225012 5778
rect 224960 5714 225012 5720
rect 214656 4140 214708 4146
rect 214656 4082 214708 4088
rect 215208 4140 215260 4146
rect 215208 4082 215260 4088
rect 222936 4140 222988 4146
rect 222936 4082 222988 4088
rect 213472 598 213868 626
rect 213472 480 213500 598
rect 214668 480 214696 4082
rect 220544 4072 220596 4078
rect 220544 4014 220596 4020
rect 219348 4004 219400 4010
rect 219348 3946 219400 3952
rect 215852 3936 215904 3942
rect 215852 3878 215904 3884
rect 215864 480 215892 3878
rect 217048 3188 217100 3194
rect 217048 3130 217100 3136
rect 217060 480 217088 3130
rect 218152 2848 218204 2854
rect 218152 2790 218204 2796
rect 218164 480 218192 2790
rect 219360 480 219388 3946
rect 220556 480 220584 4014
rect 221740 3120 221792 3126
rect 221740 3062 221792 3068
rect 221752 480 221780 3062
rect 222948 480 222976 4082
rect 226260 3670 226288 242082
rect 226352 4894 226380 244038
rect 226812 231878 226840 244174
rect 227838 244038 227944 244066
rect 226984 241732 227036 241738
rect 226984 241674 227036 241680
rect 226616 231872 226668 231878
rect 226616 231814 226668 231820
rect 226800 231872 226852 231878
rect 226800 231814 226852 231820
rect 226628 215370 226656 231814
rect 226536 215342 226656 215370
rect 226536 202910 226564 215342
rect 226524 202904 226576 202910
rect 226524 202846 226576 202852
rect 226616 202904 226668 202910
rect 226616 202846 226668 202852
rect 226628 201482 226656 202846
rect 226616 201476 226668 201482
rect 226616 201418 226668 201424
rect 226800 201476 226852 201482
rect 226800 201418 226852 201424
rect 226812 200122 226840 201418
rect 226708 200116 226760 200122
rect 226708 200058 226760 200064
rect 226800 200116 226852 200122
rect 226800 200058 226852 200064
rect 226720 190641 226748 200058
rect 226706 190632 226762 190641
rect 226706 190567 226762 190576
rect 226430 190496 226486 190505
rect 226430 190431 226432 190440
rect 226484 190431 226486 190440
rect 226800 190460 226852 190466
rect 226432 190402 226484 190408
rect 226800 190402 226852 190408
rect 226812 180849 226840 190402
rect 226614 180840 226670 180849
rect 226614 180775 226670 180784
rect 226798 180840 226854 180849
rect 226798 180775 226854 180784
rect 226628 174010 226656 180775
rect 226616 174004 226668 174010
rect 226616 173946 226668 173952
rect 226524 173868 226576 173874
rect 226524 173810 226576 173816
rect 226536 154737 226564 173810
rect 226522 154728 226578 154737
rect 226522 154663 226578 154672
rect 226522 154592 226578 154601
rect 226522 154527 226524 154536
rect 226576 154527 226578 154536
rect 226616 154556 226668 154562
rect 226524 154498 226576 154504
rect 226616 154498 226668 154504
rect 226628 144922 226656 154498
rect 226628 144894 226748 144922
rect 226720 135289 226748 144894
rect 226522 135280 226578 135289
rect 226522 135215 226578 135224
rect 226706 135280 226762 135289
rect 226706 135215 226762 135224
rect 226536 125610 226564 135215
rect 226536 125582 226656 125610
rect 226628 93838 226656 125582
rect 226616 93832 226668 93838
rect 226616 93774 226668 93780
rect 226616 92540 226668 92546
rect 226616 92482 226668 92488
rect 226628 82822 226656 92482
rect 226616 82816 226668 82822
rect 226616 82758 226668 82764
rect 226708 55276 226760 55282
rect 226708 55218 226760 55224
rect 226720 38706 226748 55218
rect 226628 38678 226748 38706
rect 226628 38604 226656 38678
rect 226536 38576 226656 38604
rect 226536 27554 226564 38576
rect 226536 27526 226656 27554
rect 226628 18034 226656 27526
rect 226536 18006 226656 18034
rect 226536 5710 226564 18006
rect 226524 5704 226576 5710
rect 226524 5646 226576 5652
rect 226340 4888 226392 4894
rect 226340 4830 226392 4836
rect 225328 3664 225380 3670
rect 225328 3606 225380 3612
rect 226248 3664 226300 3670
rect 226248 3606 226300 3612
rect 224132 3188 224184 3194
rect 224132 3130 224184 3136
rect 224144 480 224172 3130
rect 225340 480 225368 3606
rect 226996 3058 227024 241674
rect 227812 239352 227864 239358
rect 227812 239294 227864 239300
rect 227824 6186 227852 239294
rect 227812 6180 227864 6186
rect 227812 6122 227864 6128
rect 227916 4826 227944 244038
rect 228468 242010 228496 244052
rect 228744 244038 229034 244066
rect 228456 242004 228508 242010
rect 228456 241946 228508 241952
rect 228744 239358 228772 244038
rect 228732 239352 228784 239358
rect 229204 239306 229232 244174
rect 228732 239294 228784 239300
rect 229112 239278 229232 239306
rect 229006 40352 229062 40361
rect 229006 40287 229062 40296
rect 229020 39817 229048 40287
rect 229006 39808 229062 39817
rect 229006 39743 229062 39752
rect 229112 4962 229140 239278
rect 229848 231878 229876 244174
rect 230584 244038 230874 244066
rect 231136 244038 231518 244066
rect 231964 244038 232070 244066
rect 232424 244038 232714 244066
rect 233358 244038 233464 244066
rect 230480 239352 230532 239358
rect 230480 239294 230532 239300
rect 229376 231872 229428 231878
rect 229376 231814 229428 231820
rect 229836 231872 229888 231878
rect 229836 231814 229888 231820
rect 229388 215370 229416 231814
rect 229296 215342 229416 215370
rect 229296 202910 229324 215342
rect 229284 202904 229336 202910
rect 229284 202846 229336 202852
rect 229376 202904 229428 202910
rect 229376 202846 229428 202852
rect 229388 201482 229416 202846
rect 229376 201476 229428 201482
rect 229376 201418 229428 201424
rect 229468 201476 229520 201482
rect 229468 201418 229520 201424
rect 229480 173942 229508 201418
rect 229284 173936 229336 173942
rect 229284 173878 229336 173884
rect 229468 173936 229520 173942
rect 229468 173878 229520 173884
rect 229296 157570 229324 173878
rect 229204 157542 229324 157570
rect 229204 154630 229232 157542
rect 229192 154624 229244 154630
rect 229192 154566 229244 154572
rect 229284 154624 229336 154630
rect 229284 154566 229336 154572
rect 229296 149682 229324 154566
rect 229296 149654 229508 149682
rect 229480 135289 229508 149654
rect 229282 135280 229338 135289
rect 229282 135215 229338 135224
rect 229466 135280 229522 135289
rect 229466 135215 229522 135224
rect 229296 125610 229324 135215
rect 229296 125582 229416 125610
rect 229388 101402 229416 125582
rect 229296 101374 229416 101402
rect 229296 87038 229324 101374
rect 229192 87032 229244 87038
rect 229192 86974 229244 86980
rect 229284 87032 229336 87038
rect 229284 86974 229336 86980
rect 229204 85542 229232 86974
rect 229192 85536 229244 85542
rect 229192 85478 229244 85484
rect 229376 85468 229428 85474
rect 229376 85410 229428 85416
rect 229388 58002 229416 85410
rect 229284 57996 229336 58002
rect 229284 57938 229336 57944
rect 229376 57996 229428 58002
rect 229376 57938 229428 57944
rect 229296 53258 229324 57938
rect 229296 53230 229508 53258
rect 229480 39794 229508 53230
rect 229388 39766 229508 39794
rect 229388 38604 229416 39766
rect 229388 38576 229508 38604
rect 229480 29034 229508 38576
rect 229376 29028 229428 29034
rect 229376 28970 229428 28976
rect 229468 29028 229520 29034
rect 229468 28970 229520 28976
rect 229388 19378 229416 28970
rect 229284 19372 229336 19378
rect 229284 19314 229336 19320
rect 229376 19372 229428 19378
rect 229376 19314 229428 19320
rect 229296 8362 229324 19314
rect 229284 8356 229336 8362
rect 229284 8298 229336 8304
rect 230492 5030 230520 239294
rect 230584 6254 230612 244038
rect 231136 239358 231164 244038
rect 231768 242004 231820 242010
rect 231768 241946 231820 241952
rect 231124 239352 231176 239358
rect 231124 239294 231176 239300
rect 230572 6248 230624 6254
rect 230572 6190 230624 6196
rect 230480 5024 230532 5030
rect 230480 4966 230532 4972
rect 229100 4956 229152 4962
rect 229100 4898 229152 4904
rect 227904 4820 227956 4826
rect 227904 4762 227956 4768
rect 231780 3670 231808 241946
rect 231860 239352 231912 239358
rect 231860 239294 231912 239300
rect 231872 6390 231900 239294
rect 231860 6384 231912 6390
rect 231860 6326 231912 6332
rect 231964 6322 231992 244038
rect 232424 239358 232452 244038
rect 232504 241936 232556 241942
rect 232504 241878 232556 241884
rect 232412 239352 232464 239358
rect 232412 239294 232464 239300
rect 231952 6316 232004 6322
rect 231952 6258 232004 6264
rect 228916 3664 228968 3670
rect 231216 3664 231268 3670
rect 228916 3606 228968 3612
rect 231214 3632 231216 3641
rect 231308 3664 231360 3670
rect 231268 3632 231270 3641
rect 226984 3052 227036 3058
rect 226984 2994 227036 3000
rect 226524 2984 226576 2990
rect 226524 2926 226576 2932
rect 226536 480 226564 2926
rect 227720 2916 227772 2922
rect 227720 2858 227772 2864
rect 227732 480 227760 2858
rect 228928 480 228956 3606
rect 231308 3606 231360 3612
rect 231768 3664 231820 3670
rect 232516 3641 232544 241878
rect 233332 239352 233384 239358
rect 233332 239294 233384 239300
rect 233240 236700 233292 236706
rect 233240 236642 233292 236648
rect 233252 5098 233280 236642
rect 233344 5642 233372 239294
rect 233436 7614 233464 244038
rect 233528 244038 233910 244066
rect 234264 244038 234554 244066
rect 233528 236706 233556 244038
rect 234264 239358 234292 244038
rect 234252 239352 234304 239358
rect 234724 239340 234752 244174
rect 234252 239294 234304 239300
rect 234632 239312 234752 239340
rect 235460 244038 235750 244066
rect 236104 244038 236394 244066
rect 233516 236700 233568 236706
rect 233516 236642 233568 236648
rect 233424 7608 233476 7614
rect 233424 7550 233476 7556
rect 233332 5636 233384 5642
rect 233332 5578 233384 5584
rect 233240 5092 233292 5098
rect 233240 5034 233292 5040
rect 233700 4820 233752 4826
rect 233700 4762 233752 4768
rect 231768 3606 231820 3612
rect 232502 3632 232558 3641
rect 231214 3567 231270 3576
rect 230112 3052 230164 3058
rect 230112 2994 230164 3000
rect 230124 480 230152 2994
rect 231320 480 231348 3606
rect 232502 3567 232558 3576
rect 232504 2916 232556 2922
rect 232504 2858 232556 2864
rect 232516 480 232544 2858
rect 233712 480 233740 4762
rect 234632 3466 234660 239312
rect 235460 231878 235488 244038
rect 234896 231872 234948 231878
rect 234896 231814 234948 231820
rect 235448 231872 235500 231878
rect 235448 231814 235500 231820
rect 234908 215370 234936 231814
rect 234816 215342 234936 215370
rect 234816 207754 234844 215342
rect 234816 207726 234936 207754
rect 234908 193322 234936 207726
rect 234896 193316 234948 193322
rect 234896 193258 234948 193264
rect 234804 193248 234856 193254
rect 234802 193216 234804 193225
rect 234856 193216 234858 193225
rect 234802 193151 234858 193160
rect 234986 193216 235042 193225
rect 234986 193151 235042 193160
rect 235000 162897 235028 193151
rect 234802 162888 234858 162897
rect 234802 162823 234858 162832
rect 234986 162888 235042 162897
rect 234986 162823 235042 162832
rect 234816 147506 234844 162823
rect 234816 147478 234936 147506
rect 234908 144906 234936 147478
rect 234896 144900 234948 144906
rect 234896 144842 234948 144848
rect 234988 144900 235040 144906
rect 234988 144842 235040 144848
rect 235000 135289 235028 144842
rect 234802 135280 234858 135289
rect 234802 135215 234804 135224
rect 234856 135215 234858 135224
rect 234986 135280 235042 135289
rect 234986 135215 234988 135224
rect 234804 135186 234856 135192
rect 235040 135215 235042 135224
rect 234988 135186 235040 135192
rect 235000 133890 235028 135186
rect 234988 133884 235040 133890
rect 234988 133826 235040 133832
rect 234804 124296 234856 124302
rect 234804 124238 234856 124244
rect 234816 124166 234844 124238
rect 234804 124160 234856 124166
rect 234804 124102 234856 124108
rect 234804 114572 234856 114578
rect 234804 114514 234856 114520
rect 234816 106298 234844 114514
rect 234816 106270 234936 106298
rect 234908 101402 234936 106270
rect 234816 101374 234936 101402
rect 234816 87145 234844 101374
rect 234802 87136 234858 87145
rect 234802 87071 234858 87080
rect 234710 87000 234766 87009
rect 234710 86935 234766 86944
rect 234724 77314 234752 86935
rect 234712 77308 234764 77314
rect 234712 77250 234764 77256
rect 234804 77308 234856 77314
rect 234804 77250 234856 77256
rect 234816 50946 234844 77250
rect 234816 50918 234936 50946
rect 234908 48278 234936 50918
rect 234896 48272 234948 48278
rect 234896 48214 234948 48220
rect 234804 38684 234856 38690
rect 234804 38626 234856 38632
rect 234816 33810 234844 38626
rect 234724 33782 234844 33810
rect 234724 19378 234752 33782
rect 234712 19372 234764 19378
rect 234712 19314 234764 19320
rect 234804 19372 234856 19378
rect 234804 19314 234856 19320
rect 234816 5166 234844 19314
rect 236104 5574 236132 244038
rect 236564 231878 236592 244174
rect 237392 244038 237590 244066
rect 236368 231872 236420 231878
rect 236368 231814 236420 231820
rect 236552 231872 236604 231878
rect 236552 231814 236604 231820
rect 236380 215370 236408 231814
rect 236288 215342 236408 215370
rect 236288 205578 236316 215342
rect 236288 205550 236408 205578
rect 236380 198098 236408 205550
rect 236380 198070 236500 198098
rect 236472 193254 236500 198070
rect 236276 193248 236328 193254
rect 236276 193190 236328 193196
rect 236460 193248 236512 193254
rect 236460 193190 236512 193196
rect 236288 188442 236316 193190
rect 236288 188414 236408 188442
rect 236380 178786 236408 188414
rect 236380 178758 236500 178786
rect 236472 173942 236500 178758
rect 236276 173936 236328 173942
rect 236276 173878 236328 173884
rect 236460 173936 236512 173942
rect 236460 173878 236512 173884
rect 236288 164218 236316 173878
rect 236276 164212 236328 164218
rect 236276 164154 236328 164160
rect 236276 157276 236328 157282
rect 236276 157218 236328 157224
rect 236288 149682 236316 157218
rect 236288 149654 236408 149682
rect 236380 144906 236408 149654
rect 236276 144900 236328 144906
rect 236276 144842 236328 144848
rect 236368 144900 236420 144906
rect 236368 144842 236420 144848
rect 236288 130370 236316 144842
rect 236288 130342 236408 130370
rect 236380 116113 236408 130342
rect 236366 116104 236422 116113
rect 236366 116039 236422 116048
rect 236274 115968 236330 115977
rect 236274 115903 236276 115912
rect 236328 115903 236330 115912
rect 236276 115874 236328 115880
rect 236368 115864 236420 115870
rect 236368 115806 236420 115812
rect 236380 101402 236408 115806
rect 236288 101374 236408 101402
rect 236288 87038 236316 101374
rect 236184 87032 236236 87038
rect 236184 86974 236236 86980
rect 236276 87032 236328 87038
rect 236276 86974 236328 86980
rect 236196 77314 236224 86974
rect 236184 77308 236236 77314
rect 236184 77250 236236 77256
rect 236276 77308 236328 77314
rect 236276 77250 236328 77256
rect 236288 67590 236316 77250
rect 236276 67584 236328 67590
rect 236276 67526 236328 67532
rect 236368 67584 236420 67590
rect 236368 67526 236420 67532
rect 236380 48278 236408 67526
rect 236276 48272 236328 48278
rect 236276 48214 236328 48220
rect 236368 48272 236420 48278
rect 236368 48214 236420 48220
rect 236288 29102 236316 48214
rect 236276 29096 236328 29102
rect 236276 29038 236328 29044
rect 236184 29028 236236 29034
rect 236184 28970 236236 28976
rect 236196 19378 236224 28970
rect 236184 19372 236236 19378
rect 236184 19314 236236 19320
rect 236276 19372 236328 19378
rect 236276 19314 236328 19320
rect 236092 5568 236144 5574
rect 236092 5510 236144 5516
rect 234804 5160 234856 5166
rect 234804 5102 234856 5108
rect 236000 3664 236052 3670
rect 236000 3606 236052 3612
rect 234620 3460 234672 3466
rect 234620 3402 234672 3408
rect 234804 3460 234856 3466
rect 234804 3402 234856 3408
rect 234816 480 234844 3402
rect 236012 480 236040 3606
rect 236288 3602 236316 19314
rect 237392 5234 237420 244038
rect 237760 239426 237788 244174
rect 238772 244038 238878 244066
rect 239140 244038 239430 244066
rect 239692 244038 240074 244066
rect 240244 244038 240626 244066
rect 238668 241528 238720 241534
rect 238668 241470 238720 241476
rect 238680 240145 238708 241470
rect 238482 240136 238538 240145
rect 238482 240071 238538 240080
rect 238666 240136 238722 240145
rect 238666 240071 238722 240080
rect 237748 239420 237800 239426
rect 237748 239362 237800 239368
rect 237656 231872 237708 231878
rect 237656 231814 237708 231820
rect 237668 215370 237696 231814
rect 238496 230518 238524 240071
rect 238484 230512 238536 230518
rect 238484 230454 238536 230460
rect 238668 230512 238720 230518
rect 238668 230454 238720 230460
rect 238680 220833 238708 230454
rect 238482 220824 238538 220833
rect 238482 220759 238538 220768
rect 238666 220824 238722 220833
rect 238666 220759 238722 220768
rect 237576 215342 237696 215370
rect 237576 207754 237604 215342
rect 238496 211177 238524 220759
rect 238482 211168 238538 211177
rect 238482 211103 238538 211112
rect 238666 211168 238722 211177
rect 238666 211103 238722 211112
rect 237576 207726 237696 207754
rect 237668 198098 237696 207726
rect 238680 206310 238708 211103
rect 238484 206304 238536 206310
rect 238484 206246 238536 206252
rect 238668 206304 238720 206310
rect 238668 206246 238720 206252
rect 238496 201521 238524 206246
rect 238482 201512 238538 201521
rect 238482 201447 238484 201456
rect 238536 201447 238538 201456
rect 238666 201512 238722 201521
rect 238666 201447 238668 201456
rect 238484 201418 238536 201424
rect 238720 201447 238722 201456
rect 238668 201418 238720 201424
rect 237668 198070 237788 198098
rect 237760 193254 237788 198070
rect 237564 193248 237616 193254
rect 237748 193248 237800 193254
rect 237616 193196 237696 193202
rect 237564 193190 237696 193196
rect 237748 193190 237800 193196
rect 237576 193174 237696 193190
rect 237668 178786 237696 193174
rect 238496 183598 238524 201418
rect 238484 183592 238536 183598
rect 238484 183534 238536 183540
rect 238668 183592 238720 183598
rect 238668 183534 238720 183540
rect 238680 182170 238708 183534
rect 238668 182164 238720 182170
rect 238668 182106 238720 182112
rect 237668 178758 237788 178786
rect 237760 173942 237788 178758
rect 237564 173936 237616 173942
rect 237564 173878 237616 173884
rect 237748 173936 237800 173942
rect 237748 173878 237800 173884
rect 237576 164218 237604 173878
rect 238484 172576 238536 172582
rect 238484 172518 238536 172524
rect 238496 164286 238524 172518
rect 238484 164280 238536 164286
rect 238484 164222 238536 164228
rect 238668 164280 238720 164286
rect 238668 164222 238720 164228
rect 237564 164212 237616 164218
rect 237564 164154 237616 164160
rect 238680 162858 238708 164222
rect 238392 162852 238444 162858
rect 238392 162794 238444 162800
rect 238668 162852 238720 162858
rect 238668 162794 238720 162800
rect 237564 157276 237616 157282
rect 237564 157218 237616 157224
rect 237576 149682 237604 157218
rect 238404 153241 238432 162794
rect 238390 153232 238446 153241
rect 238390 153167 238446 153176
rect 238574 153232 238630 153241
rect 238574 153167 238630 153176
rect 237576 149654 237696 149682
rect 237668 144906 237696 149654
rect 238588 144974 238616 153167
rect 238576 144968 238628 144974
rect 238576 144910 238628 144916
rect 238668 144968 238720 144974
rect 238668 144910 238720 144916
rect 237564 144900 237616 144906
rect 237564 144842 237616 144848
rect 237656 144900 237708 144906
rect 237656 144842 237708 144848
rect 237576 130370 237604 144842
rect 238680 143546 238708 144910
rect 238668 143540 238720 143546
rect 238668 143482 238720 143488
rect 237576 130342 237696 130370
rect 237668 116113 237696 130342
rect 238668 125656 238720 125662
rect 238668 125598 238720 125604
rect 238680 124166 238708 125598
rect 238668 124160 238720 124166
rect 238668 124102 238720 124108
rect 237654 116104 237710 116113
rect 237654 116039 237710 116048
rect 237562 115968 237618 115977
rect 237562 115903 237564 115912
rect 237616 115903 237618 115912
rect 237564 115874 237616 115880
rect 237656 115864 237708 115870
rect 237656 115806 237708 115812
rect 237668 101402 237696 115806
rect 238576 114572 238628 114578
rect 238576 114514 238628 114520
rect 238588 106350 238616 114514
rect 238576 106344 238628 106350
rect 238576 106286 238628 106292
rect 238668 106344 238720 106350
rect 238668 106286 238720 106292
rect 238680 104854 238708 106286
rect 238668 104848 238720 104854
rect 238668 104790 238720 104796
rect 237576 101374 237696 101402
rect 237576 87145 237604 101374
rect 238668 95260 238720 95266
rect 238668 95202 238720 95208
rect 237562 87136 237618 87145
rect 237562 87071 237618 87080
rect 237470 87000 237526 87009
rect 237470 86935 237526 86944
rect 237484 77314 237512 86935
rect 238680 85542 238708 95202
rect 238668 85536 238720 85542
rect 238668 85478 238720 85484
rect 237472 77308 237524 77314
rect 237472 77250 237524 77256
rect 237564 77308 237616 77314
rect 237564 77250 237616 77256
rect 237576 67590 237604 77250
rect 238668 75948 238720 75954
rect 238668 75890 238720 75896
rect 237564 67584 237616 67590
rect 237564 67526 237616 67532
rect 237656 67584 237708 67590
rect 237656 67526 237708 67532
rect 237668 48278 237696 67526
rect 238680 66230 238708 75890
rect 238668 66224 238720 66230
rect 238668 66166 238720 66172
rect 238668 48340 238720 48346
rect 238668 48282 238720 48288
rect 237564 48272 237616 48278
rect 237564 48214 237616 48220
rect 237656 48272 237708 48278
rect 237656 48214 237708 48220
rect 237576 33810 237604 48214
rect 238680 46918 238708 48282
rect 238668 46912 238720 46918
rect 238668 46854 238720 46860
rect 238666 40624 238722 40633
rect 238666 40559 238722 40568
rect 238680 40089 238708 40559
rect 238666 40080 238722 40089
rect 238666 40015 238722 40024
rect 238668 37324 238720 37330
rect 238668 37266 238720 37272
rect 237484 33782 237604 33810
rect 237484 19378 237512 33782
rect 238680 29034 238708 37266
rect 238668 29028 238720 29034
rect 238668 28970 238720 28976
rect 238668 27736 238720 27742
rect 238668 27678 238720 27684
rect 238680 27606 238708 27678
rect 238668 27600 238720 27606
rect 238668 27542 238720 27548
rect 237472 19372 237524 19378
rect 237472 19314 237524 19320
rect 237564 19372 237616 19378
rect 237564 19314 237616 19320
rect 237576 6458 237604 19314
rect 238576 9716 238628 9722
rect 238576 9658 238628 9664
rect 237564 6452 237616 6458
rect 237564 6394 237616 6400
rect 237380 5228 237432 5234
rect 237380 5170 237432 5176
rect 237196 4888 237248 4894
rect 237196 4830 237248 4836
rect 236276 3596 236328 3602
rect 236276 3538 236328 3544
rect 237208 480 237236 4830
rect 238588 610 238616 9658
rect 238772 3738 238800 244038
rect 239140 239442 239168 244038
rect 238864 239414 239168 239442
rect 238864 5302 238892 239414
rect 239692 231878 239720 244038
rect 239128 231872 239180 231878
rect 239128 231814 239180 231820
rect 239680 231872 239732 231878
rect 239680 231814 239732 231820
rect 239140 215370 239168 231814
rect 239048 215342 239168 215370
rect 239048 205578 239076 215342
rect 239048 205550 239168 205578
rect 239140 198098 239168 205550
rect 239140 198070 239260 198098
rect 239232 193254 239260 198070
rect 239036 193248 239088 193254
rect 239034 193216 239036 193225
rect 239220 193248 239272 193254
rect 239088 193216 239090 193225
rect 239034 193151 239090 193160
rect 239218 193216 239220 193225
rect 239272 193216 239274 193225
rect 239218 193151 239274 193160
rect 239232 186266 239260 193151
rect 239140 186238 239260 186266
rect 239140 178786 239168 186238
rect 239140 178758 239260 178786
rect 239232 173942 239260 178758
rect 239036 173936 239088 173942
rect 239036 173878 239088 173884
rect 239220 173936 239272 173942
rect 239220 173878 239272 173884
rect 239048 164218 239076 173878
rect 239036 164212 239088 164218
rect 239036 164154 239088 164160
rect 239128 164212 239180 164218
rect 239128 164154 239180 164160
rect 239140 159202 239168 164154
rect 239048 159174 239168 159202
rect 239048 154562 239076 159174
rect 239036 154556 239088 154562
rect 239036 154498 239088 154504
rect 239128 154488 239180 154494
rect 239128 154430 239180 154436
rect 239140 144906 239168 154430
rect 239036 144900 239088 144906
rect 239036 144842 239088 144848
rect 239128 144900 239180 144906
rect 239128 144842 239180 144848
rect 239048 130370 239076 144842
rect 239048 130342 239260 130370
rect 239232 128330 239260 130342
rect 239140 128302 239260 128330
rect 239140 125594 239168 128302
rect 238944 125588 238996 125594
rect 238944 125530 238996 125536
rect 239128 125588 239180 125594
rect 239128 125530 239180 125536
rect 238956 118674 238984 125530
rect 238956 118646 239076 118674
rect 239048 111058 239076 118646
rect 239048 111030 239168 111058
rect 239140 101402 239168 111030
rect 239048 101374 239168 101402
rect 239048 50946 239076 101374
rect 239048 50918 239168 50946
rect 239140 19378 239168 50918
rect 240046 40624 240102 40633
rect 240046 40559 240102 40568
rect 240060 40361 240088 40559
rect 240046 40352 240102 40361
rect 240046 40287 240102 40296
rect 239036 19372 239088 19378
rect 239036 19314 239088 19320
rect 239128 19372 239180 19378
rect 239128 19314 239180 19320
rect 239048 6526 239076 19314
rect 239036 6520 239088 6526
rect 239036 6462 239088 6468
rect 238852 5296 238904 5302
rect 238852 5238 238904 5244
rect 240244 3806 240272 244038
rect 241256 241874 241284 244052
rect 241624 244038 241914 244066
rect 242176 244038 242466 244066
rect 243004 244038 243110 244066
rect 241244 241868 241296 241874
rect 241244 241810 241296 241816
rect 241428 241868 241480 241874
rect 241428 241810 241480 241816
rect 241440 3806 241468 241810
rect 241520 239352 241572 239358
rect 241520 239294 241572 239300
rect 240232 3800 240284 3806
rect 240232 3742 240284 3748
rect 240784 3800 240836 3806
rect 240784 3742 240836 3748
rect 241428 3800 241480 3806
rect 241428 3742 241480 3748
rect 238760 3732 238812 3738
rect 238760 3674 238812 3680
rect 239588 3528 239640 3534
rect 239588 3470 239640 3476
rect 238392 604 238444 610
rect 238392 546 238444 552
rect 238576 604 238628 610
rect 238576 546 238628 552
rect 238404 480 238432 546
rect 239600 480 239628 3470
rect 240796 480 240824 3742
rect 241532 3602 241560 239294
rect 241624 6594 241652 244038
rect 242176 239358 242204 244038
rect 242164 239352 242216 239358
rect 242164 239294 242216 239300
rect 241612 6588 241664 6594
rect 241612 6530 241664 6536
rect 243004 5370 243032 244038
rect 243740 242078 243768 244052
rect 244306 244038 244504 244066
rect 243728 242072 243780 242078
rect 243728 242014 243780 242020
rect 244188 242072 244240 242078
rect 244188 242014 244240 242020
rect 243544 241664 243596 241670
rect 243544 241606 243596 241612
rect 242992 5364 243044 5370
rect 242992 5306 243044 5312
rect 243176 3800 243228 3806
rect 243176 3742 243228 3748
rect 241520 3596 241572 3602
rect 241520 3538 241572 3544
rect 241980 3596 242032 3602
rect 241980 3538 242032 3544
rect 241992 480 242020 3538
rect 243188 480 243216 3742
rect 243556 3670 243584 241606
rect 244200 3806 244228 242014
rect 244372 239352 244424 239358
rect 244372 239294 244424 239300
rect 244384 5438 244412 239294
rect 244372 5432 244424 5438
rect 244372 5374 244424 5380
rect 244188 3800 244240 3806
rect 244188 3742 244240 3748
rect 244476 3738 244504 244038
rect 244568 244038 244950 244066
rect 244568 239358 244596 244038
rect 245580 242758 245608 244052
rect 245568 242752 245620 242758
rect 245568 242694 245620 242700
rect 245660 242752 245712 242758
rect 245660 242694 245712 242700
rect 245672 242570 245700 242694
rect 245580 242542 245700 242570
rect 244556 239352 244608 239358
rect 244556 239294 244608 239300
rect 244464 3732 244516 3738
rect 244464 3674 244516 3680
rect 243544 3664 243596 3670
rect 243544 3606 243596 3612
rect 244372 3256 244424 3262
rect 244372 3198 244424 3204
rect 244384 480 244412 3198
rect 245580 480 245608 242542
rect 245764 239306 245792 244174
rect 245672 239278 245792 239306
rect 246500 244038 246790 244066
rect 245672 5506 245700 239278
rect 246500 234666 246528 244038
rect 247420 242486 247448 244052
rect 247788 244038 247986 244066
rect 248524 244038 248630 244066
rect 247408 242480 247460 242486
rect 247408 242422 247460 242428
rect 247788 239358 247816 244038
rect 248328 242480 248380 242486
rect 248328 242422 248380 242428
rect 248340 240122 248368 242422
rect 248248 240094 248368 240122
rect 247224 239352 247276 239358
rect 247224 239294 247276 239300
rect 247776 239352 247828 239358
rect 247776 239294 247828 239300
rect 245936 234660 245988 234666
rect 245936 234602 245988 234608
rect 246488 234660 246540 234666
rect 246488 234602 246540 234608
rect 245948 225078 245976 234602
rect 245936 225072 245988 225078
rect 245936 225014 245988 225020
rect 247236 225010 247264 239294
rect 248248 230518 248276 240094
rect 248144 230512 248196 230518
rect 247958 230480 248014 230489
rect 247958 230415 248014 230424
rect 248142 230480 248144 230489
rect 248236 230512 248288 230518
rect 248196 230480 248198 230489
rect 248236 230454 248288 230460
rect 248142 230415 248198 230424
rect 247224 225004 247276 225010
rect 247224 224946 247276 224952
rect 245844 224936 245896 224942
rect 245844 224878 245896 224884
rect 245856 222154 245884 224878
rect 247316 224868 247368 224874
rect 247316 224810 247368 224816
rect 247328 222170 247356 224810
rect 245844 222148 245896 222154
rect 247328 222142 247448 222170
rect 245844 222090 245896 222096
rect 245936 222012 245988 222018
rect 245936 221954 245988 221960
rect 245948 205578 245976 221954
rect 247420 212566 247448 222142
rect 247972 220862 248000 230415
rect 248340 220862 248368 220893
rect 247960 220856 248012 220862
rect 248328 220856 248380 220862
rect 247960 220798 248012 220804
rect 248248 220804 248328 220810
rect 248248 220798 248380 220804
rect 248248 220782 248368 220798
rect 247316 212560 247368 212566
rect 247316 212502 247368 212508
rect 247408 212560 247460 212566
rect 247408 212502 247460 212508
rect 247328 205578 247356 212502
rect 248248 211206 248276 220782
rect 248144 211200 248196 211206
rect 248144 211142 248196 211148
rect 248236 211200 248288 211206
rect 248236 211142 248288 211148
rect 245856 205550 245976 205578
rect 247236 205550 247356 205578
rect 245856 202881 245884 205550
rect 247236 202881 247264 205550
rect 248156 202910 248184 211142
rect 248144 202904 248196 202910
rect 245842 202872 245898 202881
rect 245842 202807 245898 202816
rect 246118 202872 246174 202881
rect 246118 202807 246174 202816
rect 247038 202872 247094 202881
rect 247038 202807 247094 202816
rect 247222 202872 247278 202881
rect 248144 202846 248196 202852
rect 248328 202904 248380 202910
rect 248328 202846 248380 202852
rect 247222 202807 247278 202816
rect 246132 193254 246160 202807
rect 247052 193254 247080 202807
rect 248340 201482 248368 202846
rect 248328 201476 248380 201482
rect 248328 201418 248380 201424
rect 245936 193248 245988 193254
rect 245936 193190 245988 193196
rect 246120 193248 246172 193254
rect 246120 193190 246172 193196
rect 247040 193248 247092 193254
rect 247040 193190 247092 193196
rect 247316 193248 247368 193254
rect 247316 193190 247368 193196
rect 245948 186266 245976 193190
rect 247328 186266 247356 193190
rect 248144 191888 248196 191894
rect 248144 191830 248196 191836
rect 245856 186238 245976 186266
rect 247236 186238 247356 186266
rect 245856 183569 245884 186238
rect 247236 183569 247264 186238
rect 248156 183598 248184 191830
rect 248144 183592 248196 183598
rect 245842 183560 245898 183569
rect 245842 183495 245898 183504
rect 246118 183560 246174 183569
rect 246118 183495 246174 183504
rect 247038 183560 247094 183569
rect 247038 183495 247094 183504
rect 247222 183560 247278 183569
rect 248144 183534 248196 183540
rect 248328 183592 248380 183598
rect 248328 183534 248380 183540
rect 247222 183495 247278 183504
rect 246132 173942 246160 183495
rect 247052 173942 247080 183495
rect 248340 182170 248368 183534
rect 248144 182164 248196 182170
rect 248144 182106 248196 182112
rect 248328 182164 248380 182170
rect 248328 182106 248380 182112
rect 245936 173936 245988 173942
rect 245936 173878 245988 173884
rect 246120 173936 246172 173942
rect 246120 173878 246172 173884
rect 247040 173936 247092 173942
rect 247040 173878 247092 173884
rect 247316 173936 247368 173942
rect 247316 173878 247368 173884
rect 245948 166954 245976 173878
rect 247328 166954 247356 173878
rect 248156 172553 248184 182106
rect 248142 172544 248198 172553
rect 248142 172479 248198 172488
rect 248326 172544 248382 172553
rect 248326 172479 248382 172488
rect 245856 166926 245976 166954
rect 247236 166926 247356 166954
rect 245856 154442 245884 166926
rect 247236 164218 247264 166926
rect 247040 164212 247092 164218
rect 247040 164154 247092 164160
rect 247224 164212 247276 164218
rect 247224 164154 247276 164160
rect 247052 154601 247080 164154
rect 248340 162858 248368 172479
rect 248328 162852 248380 162858
rect 248328 162794 248380 162800
rect 247038 154592 247094 154601
rect 247038 154527 247094 154536
rect 247314 154592 247370 154601
rect 247314 154527 247370 154536
rect 245764 154414 245884 154442
rect 245764 143546 245792 154414
rect 247328 147642 247356 154527
rect 248328 153264 248380 153270
rect 248328 153206 248380 153212
rect 247236 147614 247356 147642
rect 245752 143540 245804 143546
rect 245752 143482 245804 143488
rect 245936 143472 245988 143478
rect 245936 143414 245988 143420
rect 245948 138530 245976 143414
rect 245856 138502 245976 138530
rect 245856 133906 245884 138502
rect 247236 138038 247264 147614
rect 248340 143546 248368 153206
rect 248328 143540 248380 143546
rect 248328 143482 248380 143488
rect 247224 138032 247276 138038
rect 247224 137974 247276 137980
rect 247316 137964 247368 137970
rect 247316 137906 247368 137912
rect 245856 133890 245976 133906
rect 245856 133884 245988 133890
rect 245856 133878 245936 133884
rect 245936 133826 245988 133832
rect 245948 133795 245976 133826
rect 247328 128330 247356 137906
rect 248328 133952 248380 133958
rect 248328 133894 248380 133900
rect 247236 128302 247356 128330
rect 245752 124228 245804 124234
rect 245752 124170 245804 124176
rect 245764 114753 245792 124170
rect 247236 118726 247264 128302
rect 248340 124166 248368 133894
rect 248328 124160 248380 124166
rect 248328 124102 248380 124108
rect 247224 118720 247276 118726
rect 247224 118662 247276 118668
rect 247316 118652 247368 118658
rect 247316 118594 247368 118600
rect 245750 114744 245806 114753
rect 245750 114679 245806 114688
rect 245934 114608 245990 114617
rect 245934 114543 245990 114552
rect 245948 109750 245976 114543
rect 245936 109744 245988 109750
rect 245936 109686 245988 109692
rect 247328 109018 247356 118594
rect 248328 114572 248380 114578
rect 248328 114514 248380 114520
rect 247236 108990 247356 109018
rect 245752 104916 245804 104922
rect 245752 104858 245804 104864
rect 245764 95441 245792 104858
rect 247236 99414 247264 108990
rect 248340 104854 248368 114514
rect 248328 104848 248380 104854
rect 248328 104790 248380 104796
rect 247224 99408 247276 99414
rect 247224 99350 247276 99356
rect 247316 99340 247368 99346
rect 247316 99282 247368 99288
rect 245750 95432 245806 95441
rect 245750 95367 245806 95376
rect 245934 95296 245990 95305
rect 245934 95231 245990 95240
rect 245948 90438 245976 95231
rect 245936 90432 245988 90438
rect 245936 90374 245988 90380
rect 247328 89706 247356 99282
rect 248328 95260 248380 95266
rect 248328 95202 248380 95208
rect 247144 89678 247356 89706
rect 247144 86970 247172 89678
rect 247132 86964 247184 86970
rect 247132 86906 247184 86912
rect 248340 85542 248368 95202
rect 248328 85536 248380 85542
rect 248328 85478 248380 85484
rect 246212 83224 246264 83230
rect 246212 83166 246264 83172
rect 246224 74526 246252 83166
rect 247040 77308 247092 77314
rect 247040 77250 247092 77256
rect 246212 74520 246264 74526
rect 246212 74462 246264 74468
rect 247052 70258 247080 77250
rect 248328 75948 248380 75954
rect 248328 75890 248380 75896
rect 247052 70230 247172 70258
rect 246028 64932 246080 64938
rect 246028 64874 246080 64880
rect 246040 56710 246068 64874
rect 246028 56704 246080 56710
rect 246028 56646 246080 56652
rect 247144 56642 247172 70230
rect 248340 67794 248368 75890
rect 248328 67788 248380 67794
rect 248328 67730 248380 67736
rect 248328 67652 248380 67658
rect 248328 67594 248380 67600
rect 248340 66230 248368 67594
rect 248328 66224 248380 66230
rect 248328 66166 248380 66172
rect 247132 56636 247184 56642
rect 247132 56578 247184 56584
rect 247316 56636 247368 56642
rect 247316 56578 247368 56584
rect 248328 56636 248380 56642
rect 248328 56578 248380 56584
rect 245844 56568 245896 56574
rect 245844 56510 245896 56516
rect 245856 46918 245884 56510
rect 247328 47002 247356 56578
rect 247144 46974 247356 47002
rect 247144 46918 247172 46974
rect 248340 46918 248368 56578
rect 245844 46912 245896 46918
rect 245844 46854 245896 46860
rect 247132 46912 247184 46918
rect 247132 46854 247184 46860
rect 247408 46912 247460 46918
rect 247408 46854 247460 46860
rect 248328 46912 248380 46918
rect 248328 46854 248380 46860
rect 245752 46844 245804 46850
rect 245752 46786 245804 46792
rect 245764 45558 245792 46786
rect 247420 45558 247448 46854
rect 245752 45552 245804 45558
rect 245752 45494 245804 45500
rect 247408 45552 247460 45558
rect 247408 45494 247460 45500
rect 248328 37324 248380 37330
rect 248328 37266 248380 37272
rect 247408 37256 247460 37262
rect 247408 37198 247460 37204
rect 247420 31346 247448 37198
rect 247408 31340 247460 31346
rect 247408 31282 247460 31288
rect 245844 27668 245896 27674
rect 245844 27610 245896 27616
rect 247408 27668 247460 27674
rect 247408 27610 247460 27616
rect 245856 27266 245884 27610
rect 245844 27260 245896 27266
rect 245844 27202 245896 27208
rect 247420 22114 247448 27610
rect 247328 22086 247448 22114
rect 245936 19372 245988 19378
rect 245936 19314 245988 19320
rect 245660 5500 245712 5506
rect 245660 5442 245712 5448
rect 245948 4758 245976 19314
rect 245936 4752 245988 4758
rect 245936 4694 245988 4700
rect 247328 4554 247356 22086
rect 248340 19310 248368 37266
rect 248328 19304 248380 19310
rect 248328 19246 248380 19252
rect 247960 9716 248012 9722
rect 247960 9658 248012 9664
rect 247316 4548 247368 4554
rect 247316 4490 247368 4496
rect 246764 3664 246816 3670
rect 246764 3606 246816 3612
rect 246776 480 246804 3606
rect 247972 480 248000 9658
rect 248524 4622 248552 244038
rect 249168 242214 249196 244052
rect 249826 244038 250024 244066
rect 249708 242344 249760 242350
rect 249708 242286 249760 242292
rect 249156 242208 249208 242214
rect 249156 242150 249208 242156
rect 248512 4616 248564 4622
rect 248512 4558 248564 4564
rect 249720 3806 249748 242286
rect 249892 239352 249944 239358
rect 249892 239294 249944 239300
rect 249904 4486 249932 239294
rect 249996 4690 250024 244038
rect 250088 244038 250470 244066
rect 250088 239358 250116 244038
rect 251008 241602 251036 244052
rect 251284 244038 251666 244066
rect 250996 241596 251048 241602
rect 250996 241538 251048 241544
rect 251088 241596 251140 241602
rect 251088 241538 251140 241544
rect 250444 241528 250496 241534
rect 250444 241470 250496 241476
rect 250076 239352 250128 239358
rect 250076 239294 250128 239300
rect 249984 4684 250036 4690
rect 249984 4626 250036 4632
rect 249892 4480 249944 4486
rect 249892 4422 249944 4428
rect 249156 3800 249208 3806
rect 249156 3742 249208 3748
rect 249708 3800 249760 3806
rect 249708 3742 249760 3748
rect 250352 3800 250404 3806
rect 250352 3742 250404 3748
rect 249168 480 249196 3742
rect 250364 480 250392 3742
rect 250456 3738 250484 241470
rect 251100 3806 251128 241538
rect 251284 4418 251312 244038
rect 252296 242554 252324 244052
rect 252284 242548 252336 242554
rect 252284 242490 252336 242496
rect 252848 242282 252876 244052
rect 253124 244038 253506 244066
rect 252836 242276 252888 242282
rect 252836 242218 252888 242224
rect 252468 242208 252520 242214
rect 252468 242150 252520 242156
rect 252480 58070 252508 242150
rect 253124 239306 253152 244038
rect 254136 242894 254164 244052
rect 254124 242888 254176 242894
rect 254124 242830 254176 242836
rect 254584 242548 254636 242554
rect 254584 242490 254636 242496
rect 252848 239278 253152 239306
rect 252848 225010 252876 239278
rect 252652 225004 252704 225010
rect 252652 224946 252704 224952
rect 252836 225004 252888 225010
rect 252836 224946 252888 224952
rect 252664 224890 252692 224946
rect 252664 224862 252784 224890
rect 252756 215370 252784 224862
rect 252756 215342 252876 215370
rect 252848 205698 252876 215342
rect 252652 205692 252704 205698
rect 252652 205634 252704 205640
rect 252836 205692 252888 205698
rect 252836 205634 252888 205640
rect 252664 205578 252692 205634
rect 252664 205550 252784 205578
rect 252756 196058 252784 205550
rect 252756 196030 252876 196058
rect 252848 186386 252876 196030
rect 252652 186380 252704 186386
rect 252652 186322 252704 186328
rect 252836 186380 252888 186386
rect 252836 186322 252888 186328
rect 252664 186266 252692 186322
rect 252664 186238 252784 186266
rect 252756 183569 252784 186238
rect 252558 183560 252614 183569
rect 252558 183495 252614 183504
rect 252742 183560 252798 183569
rect 252742 183495 252798 183504
rect 252572 173942 252600 183495
rect 252560 173936 252612 173942
rect 252560 173878 252612 173884
rect 252836 173936 252888 173942
rect 252836 173878 252888 173884
rect 252848 167074 252876 173878
rect 252652 167068 252704 167074
rect 252652 167010 252704 167016
rect 252836 167068 252888 167074
rect 252836 167010 252888 167016
rect 252664 166954 252692 167010
rect 252664 166926 252784 166954
rect 252756 164218 252784 166926
rect 252744 164212 252796 164218
rect 252744 164154 252796 164160
rect 252744 157344 252796 157350
rect 252744 157286 252796 157292
rect 252756 154578 252784 157286
rect 252756 154550 252876 154578
rect 252848 147694 252876 154550
rect 252652 147688 252704 147694
rect 252836 147688 252888 147694
rect 252704 147636 252784 147642
rect 252652 147630 252784 147636
rect 252836 147630 252888 147636
rect 252664 147614 252784 147630
rect 252756 144906 252784 147614
rect 252744 144900 252796 144906
rect 252744 144842 252796 144848
rect 252744 137964 252796 137970
rect 252744 137906 252796 137912
rect 252756 135266 252784 137906
rect 252756 135238 252876 135266
rect 252848 128382 252876 135238
rect 252652 128376 252704 128382
rect 252836 128376 252888 128382
rect 252704 128324 252784 128330
rect 252652 128318 252784 128324
rect 252836 128318 252888 128324
rect 252664 128302 252784 128318
rect 252756 125594 252784 128302
rect 252744 125588 252796 125594
rect 252744 125530 252796 125536
rect 252744 118652 252796 118658
rect 252744 118594 252796 118600
rect 252756 115954 252784 118594
rect 252756 115926 252876 115954
rect 252848 109070 252876 115926
rect 252652 109064 252704 109070
rect 252836 109064 252888 109070
rect 252704 109012 252784 109018
rect 252652 109006 252784 109012
rect 252836 109006 252888 109012
rect 252664 108990 252784 109006
rect 252756 106282 252784 108990
rect 252744 106276 252796 106282
rect 252744 106218 252796 106224
rect 252744 99340 252796 99346
rect 252744 99282 252796 99288
rect 252756 96642 252784 99282
rect 252756 96614 252876 96642
rect 252848 89758 252876 96614
rect 252652 89752 252704 89758
rect 252836 89752 252888 89758
rect 252704 89700 252784 89706
rect 252652 89694 252784 89700
rect 252836 89694 252888 89700
rect 252664 89678 252784 89694
rect 252756 86970 252784 89678
rect 252744 86964 252796 86970
rect 252744 86906 252796 86912
rect 252836 77308 252888 77314
rect 252836 77250 252888 77256
rect 252848 67726 252876 77250
rect 252836 67720 252888 67726
rect 252836 67662 252888 67668
rect 252744 66292 252796 66298
rect 252744 66234 252796 66240
rect 252756 60874 252784 66234
rect 252756 60846 252876 60874
rect 252468 58064 252520 58070
rect 252468 58006 252520 58012
rect 252468 57928 252520 57934
rect 252468 57870 252520 57876
rect 252376 57044 252428 57050
rect 252376 56986 252428 56992
rect 252388 51066 252416 56986
rect 252376 51060 252428 51066
rect 252376 51002 252428 51008
rect 251272 4412 251324 4418
rect 251272 4354 251324 4360
rect 252480 3806 252508 57870
rect 252848 57050 252876 60846
rect 252836 57044 252888 57050
rect 252836 56986 252888 56992
rect 252744 51060 252796 51066
rect 252744 51002 252796 51008
rect 252756 43466 252784 51002
rect 252664 43438 252784 43466
rect 252664 38690 252692 43438
rect 252652 38684 252704 38690
rect 252652 38626 252704 38632
rect 252836 38684 252888 38690
rect 252836 38626 252888 38632
rect 252848 31906 252876 38626
rect 252848 31878 252968 31906
rect 252940 31634 252968 31878
rect 252756 31606 252968 31634
rect 252756 27606 252784 31606
rect 252744 27600 252796 27606
rect 252744 27542 252796 27548
rect 252836 18012 252888 18018
rect 252836 17954 252888 17960
rect 252848 4350 252876 17954
rect 252836 4344 252888 4350
rect 252836 4286 252888 4292
rect 251088 3800 251140 3806
rect 251088 3742 251140 3748
rect 251456 3800 251508 3806
rect 251456 3742 251508 3748
rect 252468 3800 252520 3806
rect 252468 3742 252520 3748
rect 250444 3732 250496 3738
rect 250444 3674 250496 3680
rect 251468 480 251496 3742
rect 252652 3732 252704 3738
rect 252652 3674 252704 3680
rect 252664 480 252692 3674
rect 253848 3324 253900 3330
rect 253848 3266 253900 3272
rect 253860 480 253888 3266
rect 254596 3262 254624 242490
rect 254688 242418 254716 244052
rect 255346 244038 255452 244066
rect 254676 242412 254728 242418
rect 254676 242354 254728 242360
rect 255228 242412 255280 242418
rect 255228 242354 255280 242360
rect 254676 242276 254728 242282
rect 254676 242218 254728 242224
rect 254688 3330 254716 242218
rect 254676 3324 254728 3330
rect 254676 3266 254728 3272
rect 254584 3256 254636 3262
rect 254584 3198 254636 3204
rect 255240 626 255268 242354
rect 255424 4282 255452 244038
rect 255884 241738 255912 244052
rect 256528 242622 256556 244052
rect 256804 244038 257186 244066
rect 256516 242616 256568 242622
rect 256516 242558 256568 242564
rect 256700 242548 256752 242554
rect 256700 242490 256752 242496
rect 256712 242434 256740 242490
rect 256620 242406 256740 242434
rect 255872 241732 255924 241738
rect 255872 241674 255924 241680
rect 255412 4276 255464 4282
rect 255412 4218 255464 4224
rect 255056 598 255268 626
rect 256620 610 256648 242406
rect 256804 3874 256832 244038
rect 257344 241732 257396 241738
rect 257344 241674 257396 241680
rect 256792 3868 256844 3874
rect 256792 3810 256844 3816
rect 257356 2854 257384 241674
rect 257724 241534 257752 244052
rect 257988 242888 258040 242894
rect 257988 242830 258040 242836
rect 257712 241528 257764 241534
rect 257712 241470 257764 241476
rect 258000 3330 258028 242830
rect 258368 242690 258396 244052
rect 258644 244038 259026 244066
rect 258356 242684 258408 242690
rect 258356 242626 258408 242632
rect 258644 241482 258672 244038
rect 259368 242684 259420 242690
rect 259368 242626 259420 242632
rect 258276 241454 258672 241482
rect 258276 219450 258304 241454
rect 258184 219422 258304 219450
rect 258184 215286 258212 219422
rect 258172 215280 258224 215286
rect 258172 215222 258224 215228
rect 258356 215280 258408 215286
rect 258356 215222 258408 215228
rect 258368 205578 258396 215222
rect 258276 205550 258396 205578
rect 258276 202881 258304 205550
rect 258078 202872 258134 202881
rect 258078 202807 258134 202816
rect 258262 202872 258318 202881
rect 258262 202807 258318 202816
rect 258092 193254 258120 202807
rect 258080 193248 258132 193254
rect 258080 193190 258132 193196
rect 258356 193248 258408 193254
rect 258356 193190 258408 193196
rect 258368 186266 258396 193190
rect 258276 186238 258396 186266
rect 258276 183569 258304 186238
rect 258078 183560 258134 183569
rect 258078 183495 258134 183504
rect 258262 183560 258318 183569
rect 258262 183495 258318 183504
rect 258092 173942 258120 183495
rect 258080 173936 258132 173942
rect 258080 173878 258132 173884
rect 258356 173936 258408 173942
rect 258356 173878 258408 173884
rect 258368 166954 258396 173878
rect 258276 166926 258396 166954
rect 258276 164218 258304 166926
rect 258080 164212 258132 164218
rect 258080 164154 258132 164160
rect 258264 164212 258316 164218
rect 258264 164154 258316 164160
rect 258092 154601 258120 164154
rect 258078 154592 258134 154601
rect 258078 154527 258134 154536
rect 258354 154592 258410 154601
rect 258354 154527 258410 154536
rect 258368 147642 258396 154527
rect 258276 147614 258396 147642
rect 258276 140026 258304 147614
rect 258092 139998 258304 140026
rect 258092 135289 258120 139998
rect 258078 135280 258134 135289
rect 258078 135215 258134 135224
rect 258354 135280 258410 135289
rect 258354 135215 258410 135224
rect 258368 128330 258396 135215
rect 258276 128302 258396 128330
rect 258276 120714 258304 128302
rect 258092 120686 258304 120714
rect 258092 115977 258120 120686
rect 258078 115968 258134 115977
rect 258078 115903 258134 115912
rect 258354 115968 258410 115977
rect 258354 115903 258410 115912
rect 258368 109018 258396 115903
rect 258276 108990 258396 109018
rect 258276 101402 258304 108990
rect 258092 101374 258304 101402
rect 258092 96665 258120 101374
rect 258078 96656 258134 96665
rect 258078 96591 258134 96600
rect 258354 96656 258410 96665
rect 258354 96591 258410 96600
rect 258368 89706 258396 96591
rect 258184 89678 258396 89706
rect 258184 86970 258212 89678
rect 258172 86964 258224 86970
rect 258172 86906 258224 86912
rect 258080 77308 258132 77314
rect 258080 77250 258132 77256
rect 258092 70258 258120 77250
rect 258092 70230 258212 70258
rect 258184 60722 258212 70230
rect 258172 60716 258224 60722
rect 258172 60658 258224 60664
rect 258356 60716 258408 60722
rect 258356 60658 258408 60664
rect 258368 57934 258396 60658
rect 258356 57928 258408 57934
rect 258356 57870 258408 57876
rect 258172 48340 258224 48346
rect 258172 48282 258224 48288
rect 258184 45234 258212 48282
rect 258184 45206 258304 45234
rect 258276 38826 258304 45206
rect 258264 38820 258316 38826
rect 258264 38762 258316 38768
rect 258264 38684 258316 38690
rect 258264 38626 258316 38632
rect 258276 38570 258304 38626
rect 258184 38542 258304 38570
rect 258184 31634 258212 38542
rect 258184 31606 258396 31634
rect 258368 22114 258396 31606
rect 258184 22086 258396 22114
rect 258184 7002 258212 22086
rect 258172 6996 258224 7002
rect 258172 6938 258224 6944
rect 258080 6928 258132 6934
rect 258080 6870 258132 6876
rect 258092 4214 258120 6870
rect 258080 4208 258132 4214
rect 258080 4150 258132 4156
rect 259380 3398 259408 242626
rect 259564 242185 259592 244052
rect 260208 242826 260236 244052
rect 260866 244038 261064 244066
rect 260196 242820 260248 242826
rect 260196 242762 260248 242768
rect 259550 242176 259606 242185
rect 259550 242111 259606 242120
rect 261036 3942 261064 244038
rect 261404 241738 261432 244052
rect 262048 242622 262076 244052
rect 262416 244038 262706 244066
rect 262036 242616 262088 242622
rect 262036 242558 262088 242564
rect 261576 241936 261628 241942
rect 261576 241878 261628 241884
rect 261392 241732 261444 241738
rect 261392 241674 261444 241680
rect 261484 241528 261536 241534
rect 261484 241470 261536 241476
rect 261496 4078 261524 241470
rect 261484 4072 261536 4078
rect 261484 4014 261536 4020
rect 261024 3936 261076 3942
rect 261024 3878 261076 3884
rect 261024 3800 261076 3806
rect 261024 3742 261076 3748
rect 258632 3392 258684 3398
rect 258632 3334 258684 3340
rect 259368 3392 259420 3398
rect 259368 3334 259420 3340
rect 257436 3324 257488 3330
rect 257436 3266 257488 3272
rect 257988 3324 258040 3330
rect 257988 3266 258040 3272
rect 257344 2848 257396 2854
rect 257344 2790 257396 2796
rect 256240 604 256292 610
rect 255056 480 255084 598
rect 256240 546 256292 552
rect 256608 604 256660 610
rect 256608 546 256660 552
rect 256252 480 256280 546
rect 257448 480 257476 3266
rect 258644 480 258672 3334
rect 259828 3324 259880 3330
rect 259828 3266 259880 3272
rect 259840 480 259868 3266
rect 261036 480 261064 3742
rect 261588 3398 261616 241878
rect 262416 4010 262444 244038
rect 262864 241732 262916 241738
rect 262864 241674 262916 241680
rect 262404 4004 262456 4010
rect 262404 3946 262456 3952
rect 261576 3392 261628 3398
rect 261576 3334 261628 3340
rect 262220 3392 262272 3398
rect 262220 3334 262272 3340
rect 262232 480 262260 3334
rect 262876 3194 262904 241674
rect 263244 241534 263272 244052
rect 263888 241942 263916 244052
rect 264164 244038 264454 244066
rect 263876 241936 263928 241942
rect 263876 241878 263928 241884
rect 263232 241528 263284 241534
rect 263232 241470 263284 241476
rect 263508 241528 263560 241534
rect 263508 241470 263560 241476
rect 263416 3936 263468 3942
rect 263416 3878 263468 3884
rect 262864 3188 262916 3194
rect 262864 3130 262916 3136
rect 263428 480 263456 3878
rect 263520 3398 263548 241470
rect 264164 239306 264192 244038
rect 265084 241738 265112 244052
rect 265728 242146 265756 244052
rect 266004 244038 266294 244066
rect 266464 244038 266938 244066
rect 265716 242140 265768 242146
rect 265716 242082 265768 242088
rect 265072 241732 265124 241738
rect 265072 241674 265124 241680
rect 263796 239278 264192 239306
rect 263796 215286 263824 239278
rect 266004 234870 266032 244038
rect 266268 242616 266320 242622
rect 266268 242558 266320 242564
rect 265164 234864 265216 234870
rect 265164 234806 265216 234812
rect 265992 234864 266044 234870
rect 265992 234806 266044 234812
rect 265176 231849 265204 234806
rect 265162 231840 265218 231849
rect 265162 231775 265218 231784
rect 265346 231840 265402 231849
rect 265346 231775 265402 231784
rect 265360 222222 265388 231775
rect 265164 222216 265216 222222
rect 265164 222158 265216 222164
rect 265348 222216 265400 222222
rect 265348 222158 265400 222164
rect 265176 215422 265204 222158
rect 265164 215416 265216 215422
rect 265164 215358 265216 215364
rect 263784 215280 263836 215286
rect 263784 215222 263836 215228
rect 263784 212560 263836 212566
rect 263784 212502 263836 212508
rect 265072 212560 265124 212566
rect 265072 212502 265124 212508
rect 263796 202881 263824 212502
rect 265084 205714 265112 212502
rect 264992 205686 265112 205714
rect 264992 205578 265020 205686
rect 264992 205550 265112 205578
rect 263598 202872 263654 202881
rect 263598 202807 263654 202816
rect 263782 202872 263838 202881
rect 263782 202807 263838 202816
rect 263612 193254 263640 202807
rect 263600 193248 263652 193254
rect 263600 193190 263652 193196
rect 263784 193248 263836 193254
rect 263784 193190 263836 193196
rect 263796 183569 263824 193190
rect 265084 186402 265112 205550
rect 264992 186374 265112 186402
rect 264992 186266 265020 186374
rect 264992 186238 265112 186266
rect 263598 183560 263654 183569
rect 263598 183495 263654 183504
rect 263782 183560 263838 183569
rect 263782 183495 263838 183504
rect 263612 173942 263640 183495
rect 263600 173936 263652 173942
rect 263600 173878 263652 173884
rect 263784 173936 263836 173942
rect 263784 173878 263836 173884
rect 263796 157434 263824 173878
rect 265084 167006 265112 186238
rect 265072 167000 265124 167006
rect 265072 166942 265124 166948
rect 265072 166864 265124 166870
rect 265072 166806 265124 166812
rect 265084 162858 265112 166806
rect 265072 162852 265124 162858
rect 265072 162794 265124 162800
rect 265256 162852 265308 162858
rect 265256 162794 265308 162800
rect 263704 157406 263824 157434
rect 263704 157298 263732 157406
rect 263704 157270 263824 157298
rect 263796 154562 263824 157270
rect 263784 154556 263836 154562
rect 263784 154498 263836 154504
rect 263784 148368 263836 148374
rect 263784 148310 263836 148316
rect 263796 143721 263824 148310
rect 265268 144945 265296 162794
rect 265070 144936 265126 144945
rect 265070 144871 265126 144880
rect 265254 144936 265310 144945
rect 265254 144871 265310 144880
rect 265084 144786 265112 144871
rect 265084 144758 265296 144786
rect 263782 143712 263838 143721
rect 263782 143647 263838 143656
rect 263782 143576 263838 143585
rect 263782 143511 263838 143520
rect 263796 142118 263824 143511
rect 263784 142112 263836 142118
rect 263784 142054 263836 142060
rect 265268 135289 265296 144758
rect 265070 135280 265126 135289
rect 265070 135215 265126 135224
rect 265254 135280 265310 135289
rect 265254 135215 265310 135224
rect 263784 132524 263836 132530
rect 263784 132466 263836 132472
rect 263796 124386 263824 132466
rect 265084 128874 265112 135215
rect 263704 124358 263824 124386
rect 264992 128846 265112 128874
rect 263704 124250 263732 124358
rect 263704 124222 263824 124250
rect 263796 122806 263824 124222
rect 264992 122806 265020 128846
rect 263784 122800 263836 122806
rect 263784 122742 263836 122748
rect 264980 122800 265032 122806
rect 264980 122742 265032 122748
rect 263784 114300 263836 114306
rect 263784 114242 263836 114248
rect 263796 104854 263824 114242
rect 265072 113212 265124 113218
rect 265072 113154 265124 113160
rect 265084 110922 265112 113154
rect 264992 110894 265112 110922
rect 263784 104848 263836 104854
rect 263784 104790 263836 104796
rect 263784 96892 263836 96898
rect 263784 96834 263836 96840
rect 263796 67833 263824 96834
rect 264992 89758 265020 110894
rect 264980 89752 265032 89758
rect 264980 89694 265032 89700
rect 265072 89684 265124 89690
rect 265072 89626 265124 89632
rect 265084 77314 265112 89626
rect 265072 77308 265124 77314
rect 265072 77250 265124 77256
rect 265072 77172 265124 77178
rect 265072 77114 265124 77120
rect 263782 67824 263838 67833
rect 265084 67794 265112 77114
rect 263782 67759 263838 67768
rect 265072 67788 265124 67794
rect 265072 67730 265124 67736
rect 263782 67688 263838 67697
rect 263782 67623 263838 67632
rect 265072 67652 265124 67658
rect 263796 66230 263824 67623
rect 265072 67594 265124 67600
rect 265084 66230 265112 67594
rect 263784 66224 263836 66230
rect 263784 66166 263836 66172
rect 265072 66224 265124 66230
rect 265072 66166 265124 66172
rect 265072 60716 265124 60722
rect 265072 60658 265124 60664
rect 265084 51082 265112 60658
rect 264992 51054 265112 51082
rect 263692 48340 263744 48346
rect 263692 48282 263744 48288
rect 263704 48249 263732 48282
rect 263690 48240 263746 48249
rect 263690 48175 263746 48184
rect 263782 48104 263838 48113
rect 263782 48039 263838 48048
rect 263796 22114 263824 48039
rect 264992 38690 265020 51054
rect 264980 38684 265032 38690
rect 264980 38626 265032 38632
rect 265072 38684 265124 38690
rect 265072 38626 265124 38632
rect 265084 29102 265112 38626
rect 264980 29096 265032 29102
rect 264980 29038 265032 29044
rect 265072 29096 265124 29102
rect 265072 29038 265124 29044
rect 264992 27606 265020 29038
rect 264980 27600 265032 27606
rect 264980 27542 265032 27548
rect 263704 22086 263824 22114
rect 263704 4146 263732 22086
rect 265072 18012 265124 18018
rect 265072 17954 265124 17960
rect 265084 12458 265112 17954
rect 264992 12430 265112 12458
rect 263692 4140 263744 4146
rect 263692 4082 263744 4088
rect 264612 4004 264664 4010
rect 264612 3946 264664 3952
rect 263508 3392 263560 3398
rect 263508 3334 263560 3340
rect 264624 480 264652 3946
rect 264992 2990 265020 12430
rect 266280 4146 266308 242558
rect 265808 4140 265860 4146
rect 265808 4082 265860 4088
rect 266268 4140 266320 4146
rect 266268 4082 266320 4088
rect 264980 2984 265032 2990
rect 264980 2926 265032 2932
rect 265820 480 265848 4082
rect 266464 3126 266492 244038
rect 267568 242826 267596 244052
rect 267844 244038 268134 244066
rect 267556 242820 267608 242826
rect 267556 242762 267608 242768
rect 267648 242140 267700 242146
rect 267648 242082 267700 242088
rect 267660 3126 267688 242082
rect 266452 3120 266504 3126
rect 266452 3062 266504 3068
rect 267004 3120 267056 3126
rect 267004 3062 267056 3068
rect 267648 3120 267700 3126
rect 267648 3062 267700 3068
rect 267016 480 267044 3062
rect 267844 3058 267872 244038
rect 268476 242072 268528 242078
rect 268476 242014 268528 242020
rect 268488 241754 268516 242014
rect 268764 242010 268792 244052
rect 269316 244038 269422 244066
rect 269592 244038 269974 244066
rect 268752 242004 268804 242010
rect 268752 241946 268804 241952
rect 269028 242004 269080 242010
rect 269028 241946 269080 241952
rect 268396 241726 268516 241754
rect 268396 4162 268424 241726
rect 268474 241632 268530 241641
rect 268474 241567 268530 241576
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 268304 4134 268424 4162
rect 267832 3052 267884 3058
rect 267832 2994 267884 3000
rect 268120 480 268148 4082
rect 268304 4078 268332 4134
rect 268292 4072 268344 4078
rect 268292 4014 268344 4020
rect 268488 3466 268516 241567
rect 269040 4146 269068 241946
rect 269212 238740 269264 238746
rect 269212 238682 269264 238688
rect 269224 4826 269252 238682
rect 269212 4820 269264 4826
rect 269212 4762 269264 4768
rect 269316 4298 269344 244038
rect 269592 238746 269620 244038
rect 270408 241732 270460 241738
rect 270408 241674 270460 241680
rect 269580 238740 269632 238746
rect 269580 238682 269632 238688
rect 269224 4270 269344 4298
rect 269028 4140 269080 4146
rect 269028 4082 269080 4088
rect 268476 3460 268528 3466
rect 268476 3402 268528 3408
rect 269224 2922 269252 4270
rect 270420 4146 270448 241674
rect 270604 241641 270632 244052
rect 271248 241670 271276 244052
rect 271524 244038 271814 244066
rect 271236 241664 271288 241670
rect 270590 241632 270646 241641
rect 271236 241606 271288 241612
rect 270590 241567 270646 241576
rect 271524 239358 271552 244038
rect 271788 241936 271840 241942
rect 271788 241878 271840 241884
rect 270500 239352 270552 239358
rect 270500 239294 270552 239300
rect 271512 239352 271564 239358
rect 271512 239294 271564 239300
rect 270512 234598 270540 239294
rect 270500 234592 270552 234598
rect 270500 234534 270552 234540
rect 270684 234592 270736 234598
rect 270684 234534 270736 234540
rect 270696 231849 270724 234534
rect 270498 231840 270554 231849
rect 270498 231775 270554 231784
rect 270682 231840 270738 231849
rect 270682 231775 270738 231784
rect 270512 224346 270540 231775
rect 270512 224318 270724 224346
rect 270696 215422 270724 224318
rect 270684 215416 270736 215422
rect 270684 215358 270736 215364
rect 270592 212560 270644 212566
rect 270592 212502 270644 212508
rect 270604 205714 270632 212502
rect 270512 205686 270632 205714
rect 270512 205578 270540 205686
rect 270512 205550 270632 205578
rect 270604 186402 270632 205550
rect 270512 186374 270632 186402
rect 270512 186266 270540 186374
rect 270512 186238 270632 186266
rect 270604 167006 270632 186238
rect 270592 167000 270644 167006
rect 270592 166942 270644 166948
rect 270592 166864 270644 166870
rect 270592 166806 270644 166812
rect 270604 162858 270632 166806
rect 270592 162852 270644 162858
rect 270592 162794 270644 162800
rect 270776 162852 270828 162858
rect 270776 162794 270828 162800
rect 270788 144945 270816 162794
rect 270498 144936 270554 144945
rect 270498 144871 270554 144880
rect 270774 144936 270830 144945
rect 270774 144871 270830 144880
rect 270512 135266 270540 144871
rect 270512 135238 270632 135266
rect 270604 128330 270632 135238
rect 270512 128302 270632 128330
rect 270512 115954 270540 128302
rect 270512 115926 270632 115954
rect 270604 109698 270632 115926
rect 270512 109670 270632 109698
rect 270512 103494 270540 109670
rect 270500 103488 270552 103494
rect 270500 103430 270552 103436
rect 270592 93900 270644 93906
rect 270592 93842 270644 93848
rect 270604 90386 270632 93842
rect 270512 90358 270632 90386
rect 270512 85542 270540 90358
rect 270500 85536 270552 85542
rect 270500 85478 270552 85484
rect 270592 75948 270644 75954
rect 270592 75890 270644 75896
rect 270604 70394 270632 75890
rect 270512 70366 270632 70394
rect 270512 70258 270540 70366
rect 270512 70230 270632 70258
rect 270604 51202 270632 70230
rect 270592 51196 270644 51202
rect 270592 51138 270644 51144
rect 270592 48340 270644 48346
rect 270592 48282 270644 48288
rect 270604 31890 270632 48282
rect 270592 31884 270644 31890
rect 270592 31826 270644 31832
rect 270592 27668 270644 27674
rect 270592 27610 270644 27616
rect 270604 19378 270632 27610
rect 270592 19372 270644 19378
rect 270592 19314 270644 19320
rect 270592 9716 270644 9722
rect 270592 9658 270644 9664
rect 270604 4894 270632 9658
rect 270592 4888 270644 4894
rect 270592 4830 270644 4836
rect 269304 4140 269356 4146
rect 269304 4082 269356 4088
rect 270408 4140 270460 4146
rect 270408 4082 270460 4088
rect 269212 2916 269264 2922
rect 269212 2858 269264 2864
rect 269316 480 269344 4082
rect 270500 3460 270552 3466
rect 270500 3402 270552 3408
rect 270512 480 270540 3402
rect 271800 626 271828 241878
rect 272444 241806 272472 244052
rect 272812 244038 273010 244066
rect 272432 241800 272484 241806
rect 272432 241742 272484 241748
rect 272812 239358 272840 244038
rect 273640 241874 273668 244052
rect 273916 244038 274298 244066
rect 273628 241868 273680 241874
rect 273628 241810 273680 241816
rect 273168 241800 273220 241806
rect 273168 241742 273220 241748
rect 272064 239352 272116 239358
rect 272064 239294 272116 239300
rect 272800 239352 272852 239358
rect 272800 239294 272852 239300
rect 272076 215286 272104 239294
rect 272064 215280 272116 215286
rect 272064 215222 272116 215228
rect 272064 212560 272116 212566
rect 272064 212502 272116 212508
rect 272076 202881 272104 212502
rect 271878 202872 271934 202881
rect 271878 202807 271934 202816
rect 272062 202872 272118 202881
rect 272062 202807 272118 202816
rect 271892 193254 271920 202807
rect 271880 193248 271932 193254
rect 271880 193190 271932 193196
rect 272064 193248 272116 193254
rect 272064 193190 272116 193196
rect 272076 183569 272104 193190
rect 271878 183560 271934 183569
rect 271878 183495 271934 183504
rect 272062 183560 272118 183569
rect 272062 183495 272118 183504
rect 271892 173942 271920 183495
rect 271880 173936 271932 173942
rect 271880 173878 271932 173884
rect 272064 173936 272116 173942
rect 272064 173878 272116 173884
rect 272076 157434 272104 173878
rect 271984 157406 272104 157434
rect 271984 157298 272012 157406
rect 271984 157270 272104 157298
rect 272076 154562 272104 157270
rect 271880 154556 271932 154562
rect 271880 154498 271932 154504
rect 272064 154556 272116 154562
rect 272064 154498 272116 154504
rect 271892 144945 271920 154498
rect 271878 144936 271934 144945
rect 271878 144871 271934 144880
rect 272062 144936 272118 144945
rect 272062 144871 272118 144880
rect 272076 135250 272104 144871
rect 271880 135244 271932 135250
rect 271880 135186 271932 135192
rect 272064 135244 272116 135250
rect 272064 135186 272116 135192
rect 271892 125633 271920 135186
rect 271878 125624 271934 125633
rect 271878 125559 271934 125568
rect 272062 125624 272118 125633
rect 272062 125559 272118 125568
rect 272076 116090 272104 125559
rect 271984 116062 272104 116090
rect 271984 115954 272012 116062
rect 271984 115926 272104 115954
rect 272076 114510 272104 115926
rect 271972 114504 272024 114510
rect 271972 114446 272024 114452
rect 272064 114504 272116 114510
rect 272064 114446 272116 114452
rect 271984 104938 272012 114446
rect 271984 104910 272104 104938
rect 272076 103494 272104 104910
rect 272064 103488 272116 103494
rect 272064 103430 272116 103436
rect 272064 93900 272116 93906
rect 272064 93842 272116 93848
rect 272076 85542 272104 93842
rect 272064 85536 272116 85542
rect 272064 85478 272116 85484
rect 272064 75948 272116 75954
rect 272064 75890 272116 75896
rect 272076 51134 272104 75890
rect 272064 51128 272116 51134
rect 272064 51070 272116 51076
rect 271880 48340 271932 48346
rect 271880 48282 271932 48288
rect 271892 41290 271920 48282
rect 271892 41262 272104 41290
rect 272076 28966 272104 41262
rect 271972 28960 272024 28966
rect 271972 28902 272024 28908
rect 272064 28960 272116 28966
rect 272064 28902 272116 28908
rect 271984 3534 272012 28902
rect 271972 3528 272024 3534
rect 271972 3470 272024 3476
rect 273180 626 273208 241742
rect 273916 239340 273944 244038
rect 274548 241664 274600 241670
rect 274548 241606 274600 241612
rect 273272 239312 273944 239340
rect 273272 234546 273300 239312
rect 273272 234518 273392 234546
rect 273364 205714 273392 234518
rect 273272 205686 273392 205714
rect 273272 205578 273300 205686
rect 273272 205550 273392 205578
rect 273364 186402 273392 205550
rect 273272 186374 273392 186402
rect 273272 186266 273300 186374
rect 273272 186238 273392 186266
rect 273364 167090 273392 186238
rect 273272 167062 273392 167090
rect 273272 166954 273300 167062
rect 273272 166926 273392 166954
rect 273364 147778 273392 166926
rect 273272 147750 273392 147778
rect 273272 147642 273300 147750
rect 273272 147614 273392 147642
rect 273364 128466 273392 147614
rect 273272 128438 273392 128466
rect 273272 128330 273300 128438
rect 273272 128302 273392 128330
rect 273364 109154 273392 128302
rect 273272 109126 273392 109154
rect 273272 109018 273300 109126
rect 273272 108990 273392 109018
rect 273364 89842 273392 108990
rect 273272 89814 273392 89842
rect 273272 89706 273300 89814
rect 273272 89678 273392 89706
rect 273364 70394 273392 89678
rect 273272 70366 273392 70394
rect 273272 70258 273300 70366
rect 273272 70230 273392 70258
rect 273364 51082 273392 70230
rect 273272 51054 273392 51082
rect 273272 50946 273300 51054
rect 273272 50918 273392 50946
rect 273364 31890 273392 50918
rect 273352 31884 273404 31890
rect 273352 31826 273404 31832
rect 273352 27668 273404 27674
rect 273352 27610 273404 27616
rect 273364 19258 273392 27610
rect 273272 19230 273392 19258
rect 273272 3670 273300 19230
rect 274560 4146 274588 241606
rect 274836 241534 274864 244052
rect 275480 242078 275508 244052
rect 275468 242072 275520 242078
rect 275468 242014 275520 242020
rect 275928 242072 275980 242078
rect 275928 242014 275980 242020
rect 274824 241528 274876 241534
rect 274824 241470 274876 241476
rect 274088 4140 274140 4146
rect 274088 4082 274140 4088
rect 274548 4140 274600 4146
rect 274548 4082 274600 4088
rect 273260 3664 273312 3670
rect 273260 3606 273312 3612
rect 271708 598 271828 626
rect 272904 598 273208 626
rect 271708 480 271736 598
rect 272904 480 272932 598
rect 274100 480 274128 4082
rect 275940 3058 275968 242014
rect 276124 241602 276152 244052
rect 276492 244038 276690 244066
rect 276112 241596 276164 241602
rect 276112 241538 276164 241544
rect 276492 239358 276520 244038
rect 277320 242486 277348 244052
rect 277308 242480 277360 242486
rect 277308 242422 277360 242428
rect 277400 242480 277452 242486
rect 277400 242422 277452 242428
rect 277412 242298 277440 242422
rect 277964 242350 277992 244052
rect 277320 242270 277440 242298
rect 277952 242344 278004 242350
rect 277952 242286 278004 242292
rect 276020 239352 276072 239358
rect 276020 239294 276072 239300
rect 276480 239352 276532 239358
rect 276480 239294 276532 239300
rect 276032 234546 276060 239294
rect 276032 234518 276152 234546
rect 276124 205714 276152 234518
rect 276032 205686 276152 205714
rect 276032 205578 276060 205686
rect 276032 205550 276152 205578
rect 276124 186402 276152 205550
rect 276032 186374 276152 186402
rect 276032 186266 276060 186374
rect 276032 186238 276152 186266
rect 276124 167090 276152 186238
rect 276032 167062 276152 167090
rect 276032 166954 276060 167062
rect 276032 166926 276152 166954
rect 276124 147778 276152 166926
rect 276032 147750 276152 147778
rect 276032 147642 276060 147750
rect 276032 147614 276152 147642
rect 276124 128466 276152 147614
rect 276032 128438 276152 128466
rect 276032 128330 276060 128438
rect 276032 128302 276152 128330
rect 276124 109154 276152 128302
rect 276032 109126 276152 109154
rect 276032 109018 276060 109126
rect 276032 108990 276152 109018
rect 276124 89842 276152 108990
rect 276032 89814 276152 89842
rect 276032 89706 276060 89814
rect 276032 89678 276152 89706
rect 276124 70394 276152 89678
rect 276032 70366 276152 70394
rect 276032 70258 276060 70366
rect 276032 70230 276152 70258
rect 276124 51082 276152 70230
rect 276032 51054 276152 51082
rect 276032 50946 276060 51054
rect 276032 50918 276152 50946
rect 276124 31770 276152 50918
rect 276032 31742 276152 31770
rect 276032 31634 276060 31742
rect 276032 31606 276152 31634
rect 276124 14498 276152 31606
rect 276032 14470 276152 14498
rect 276032 4078 276060 14470
rect 276020 4072 276072 4078
rect 276020 4014 276072 4020
rect 277320 3466 277348 242270
rect 278516 241874 278544 244052
rect 279160 242214 279188 244052
rect 279436 244038 279818 244066
rect 279148 242208 279200 242214
rect 279148 242150 279200 242156
rect 278504 241868 278556 241874
rect 278504 241810 278556 241816
rect 279436 239340 279464 244038
rect 280356 242758 280384 244052
rect 280344 242752 280396 242758
rect 280344 242694 280396 242700
rect 281000 242418 281028 244052
rect 281552 242554 281580 244052
rect 282196 242826 282224 244052
rect 282184 242820 282236 242826
rect 282184 242762 282236 242768
rect 282840 242690 282868 244052
rect 282828 242684 282880 242690
rect 282828 242626 282880 242632
rect 281540 242548 281592 242554
rect 281540 242490 281592 242496
rect 280988 242412 281040 242418
rect 280988 242354 281040 242360
rect 281448 242276 281500 242282
rect 281448 242218 281500 242224
rect 280068 242208 280120 242214
rect 280068 242150 280120 242156
rect 278792 239312 279464 239340
rect 278792 234546 278820 239312
rect 278792 234518 279004 234546
rect 278976 225078 279004 234518
rect 278964 225072 279016 225078
rect 278964 225014 279016 225020
rect 278872 222216 278924 222222
rect 278872 222158 278924 222164
rect 278884 215354 278912 222158
rect 278872 215348 278924 215354
rect 278872 215290 278924 215296
rect 278872 215212 278924 215218
rect 278872 215154 278924 215160
rect 278884 205714 278912 215154
rect 278792 205686 278912 205714
rect 278792 205578 278820 205686
rect 278792 205550 278912 205578
rect 278884 186402 278912 205550
rect 278792 186374 278912 186402
rect 278792 186266 278820 186374
rect 278792 186238 278912 186266
rect 278884 167090 278912 186238
rect 278792 167062 278912 167090
rect 278792 166954 278820 167062
rect 278792 166926 278912 166954
rect 278884 147778 278912 166926
rect 278792 147750 278912 147778
rect 278792 147642 278820 147750
rect 278792 147614 278912 147642
rect 278884 128466 278912 147614
rect 278792 128438 278912 128466
rect 278792 128330 278820 128438
rect 278792 128302 278912 128330
rect 278884 109154 278912 128302
rect 278792 109126 278912 109154
rect 278792 109018 278820 109126
rect 278792 108990 278912 109018
rect 278884 89842 278912 108990
rect 278792 89814 278912 89842
rect 278792 89706 278820 89814
rect 278792 89678 278912 89706
rect 278884 70394 278912 89678
rect 278792 70366 278912 70394
rect 278792 70258 278820 70366
rect 278792 70230 278912 70258
rect 278884 60722 278912 70230
rect 278872 60716 278924 60722
rect 278872 60658 278924 60664
rect 278964 60648 279016 60654
rect 278964 60590 279016 60596
rect 278976 41562 279004 60590
rect 278884 41534 279004 41562
rect 278884 41426 278912 41534
rect 278792 41398 278912 41426
rect 278792 41290 278820 41398
rect 278792 41262 278912 41290
rect 278884 22114 278912 41262
rect 278792 22086 278912 22114
rect 278792 21978 278820 22086
rect 278792 21950 278912 21978
rect 278884 3738 278912 21950
rect 278872 3732 278924 3738
rect 278872 3674 278924 3680
rect 277676 3596 277728 3602
rect 277676 3538 277728 3544
rect 276480 3460 276532 3466
rect 276480 3402 276532 3408
rect 277308 3460 277360 3466
rect 277308 3402 277360 3408
rect 275284 3052 275336 3058
rect 275284 2994 275336 3000
rect 275928 3052 275980 3058
rect 275928 2994 275980 3000
rect 275296 480 275324 2994
rect 276492 480 276520 3402
rect 277688 480 277716 3538
rect 278872 3460 278924 3466
rect 278872 3402 278924 3408
rect 278884 480 278912 3402
rect 280080 480 280108 242150
rect 280804 241528 280856 241534
rect 280804 241470 280856 241476
rect 280816 3330 280844 241470
rect 280804 3324 280856 3330
rect 280804 3266 280856 3272
rect 281460 610 281488 242218
rect 283392 241534 283420 244052
rect 283380 241528 283432 241534
rect 283380 241470 283432 241476
rect 283576 241346 283604 244174
rect 284680 242622 284708 244052
rect 284956 244038 285246 244066
rect 285784 244038 285890 244066
rect 284956 242978 284984 244038
rect 284772 242950 284984 242978
rect 284668 242616 284720 242622
rect 284668 242558 284720 242564
rect 284208 242344 284260 242350
rect 284208 242286 284260 242292
rect 283024 241318 283604 241346
rect 283024 3874 283052 241318
rect 283012 3868 283064 3874
rect 283012 3810 283064 3816
rect 282460 3664 282512 3670
rect 282460 3606 282512 3612
rect 281264 604 281316 610
rect 281264 546 281316 552
rect 281448 604 281500 610
rect 281448 546 281500 552
rect 281276 480 281304 546
rect 282472 480 282500 3606
rect 284220 2990 284248 242286
rect 284772 241346 284800 242950
rect 284944 242820 284996 242826
rect 284944 242762 284996 242768
rect 284312 241318 284800 241346
rect 284312 234546 284340 241318
rect 284312 234518 284432 234546
rect 284404 225026 284432 234518
rect 284404 224998 284524 225026
rect 284496 205698 284524 224998
rect 284300 205692 284352 205698
rect 284300 205634 284352 205640
rect 284484 205692 284536 205698
rect 284484 205634 284536 205640
rect 284312 205578 284340 205634
rect 284312 205550 284432 205578
rect 284404 196058 284432 205550
rect 284404 196030 284524 196058
rect 284496 186386 284524 196030
rect 284300 186380 284352 186386
rect 284300 186322 284352 186328
rect 284484 186380 284536 186386
rect 284484 186322 284536 186328
rect 284312 186266 284340 186322
rect 284312 186238 284432 186266
rect 284404 183569 284432 186238
rect 284390 183560 284446 183569
rect 284390 183495 284446 183504
rect 284666 183560 284722 183569
rect 284666 183495 284722 183504
rect 284680 173942 284708 183495
rect 284484 173936 284536 173942
rect 284484 173878 284536 173884
rect 284668 173936 284720 173942
rect 284668 173878 284720 173884
rect 284496 167074 284524 173878
rect 284300 167068 284352 167074
rect 284300 167010 284352 167016
rect 284484 167068 284536 167074
rect 284484 167010 284536 167016
rect 284312 166954 284340 167010
rect 284312 166926 284432 166954
rect 284404 164218 284432 166926
rect 284392 164212 284444 164218
rect 284392 164154 284444 164160
rect 284392 157344 284444 157350
rect 284392 157286 284444 157292
rect 284404 154578 284432 157286
rect 284404 154550 284524 154578
rect 284496 147694 284524 154550
rect 284300 147688 284352 147694
rect 284484 147688 284536 147694
rect 284352 147636 284432 147642
rect 284300 147630 284432 147636
rect 284484 147630 284536 147636
rect 284312 147614 284432 147630
rect 284404 144906 284432 147614
rect 284392 144900 284444 144906
rect 284392 144842 284444 144848
rect 284392 137964 284444 137970
rect 284392 137906 284444 137912
rect 284404 135266 284432 137906
rect 284404 135238 284524 135266
rect 284496 128382 284524 135238
rect 284300 128376 284352 128382
rect 284484 128376 284536 128382
rect 284352 128324 284432 128330
rect 284300 128318 284432 128324
rect 284484 128318 284536 128324
rect 284312 128302 284432 128318
rect 284404 125594 284432 128302
rect 284392 125588 284444 125594
rect 284392 125530 284444 125536
rect 284392 118652 284444 118658
rect 284392 118594 284444 118600
rect 284404 115954 284432 118594
rect 284404 115926 284524 115954
rect 284496 109070 284524 115926
rect 284300 109064 284352 109070
rect 284484 109064 284536 109070
rect 284352 109012 284432 109018
rect 284300 109006 284432 109012
rect 284484 109006 284536 109012
rect 284312 108990 284432 109006
rect 284404 106282 284432 108990
rect 284392 106276 284444 106282
rect 284392 106218 284444 106224
rect 284392 99340 284444 99346
rect 284392 99282 284444 99288
rect 284404 96642 284432 99282
rect 284404 96614 284524 96642
rect 284496 89758 284524 96614
rect 284300 89752 284352 89758
rect 284484 89752 284536 89758
rect 284352 89700 284432 89706
rect 284300 89694 284432 89700
rect 284484 89694 284536 89700
rect 284312 89678 284432 89694
rect 284404 86970 284432 89678
rect 284392 86964 284444 86970
rect 284392 86906 284444 86912
rect 284484 77308 284536 77314
rect 284484 77250 284536 77256
rect 284496 66298 284524 77250
rect 284392 66292 284444 66298
rect 284392 66234 284444 66240
rect 284484 66292 284536 66298
rect 284484 66234 284536 66240
rect 284404 60858 284432 66234
rect 284392 60852 284444 60858
rect 284392 60794 284444 60800
rect 284392 60716 284444 60722
rect 284392 60658 284444 60664
rect 284404 51134 284432 60658
rect 284392 51128 284444 51134
rect 284392 51070 284444 51076
rect 284300 51060 284352 51066
rect 284300 51002 284352 51008
rect 284312 48278 284340 51002
rect 284300 48272 284352 48278
rect 284300 48214 284352 48220
rect 284484 41404 284536 41410
rect 284484 41346 284536 41352
rect 284496 38622 284524 41346
rect 284484 38616 284536 38622
rect 284484 38558 284536 38564
rect 284392 29028 284444 29034
rect 284392 28970 284444 28976
rect 284404 24154 284432 28970
rect 284404 24126 284524 24154
rect 284496 3942 284524 24126
rect 284484 3936 284536 3942
rect 284484 3878 284536 3884
rect 284956 3398 284984 242762
rect 285784 4010 285812 244038
rect 286520 242894 286548 244052
rect 286508 242888 286560 242894
rect 286508 242830 286560 242836
rect 286324 242684 286376 242690
rect 286324 242626 286376 242632
rect 285772 4004 285824 4010
rect 285772 3946 285824 3952
rect 285956 3732 286008 3738
rect 285956 3674 286008 3680
rect 284944 3392 284996 3398
rect 284944 3334 284996 3340
rect 284760 3324 284812 3330
rect 284760 3266 284812 3272
rect 283656 2984 283708 2990
rect 283656 2926 283708 2932
rect 284208 2984 284260 2990
rect 284208 2926 284260 2932
rect 283668 480 283696 2926
rect 284772 480 284800 3266
rect 285968 480 285996 3674
rect 286336 3602 286364 242626
rect 287072 242146 287100 244052
rect 287060 242140 287112 242146
rect 287060 242082 287112 242088
rect 287716 242010 287744 244052
rect 287992 244038 288282 244066
rect 287704 242004 287756 242010
rect 287704 241946 287756 241952
rect 287992 241738 288020 244038
rect 288912 242826 288940 244052
rect 288900 242820 288952 242826
rect 288900 242762 288952 242768
rect 288256 242548 288308 242554
rect 288256 242490 288308 242496
rect 287980 241732 288032 241738
rect 287980 241674 288032 241680
rect 286324 3596 286376 3602
rect 286324 3538 286376 3544
rect 288268 3058 288296 242490
rect 288348 242412 288400 242418
rect 288348 242354 288400 242360
rect 287152 3052 287204 3058
rect 287152 2994 287204 3000
rect 288256 3052 288308 3058
rect 288256 2994 288308 3000
rect 287164 480 287192 2994
rect 288360 480 288388 242354
rect 289556 241942 289584 244052
rect 289544 241936 289596 241942
rect 289544 241878 289596 241884
rect 290108 241806 290136 244052
rect 290096 241800 290148 241806
rect 290096 241742 290148 241748
rect 290752 241670 290780 244052
rect 291396 242078 291424 244052
rect 291948 242486 291976 244052
rect 292592 242690 292620 244052
rect 292580 242684 292632 242690
rect 292580 242626 292632 242632
rect 291936 242480 291988 242486
rect 291936 242422 291988 242428
rect 292488 242480 292540 242486
rect 292488 242422 292540 242428
rect 291384 242072 291436 242078
rect 291384 242014 291436 242020
rect 291108 241800 291160 241806
rect 291108 241742 291160 241748
rect 290740 241664 290792 241670
rect 290740 241606 290792 241612
rect 290464 241596 290516 241602
rect 290464 241538 290516 241544
rect 289544 3460 289596 3466
rect 289544 3402 289596 3408
rect 289556 480 289584 3402
rect 290476 3330 290504 241538
rect 290464 3324 290516 3330
rect 290464 3266 290516 3272
rect 291120 2854 291148 241742
rect 291844 241528 291896 241534
rect 291844 241470 291896 241476
rect 291856 3398 291884 241470
rect 292500 4146 292528 242422
rect 293236 241534 293264 244052
rect 293788 242214 293816 244052
rect 294432 242282 294460 244052
rect 294616 244038 295090 244066
rect 294420 242276 294472 242282
rect 294420 242218 294472 242224
rect 293776 242208 293828 242214
rect 293776 242150 293828 242156
rect 293224 241528 293276 241534
rect 293224 241470 293276 241476
rect 294616 241346 294644 244038
rect 294788 242752 294840 242758
rect 294788 242694 294840 242700
rect 294156 241318 294644 241346
rect 291936 4140 291988 4146
rect 291936 4082 291988 4088
rect 292488 4140 292540 4146
rect 292488 4082 292540 4088
rect 291844 3392 291896 3398
rect 291844 3334 291896 3340
rect 291108 2848 291160 2854
rect 291108 2790 291160 2796
rect 290740 604 290792 610
rect 290740 546 290792 552
rect 290752 480 290780 546
rect 291948 480 291976 4082
rect 294156 3670 294184 241318
rect 294800 238762 294828 242694
rect 295628 242350 295656 244052
rect 295616 242344 295668 242350
rect 295616 242286 295668 242292
rect 296272 241602 296300 244052
rect 296824 242758 296852 244052
rect 296812 242752 296864 242758
rect 296812 242694 296864 242700
rect 297468 242554 297496 244052
rect 297456 242548 297508 242554
rect 297456 242490 297508 242496
rect 298112 242418 298140 244052
rect 298100 242412 298152 242418
rect 298100 242354 298152 242360
rect 296260 241596 296312 241602
rect 296260 241538 296312 241544
rect 297456 241596 297508 241602
rect 297456 241538 297508 241544
rect 297364 241528 297416 241534
rect 297364 241470 297416 241476
rect 294616 238734 294828 238762
rect 294616 3738 294644 238734
rect 295524 4140 295576 4146
rect 295524 4082 295576 4088
rect 294604 3732 294656 3738
rect 294604 3674 294656 3680
rect 294144 3664 294196 3670
rect 294144 3606 294196 3612
rect 294328 3392 294380 3398
rect 294328 3334 294380 3340
rect 293132 3052 293184 3058
rect 293132 2994 293184 3000
rect 293144 480 293172 2994
rect 294340 480 294368 3334
rect 295536 480 295564 4082
rect 297376 3466 297404 241470
rect 297364 3460 297416 3466
rect 297364 3402 297416 3408
rect 297468 3398 297496 241538
rect 298664 241534 298692 244052
rect 299308 241806 299336 244052
rect 299952 242486 299980 244052
rect 299940 242480 299992 242486
rect 299940 242422 299992 242428
rect 299296 241800 299348 241806
rect 299296 241742 299348 241748
rect 298744 241664 298796 241670
rect 298744 241606 298796 241612
rect 298652 241528 298704 241534
rect 298652 241470 298704 241476
rect 298756 4146 298784 241606
rect 300504 241534 300532 244052
rect 301148 241602 301176 244052
rect 301792 241670 301820 244052
rect 302358 244038 302464 244066
rect 301780 241664 301832 241670
rect 301780 241606 301832 241612
rect 301136 241596 301188 241602
rect 301136 241538 301188 241544
rect 301504 241596 301556 241602
rect 301504 241538 301556 241544
rect 298836 241528 298888 241534
rect 298836 241470 298888 241476
rect 300492 241528 300544 241534
rect 300492 241470 300544 241476
rect 298744 4140 298796 4146
rect 298744 4082 298796 4088
rect 297916 3460 297968 3466
rect 297916 3402 297968 3408
rect 297456 3392 297508 3398
rect 297456 3334 297508 3340
rect 296720 2916 296772 2922
rect 296720 2858 296772 2864
rect 296732 480 296760 2858
rect 297928 480 297956 3402
rect 298848 3058 298876 241470
rect 300308 3664 300360 3670
rect 300308 3606 300360 3612
rect 299112 3188 299164 3194
rect 299112 3130 299164 3136
rect 298836 3052 298888 3058
rect 298836 2994 298888 3000
rect 299124 480 299152 3130
rect 300320 480 300348 3606
rect 301412 3528 301464 3534
rect 301412 3470 301464 3476
rect 301424 480 301452 3470
rect 301516 3194 301544 241538
rect 301596 241528 301648 241534
rect 301596 241470 301648 241476
rect 301608 3466 301636 241470
rect 302146 40216 302202 40225
rect 302330 40216 302386 40225
rect 302202 40174 302330 40202
rect 302146 40151 302202 40160
rect 302330 40151 302386 40160
rect 302146 16824 302202 16833
rect 302330 16824 302386 16833
rect 302202 16782 302330 16810
rect 302146 16759 302202 16768
rect 302330 16759 302386 16768
rect 301596 3460 301648 3466
rect 301596 3402 301648 3408
rect 301504 3188 301556 3194
rect 301504 3130 301556 3136
rect 302436 2922 302464 244038
rect 302884 241664 302936 241670
rect 302884 241606 302936 241612
rect 302608 4072 302660 4078
rect 302608 4014 302660 4020
rect 302424 2916 302476 2922
rect 302424 2858 302476 2864
rect 302620 480 302648 4014
rect 302896 3534 302924 241606
rect 302988 241534 303016 244052
rect 303632 241602 303660 244052
rect 303620 241596 303672 241602
rect 303620 241538 303672 241544
rect 302976 241528 303028 241534
rect 302976 241470 303028 241476
rect 303816 241466 303844 244174
rect 304828 241670 304856 244052
rect 304816 241664 304868 241670
rect 304816 241606 304868 241612
rect 305380 241602 305408 244052
rect 304264 241596 304316 241602
rect 304264 241538 304316 241544
rect 305368 241596 305420 241602
rect 305368 241538 305420 241544
rect 303804 241460 303856 241466
rect 303804 241402 303856 241408
rect 303896 231872 303948 231878
rect 303896 231814 303948 231820
rect 303908 144906 303936 231814
rect 303896 144900 303948 144906
rect 303896 144842 303948 144848
rect 303988 144900 304040 144906
rect 303988 144842 304040 144848
rect 304000 137986 304028 144842
rect 303908 137958 304028 137986
rect 303908 125594 303936 137958
rect 303896 125588 303948 125594
rect 303896 125530 303948 125536
rect 303988 125588 304040 125594
rect 303988 125530 304040 125536
rect 304000 118674 304028 125530
rect 303908 118646 304028 118674
rect 303908 106298 303936 118646
rect 303908 106270 304028 106298
rect 304000 96665 304028 106270
rect 303618 96656 303674 96665
rect 303986 96656 304042 96665
rect 303618 96591 303620 96600
rect 303672 96591 303674 96600
rect 303712 96620 303764 96626
rect 303620 96562 303672 96568
rect 303986 96591 304042 96600
rect 303712 96562 303764 96568
rect 303724 86986 303752 96562
rect 303724 86958 303844 86986
rect 303816 77330 303844 86958
rect 303816 77302 303936 77330
rect 303908 77246 303936 77302
rect 303896 77240 303948 77246
rect 303896 77182 303948 77188
rect 303896 70236 303948 70242
rect 303896 70178 303948 70184
rect 303908 58002 303936 70178
rect 303620 57996 303672 58002
rect 303620 57938 303672 57944
rect 303896 57996 303948 58002
rect 303896 57938 303948 57944
rect 303632 3670 303660 57938
rect 303804 4140 303856 4146
rect 303804 4082 303856 4088
rect 303620 3664 303672 3670
rect 303620 3606 303672 3612
rect 302884 3528 302936 3534
rect 302884 3470 302936 3476
rect 303816 480 303844 4082
rect 304276 4078 304304 241538
rect 306024 241534 306052 244052
rect 306392 244038 306682 244066
rect 306392 241584 306420 244038
rect 306208 241556 306420 241584
rect 304908 241528 304960 241534
rect 304908 241470 304960 241476
rect 306012 241528 306064 241534
rect 306012 241470 306064 241476
rect 304920 4146 304948 241470
rect 306208 4146 306236 241556
rect 307220 241534 307248 244052
rect 307772 244038 307878 244066
rect 308048 244038 308522 244066
rect 307208 241528 307260 241534
rect 307208 241470 307260 241476
rect 306288 241460 306340 241466
rect 306288 241402 306340 241408
rect 304908 4140 304960 4146
rect 304908 4082 304960 4088
rect 305000 4140 305052 4146
rect 305000 4082 305052 4088
rect 306196 4140 306248 4146
rect 306196 4082 306248 4088
rect 304264 4072 304316 4078
rect 304264 4014 304316 4020
rect 305012 480 305040 4082
rect 306300 4026 306328 241402
rect 307668 67584 307720 67590
rect 307668 67526 307720 67532
rect 307680 58041 307708 67526
rect 307666 58032 307722 58041
rect 307666 57967 307722 57976
rect 307772 4026 307800 244038
rect 308048 225010 308076 244038
rect 309060 241584 309088 244052
rect 309060 241556 309364 241584
rect 307852 225004 307904 225010
rect 307852 224946 307904 224952
rect 308036 225004 308088 225010
rect 308036 224946 308088 224952
rect 307864 224890 307892 224946
rect 307864 224862 307984 224890
rect 307956 215370 307984 224862
rect 307956 215342 308076 215370
rect 308048 205698 308076 215342
rect 307852 205692 307904 205698
rect 307852 205634 307904 205640
rect 308036 205692 308088 205698
rect 308036 205634 308088 205640
rect 307864 205578 307892 205634
rect 307864 205550 307984 205578
rect 307956 196058 307984 205550
rect 307956 196030 308076 196058
rect 308048 186386 308076 196030
rect 307852 186380 307904 186386
rect 307852 186322 307904 186328
rect 308036 186380 308088 186386
rect 308036 186322 308088 186328
rect 307864 186266 307892 186322
rect 307864 186238 307984 186266
rect 307956 183569 307984 186238
rect 307942 183560 307998 183569
rect 307942 183495 307998 183504
rect 308218 183560 308274 183569
rect 308218 183495 308274 183504
rect 308232 173942 308260 183495
rect 308036 173936 308088 173942
rect 308036 173878 308088 173884
rect 308220 173936 308272 173942
rect 308220 173878 308272 173884
rect 308048 167074 308076 173878
rect 307852 167068 307904 167074
rect 307852 167010 307904 167016
rect 308036 167068 308088 167074
rect 308036 167010 308088 167016
rect 307864 166954 307892 167010
rect 307864 166926 307984 166954
rect 307956 164218 307984 166926
rect 307944 164212 307996 164218
rect 307944 164154 307996 164160
rect 307944 157344 307996 157350
rect 307944 157286 307996 157292
rect 307956 154578 307984 157286
rect 307956 154550 308076 154578
rect 308048 147694 308076 154550
rect 307852 147688 307904 147694
rect 308036 147688 308088 147694
rect 307904 147636 307984 147642
rect 307852 147630 307984 147636
rect 308036 147630 308088 147636
rect 307864 147614 307984 147630
rect 307956 144906 307984 147614
rect 307944 144900 307996 144906
rect 307944 144842 307996 144848
rect 307944 137964 307996 137970
rect 307944 137906 307996 137912
rect 307956 135266 307984 137906
rect 307956 135238 308076 135266
rect 308048 128382 308076 135238
rect 307852 128376 307904 128382
rect 308036 128376 308088 128382
rect 307904 128324 307984 128330
rect 307852 128318 307984 128324
rect 308036 128318 308088 128324
rect 307864 128302 307984 128318
rect 307956 125594 307984 128302
rect 307944 125588 307996 125594
rect 307944 125530 307996 125536
rect 307944 118652 307996 118658
rect 307944 118594 307996 118600
rect 307956 115954 307984 118594
rect 307956 115926 308076 115954
rect 308048 109070 308076 115926
rect 307852 109064 307904 109070
rect 308036 109064 308088 109070
rect 307904 109012 307984 109018
rect 307852 109006 307984 109012
rect 308036 109006 308088 109012
rect 307864 108990 307984 109006
rect 307956 106282 307984 108990
rect 307944 106276 307996 106282
rect 307944 106218 307996 106224
rect 307944 99340 307996 99346
rect 307944 99282 307996 99288
rect 307956 96642 307984 99282
rect 307956 96614 308076 96642
rect 308048 89758 308076 96614
rect 307852 89752 307904 89758
rect 308036 89752 308088 89758
rect 307904 89700 307984 89706
rect 307852 89694 307984 89700
rect 308036 89694 308088 89700
rect 307864 89678 307984 89694
rect 307956 86970 307984 89678
rect 307944 86964 307996 86970
rect 307944 86906 307996 86912
rect 308036 77308 308088 77314
rect 308036 77250 308088 77256
rect 308048 67726 308076 77250
rect 307944 67720 307996 67726
rect 307944 67662 307996 67668
rect 308036 67720 308088 67726
rect 308036 67662 308088 67668
rect 307956 67590 307984 67662
rect 307944 67584 307996 67590
rect 307944 67526 307996 67532
rect 307850 58032 307906 58041
rect 307850 57967 307906 57976
rect 307864 57934 307892 57967
rect 307852 57928 307904 57934
rect 307852 57870 307904 57876
rect 307944 48340 307996 48346
rect 307944 48282 307996 48288
rect 307956 48249 307984 48282
rect 307942 48240 307998 48249
rect 307942 48175 307998 48184
rect 308034 38720 308090 38729
rect 308034 38655 308090 38664
rect 308048 38622 308076 38655
rect 308036 38616 308088 38622
rect 308036 38558 308088 38564
rect 307944 29028 307996 29034
rect 307944 28970 307996 28976
rect 307956 28914 307984 28970
rect 307956 28886 308076 28914
rect 308048 21978 308076 28886
rect 307956 21950 308076 21978
rect 307956 12458 307984 21950
rect 309336 14498 309364 241556
rect 309704 241534 309732 244052
rect 310348 241602 310376 244052
rect 310336 241596 310388 241602
rect 310336 241538 310388 241544
rect 310900 241534 310928 244052
rect 311558 244038 311848 244066
rect 309692 241528 309744 241534
rect 309692 241470 309744 241476
rect 310428 241528 310480 241534
rect 310428 241470 310480 241476
rect 310888 241528 310940 241534
rect 310888 241470 310940 241476
rect 309336 14470 309456 14498
rect 307956 12430 308076 12458
rect 308048 4146 308076 12430
rect 309428 9722 309456 14470
rect 309416 9716 309468 9722
rect 309416 9658 309468 9664
rect 309784 9716 309836 9722
rect 309784 9658 309836 9664
rect 308036 4140 308088 4146
rect 308036 4082 308088 4088
rect 308588 4140 308640 4146
rect 308588 4082 308640 4088
rect 306208 3998 306328 4026
rect 307404 3998 307800 4026
rect 306208 480 306236 3998
rect 307404 480 307432 3998
rect 308600 480 308628 4082
rect 309796 480 309824 9658
rect 310440 4146 310468 241470
rect 310428 4140 310480 4146
rect 310428 4082 310480 4088
rect 310980 4140 311032 4146
rect 310980 4082 311032 4088
rect 310992 480 311020 4082
rect 311820 3466 311848 244038
rect 312188 241602 312216 244052
rect 312740 242894 312768 244052
rect 312728 242888 312780 242894
rect 312728 242830 312780 242836
rect 313384 242622 313412 244052
rect 313936 242690 313964 244052
rect 314580 242758 314608 244052
rect 314568 242752 314620 242758
rect 314568 242694 314620 242700
rect 313924 242684 313976 242690
rect 313924 242626 313976 242632
rect 313372 242616 313424 242622
rect 313372 242558 313424 242564
rect 315224 242350 315252 244052
rect 315790 244038 315988 244066
rect 315212 242344 315264 242350
rect 315212 242286 315264 242292
rect 311900 241596 311952 241602
rect 311900 241538 311952 241544
rect 312176 241596 312228 241602
rect 312176 241538 312228 241544
rect 314844 241596 314896 241602
rect 314844 241538 314896 241544
rect 311808 3460 311860 3466
rect 311808 3402 311860 3408
rect 311912 3346 311940 241538
rect 312544 241528 312596 241534
rect 312544 241470 312596 241476
rect 312556 3534 312584 241470
rect 312544 3528 312596 3534
rect 312544 3470 312596 3476
rect 313372 3528 313424 3534
rect 313372 3470 313424 3476
rect 314856 3482 314884 241538
rect 311912 3318 312216 3346
rect 312188 480 312216 3318
rect 313384 480 313412 3470
rect 314568 3460 314620 3466
rect 314856 3454 315804 3482
rect 315960 3466 315988 244038
rect 316040 242888 316092 242894
rect 316040 242830 316092 242836
rect 314568 3402 314620 3408
rect 314580 480 314608 3402
rect 315776 480 315804 3454
rect 315948 3460 316000 3466
rect 315948 3402 316000 3408
rect 316052 3346 316080 242830
rect 316420 241602 316448 244052
rect 316776 242752 316828 242758
rect 316776 242694 316828 242700
rect 316684 242616 316736 242622
rect 316684 242558 316736 242564
rect 316408 241596 316460 241602
rect 316408 241538 316460 241544
rect 316696 3602 316724 242558
rect 316788 3670 316816 242694
rect 317064 241670 317092 244052
rect 317616 242282 317644 244052
rect 317604 242276 317656 242282
rect 317604 242218 317656 242224
rect 318260 242214 318288 244052
rect 318248 242208 318300 242214
rect 318248 242150 318300 242156
rect 318904 241738 318932 244052
rect 319470 244038 320036 244066
rect 319076 242684 319128 242690
rect 319076 242626 319128 242632
rect 318892 241732 318944 241738
rect 318892 241674 318944 241680
rect 317052 241664 317104 241670
rect 317052 241606 317104 241612
rect 318798 16824 318854 16833
rect 318798 16759 318800 16768
rect 318852 16759 318854 16768
rect 318800 16730 318852 16736
rect 316776 3664 316828 3670
rect 316776 3606 316828 3612
rect 316684 3596 316736 3602
rect 316684 3538 316736 3544
rect 318064 3596 318116 3602
rect 318064 3538 318116 3544
rect 316052 3318 317000 3346
rect 316972 480 317000 3318
rect 318076 480 318104 3538
rect 319088 626 319116 242626
rect 320008 3874 320036 244038
rect 319996 3868 320048 3874
rect 319996 3810 320048 3816
rect 320100 3806 320128 244052
rect 320652 241534 320680 244052
rect 321310 244038 321416 244066
rect 320824 241596 320876 241602
rect 320824 241538 320876 241544
rect 320640 241528 320692 241534
rect 320640 241470 320692 241476
rect 320088 3800 320140 3806
rect 320088 3742 320140 3748
rect 320456 3664 320508 3670
rect 320456 3606 320508 3612
rect 319088 598 319208 626
rect 319180 592 319208 598
rect 319180 564 319300 592
rect 319272 480 319300 564
rect 320468 480 320496 3606
rect 320836 3262 320864 241538
rect 321282 40216 321338 40225
rect 321282 40151 321284 40160
rect 321336 40151 321338 40160
rect 321284 40122 321336 40128
rect 321388 3738 321416 244038
rect 321652 242344 321704 242350
rect 321652 242286 321704 242292
rect 321468 241528 321520 241534
rect 321468 241470 321520 241476
rect 321480 4078 321508 241470
rect 321558 40216 321614 40225
rect 321558 40151 321560 40160
rect 321612 40151 321614 40160
rect 321560 40122 321612 40128
rect 321558 16824 321614 16833
rect 321558 16759 321560 16768
rect 321612 16759 321614 16768
rect 321560 16730 321612 16736
rect 321468 4072 321520 4078
rect 321468 4014 321520 4020
rect 321376 3732 321428 3738
rect 321376 3674 321428 3680
rect 320824 3256 320876 3262
rect 320824 3198 320876 3204
rect 321664 480 321692 242286
rect 321940 241534 321968 244052
rect 322506 244038 322796 244066
rect 322204 241664 322256 241670
rect 322204 241606 322256 241612
rect 321928 241528 321980 241534
rect 321928 241470 321980 241476
rect 322216 3534 322244 241606
rect 322768 3670 322796 244038
rect 323136 241534 323164 244052
rect 323794 244038 324268 244066
rect 323584 241732 323636 241738
rect 323584 241674 323636 241680
rect 322848 241528 322900 241534
rect 322848 241470 322900 241476
rect 323124 241528 323176 241534
rect 323124 241470 323176 241476
rect 322756 3664 322808 3670
rect 322756 3606 322808 3612
rect 322860 3618 322888 241470
rect 322860 3590 322980 3618
rect 322204 3528 322256 3534
rect 322204 3470 322256 3476
rect 322848 3460 322900 3466
rect 322848 3402 322900 3408
rect 322860 480 322888 3402
rect 322952 3398 322980 3590
rect 322940 3392 322992 3398
rect 322940 3334 322992 3340
rect 323596 3330 323624 241674
rect 324136 241528 324188 241534
rect 324136 241470 324188 241476
rect 324148 4146 324176 241470
rect 324136 4140 324188 4146
rect 324136 4082 324188 4088
rect 324240 3602 324268 244038
rect 324332 241534 324360 244052
rect 324976 242350 325004 244052
rect 325620 242622 325648 244052
rect 325608 242616 325660 242622
rect 325608 242558 325660 242564
rect 324964 242344 325016 242350
rect 324964 242286 325016 242292
rect 325792 242276 325844 242282
rect 325792 242218 325844 242224
rect 324320 241528 324372 241534
rect 324320 241470 324372 241476
rect 325608 241528 325660 241534
rect 325608 241470 325660 241476
rect 324228 3596 324280 3602
rect 324228 3538 324280 3544
rect 325620 3534 325648 241470
rect 325240 3528 325292 3534
rect 325240 3470 325292 3476
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 323584 3324 323636 3330
rect 323584 3266 323636 3272
rect 324044 3256 324096 3262
rect 324044 3198 324096 3204
rect 324056 480 324084 3198
rect 325252 480 325280 3470
rect 325804 610 325832 242218
rect 326172 241534 326200 244052
rect 326816 242418 326844 244052
rect 326804 242412 326856 242418
rect 326804 242354 326856 242360
rect 327264 242208 327316 242214
rect 327264 242150 327316 242156
rect 326160 241528 326212 241534
rect 326160 241470 326212 241476
rect 326988 241528 327040 241534
rect 326988 241470 327040 241476
rect 327000 3466 327028 241470
rect 326988 3460 327040 3466
rect 326988 3402 327040 3408
rect 327276 626 327304 242150
rect 327460 241534 327488 244052
rect 328026 244038 328316 244066
rect 327448 241528 327500 241534
rect 327448 241470 327500 241476
rect 328288 3942 328316 244038
rect 328656 242690 328684 244052
rect 328644 242684 328696 242690
rect 328644 242626 328696 242632
rect 329208 241602 329236 244052
rect 329852 242758 329880 244052
rect 330510 244038 330800 244066
rect 331062 244038 331168 244066
rect 329840 242752 329892 242758
rect 329840 242694 329892 242700
rect 330484 242344 330536 242350
rect 330484 242286 330536 242292
rect 329196 241596 329248 241602
rect 329196 241538 329248 241544
rect 328368 241528 328420 241534
rect 328368 241470 328420 241476
rect 328380 4010 328408 241470
rect 328368 4004 328420 4010
rect 328368 3946 328420 3952
rect 328276 3936 328328 3942
rect 328276 3878 328328 3884
rect 330024 3868 330076 3874
rect 330024 3810 330076 3816
rect 328828 3324 328880 3330
rect 328828 3266 328880 3272
rect 325792 604 325844 610
rect 325792 546 325844 552
rect 326436 604 326488 610
rect 327276 598 327672 626
rect 326436 546 326488 552
rect 326448 480 326476 546
rect 327644 480 327672 598
rect 328840 480 328868 3266
rect 330036 480 330064 3810
rect 330496 3330 330524 242286
rect 330772 241738 330800 244038
rect 330760 241732 330812 241738
rect 330760 241674 330812 241680
rect 331140 3874 331168 244038
rect 331692 242826 331720 244052
rect 331680 242820 331732 242826
rect 331680 242762 331732 242768
rect 332336 242214 332364 244052
rect 332324 242208 332376 242214
rect 332324 242150 332376 242156
rect 332888 241534 332916 244052
rect 333532 242554 333560 244052
rect 333520 242548 333572 242554
rect 333520 242490 333572 242496
rect 334176 241806 334204 244052
rect 334742 244038 335308 244066
rect 334164 241800 334216 241806
rect 334164 241742 334216 241748
rect 333244 241596 333296 241602
rect 333244 241538 333296 241544
rect 332876 241528 332928 241534
rect 332876 241470 332928 241476
rect 333256 4078 333284 241538
rect 333888 241528 333940 241534
rect 333888 241470 333940 241476
rect 332416 4072 332468 4078
rect 332416 4014 332468 4020
rect 333244 4072 333296 4078
rect 333244 4014 333296 4020
rect 331128 3868 331180 3874
rect 331128 3810 331180 3816
rect 331220 3800 331272 3806
rect 331220 3742 331272 3748
rect 330484 3324 330536 3330
rect 330484 3266 330536 3272
rect 331232 480 331260 3742
rect 332428 480 332456 4014
rect 333900 3806 333928 241470
rect 333888 3800 333940 3806
rect 333888 3742 333940 3748
rect 335280 3738 335308 244038
rect 335372 241942 335400 244052
rect 336016 242350 336044 244052
rect 336004 242344 336056 242350
rect 336004 242286 336056 242292
rect 335360 241936 335412 241942
rect 335360 241878 335412 241884
rect 336568 241602 336596 244052
rect 337212 241670 337240 244052
rect 337764 242282 337792 244052
rect 337752 242276 337804 242282
rect 337752 242218 337804 242224
rect 337200 241664 337252 241670
rect 337200 241606 337252 241612
rect 336556 241596 336608 241602
rect 336556 241538 336608 241544
rect 338408 241534 338436 244052
rect 338764 242616 338816 242622
rect 338764 242558 338816 242564
rect 338396 241528 338448 241534
rect 338396 241470 338448 241476
rect 338212 16856 338264 16862
rect 338210 16824 338212 16833
rect 338264 16824 338266 16833
rect 338210 16759 338266 16768
rect 337108 4140 337160 4146
rect 337108 4082 337160 4088
rect 333612 3732 333664 3738
rect 333612 3674 333664 3680
rect 335268 3732 335320 3738
rect 335268 3674 335320 3680
rect 333624 480 333652 3674
rect 335912 3664 335964 3670
rect 335912 3606 335964 3612
rect 334716 3392 334768 3398
rect 334716 3334 334768 3340
rect 334728 480 334756 3334
rect 335924 480 335952 3606
rect 337120 480 337148 4082
rect 338304 3596 338356 3602
rect 338304 3538 338356 3544
rect 338316 480 338344 3538
rect 338776 3058 338804 242558
rect 339052 241670 339080 244052
rect 339604 241874 339632 244052
rect 340262 244038 340828 244066
rect 340144 242752 340196 242758
rect 340144 242694 340196 242700
rect 339592 241868 339644 241874
rect 339592 241810 339644 241816
rect 339040 241664 339092 241670
rect 339040 241606 339092 241612
rect 338856 241596 338908 241602
rect 338856 241538 338908 241544
rect 338868 4146 338896 241538
rect 339408 241528 339460 241534
rect 339408 241470 339460 241476
rect 338856 4140 338908 4146
rect 338856 4082 338908 4088
rect 339420 3670 339448 241470
rect 339408 3664 339460 3670
rect 339408 3606 339460 3612
rect 339500 3528 339552 3534
rect 339500 3470 339552 3476
rect 338764 3052 338816 3058
rect 338764 2994 338816 3000
rect 339512 480 339540 3470
rect 340156 3398 340184 242694
rect 340696 40248 340748 40254
rect 340694 40216 340696 40225
rect 340748 40216 340750 40225
rect 340694 40151 340750 40160
rect 340800 3602 340828 244038
rect 340892 241534 340920 244052
rect 341444 242894 341472 244052
rect 341432 242888 341484 242894
rect 341432 242830 341484 242836
rect 341524 242820 341576 242826
rect 341524 242762 341576 242768
rect 340880 241528 340932 241534
rect 340880 241470 340932 241476
rect 340972 40248 341024 40254
rect 340970 40216 340972 40225
rect 341024 40216 341026 40225
rect 340970 40151 341026 40160
rect 340788 3596 340840 3602
rect 340788 3538 340840 3544
rect 340144 3392 340196 3398
rect 340144 3334 340196 3340
rect 340696 3324 340748 3330
rect 340696 3266 340748 3272
rect 340708 480 340736 3266
rect 341536 3194 341564 242762
rect 342088 242690 342116 244052
rect 342076 242684 342128 242690
rect 342076 242626 342128 242632
rect 342732 242078 342760 244052
rect 343284 242758 343312 244052
rect 343272 242752 343324 242758
rect 343272 242694 343324 242700
rect 342904 242412 342956 242418
rect 342904 242354 342956 242360
rect 342720 242072 342772 242078
rect 342720 242014 342772 242020
rect 342628 16856 342680 16862
rect 342626 16824 342628 16833
rect 342680 16824 342682 16833
rect 342626 16759 342682 16768
rect 342916 4146 342944 242354
rect 343928 242146 343956 244052
rect 344586 244038 344968 244066
rect 343916 242140 343968 242146
rect 343916 242082 343968 242088
rect 342904 4140 342956 4146
rect 342904 4082 342956 4088
rect 344284 4140 344336 4146
rect 344284 4082 344336 4088
rect 343088 3460 343140 3466
rect 343088 3402 343140 3408
rect 341524 3188 341576 3194
rect 341524 3130 341576 3136
rect 341892 3052 341944 3058
rect 341892 2994 341944 3000
rect 341904 480 341932 2994
rect 343100 480 343128 3402
rect 344296 480 344324 4082
rect 344940 3466 344968 244038
rect 345124 242826 345152 244052
rect 345112 242820 345164 242826
rect 345112 242762 345164 242768
rect 345664 241732 345716 241738
rect 345664 241674 345716 241680
rect 345676 4146 345704 241674
rect 346228 239306 346256 244174
rect 346320 242894 346348 244052
rect 346964 243234 346992 244052
rect 347622 244038 347728 244066
rect 346952 243228 347004 243234
rect 346952 243170 347004 243176
rect 346308 242888 346360 242894
rect 346308 242830 346360 242836
rect 346228 239278 346348 239306
rect 346320 225010 346348 239278
rect 346124 225004 346176 225010
rect 346124 224946 346176 224952
rect 346308 225004 346360 225010
rect 346308 224946 346360 224952
rect 346136 224890 346164 224946
rect 346136 224862 346256 224890
rect 346228 215370 346256 224862
rect 346228 215342 346348 215370
rect 346320 205698 346348 215342
rect 346124 205692 346176 205698
rect 346124 205634 346176 205640
rect 346308 205692 346360 205698
rect 346308 205634 346360 205640
rect 346136 205578 346164 205634
rect 346136 205550 346256 205578
rect 346228 196058 346256 205550
rect 346228 196030 346348 196058
rect 346320 186386 346348 196030
rect 346124 186380 346176 186386
rect 346124 186322 346176 186328
rect 346308 186380 346360 186386
rect 346308 186322 346360 186328
rect 346136 186266 346164 186322
rect 346136 186238 346256 186266
rect 346228 183569 346256 186238
rect 346030 183560 346086 183569
rect 346030 183495 346086 183504
rect 346214 183560 346270 183569
rect 346214 183495 346270 183504
rect 346044 173942 346072 183495
rect 346032 173936 346084 173942
rect 346032 173878 346084 173884
rect 346308 173936 346360 173942
rect 346308 173878 346360 173884
rect 346320 167074 346348 173878
rect 346124 167068 346176 167074
rect 346124 167010 346176 167016
rect 346308 167068 346360 167074
rect 346308 167010 346360 167016
rect 346136 166954 346164 167010
rect 346136 166926 346256 166954
rect 346228 164218 346256 166926
rect 346216 164212 346268 164218
rect 346216 164154 346268 164160
rect 346216 157344 346268 157350
rect 346216 157286 346268 157292
rect 346228 154578 346256 157286
rect 346228 154550 346348 154578
rect 346320 147694 346348 154550
rect 346124 147688 346176 147694
rect 346308 147688 346360 147694
rect 346176 147636 346256 147642
rect 346124 147630 346256 147636
rect 346308 147630 346360 147636
rect 346136 147614 346256 147630
rect 346228 144906 346256 147614
rect 346216 144900 346268 144906
rect 346216 144842 346268 144848
rect 346216 137964 346268 137970
rect 346216 137906 346268 137912
rect 346228 135266 346256 137906
rect 346228 135238 346348 135266
rect 346320 128382 346348 135238
rect 346124 128376 346176 128382
rect 346308 128376 346360 128382
rect 346176 128324 346256 128330
rect 346124 128318 346256 128324
rect 346308 128318 346360 128324
rect 346136 128302 346256 128318
rect 346228 125594 346256 128302
rect 346216 125588 346268 125594
rect 346216 125530 346268 125536
rect 346216 118652 346268 118658
rect 346216 118594 346268 118600
rect 346228 115954 346256 118594
rect 346228 115926 346348 115954
rect 346320 109070 346348 115926
rect 346124 109064 346176 109070
rect 346308 109064 346360 109070
rect 346176 109012 346256 109018
rect 346124 109006 346256 109012
rect 346308 109006 346360 109012
rect 346136 108990 346256 109006
rect 346228 106282 346256 108990
rect 346216 106276 346268 106282
rect 346216 106218 346268 106224
rect 346216 99340 346268 99346
rect 346216 99282 346268 99288
rect 346228 96642 346256 99282
rect 346228 96614 346348 96642
rect 346320 89758 346348 96614
rect 346124 89752 346176 89758
rect 346308 89752 346360 89758
rect 346176 89700 346256 89706
rect 346124 89694 346256 89700
rect 346308 89694 346360 89700
rect 346136 89678 346256 89694
rect 346228 86970 346256 89678
rect 346216 86964 346268 86970
rect 346216 86906 346268 86912
rect 346308 77308 346360 77314
rect 346308 77250 346360 77256
rect 346320 77217 346348 77250
rect 346122 77208 346178 77217
rect 346122 77143 346178 77152
rect 346306 77208 346362 77217
rect 346306 77143 346362 77152
rect 346136 70446 346164 77143
rect 346124 70440 346176 70446
rect 346124 70382 346176 70388
rect 346216 70372 346268 70378
rect 346216 70314 346268 70320
rect 346228 60738 346256 70314
rect 346228 60710 346348 60738
rect 346320 48346 346348 60710
rect 346216 48340 346268 48346
rect 346216 48282 346268 48288
rect 346308 48340 346360 48346
rect 346308 48282 346360 48288
rect 346228 48226 346256 48282
rect 346136 48198 346256 48226
rect 346136 41426 346164 48198
rect 346136 41398 346256 41426
rect 346228 38706 346256 41398
rect 346136 38678 346256 38706
rect 346136 31822 346164 38678
rect 346124 31816 346176 31822
rect 346124 31758 346176 31764
rect 346216 31680 346268 31686
rect 346216 31622 346268 31628
rect 346228 27606 346256 31622
rect 346216 27600 346268 27606
rect 346216 27542 346268 27548
rect 346216 22092 346268 22098
rect 346216 22034 346268 22040
rect 346228 4214 346256 22034
rect 347700 4282 347728 244038
rect 347964 242480 348016 242486
rect 347964 242422 348016 242428
rect 347688 4276 347740 4282
rect 347688 4218 347740 4224
rect 346216 4208 346268 4214
rect 346216 4150 346268 4156
rect 345664 4140 345716 4146
rect 345664 4082 345716 4088
rect 345480 4004 345532 4010
rect 345480 3946 345532 3952
rect 344928 3460 344980 3466
rect 344928 3402 344980 3408
rect 345492 480 345520 3946
rect 346676 3936 346728 3942
rect 346676 3878 346728 3884
rect 346688 480 346716 3878
rect 347976 626 348004 242422
rect 348160 241534 348188 244052
rect 348804 242214 348832 244052
rect 348792 242208 348844 242214
rect 348792 242150 348844 242156
rect 349448 241738 349476 244052
rect 350000 242486 350028 244052
rect 350658 244038 351040 244066
rect 351302 244038 351776 244066
rect 349988 242480 350040 242486
rect 349988 242422 350040 242428
rect 350816 241936 350868 241942
rect 350816 241878 350868 241884
rect 349436 241732 349488 241738
rect 349436 241674 349488 241680
rect 350448 241732 350500 241738
rect 350448 241674 350500 241680
rect 348148 241528 348200 241534
rect 348148 241470 348200 241476
rect 349068 241528 349120 241534
rect 349068 241470 349120 241476
rect 349080 4078 349108 241470
rect 350460 4350 350488 241674
rect 350448 4344 350500 4350
rect 350448 4286 350500 4292
rect 349068 4072 349120 4078
rect 349068 4014 349120 4020
rect 349068 3392 349120 3398
rect 349068 3334 349120 3340
rect 347884 598 348004 626
rect 347884 480 347912 598
rect 349080 480 349108 3334
rect 350264 3324 350316 3330
rect 350264 3266 350316 3272
rect 350276 480 350304 3266
rect 350828 610 350856 241878
rect 351012 234666 351040 244038
rect 351748 239306 351776 244038
rect 351840 242690 351868 244052
rect 351828 242684 351880 242690
rect 351828 242626 351880 242632
rect 352484 241534 352512 244052
rect 353050 244038 353156 244066
rect 352472 241528 352524 241534
rect 352472 241470 352524 241476
rect 351748 239278 351868 239306
rect 351000 234660 351052 234666
rect 351000 234602 351052 234608
rect 351736 234660 351788 234666
rect 351736 234602 351788 234608
rect 351748 4418 351776 234602
rect 351840 4486 351868 239278
rect 353128 6458 353156 244038
rect 353680 242185 353708 244052
rect 354338 244038 354628 244066
rect 353666 242176 353722 242185
rect 353666 242111 353722 242120
rect 353208 241528 353260 241534
rect 353208 241470 353260 241476
rect 353116 6452 353168 6458
rect 353116 6394 353168 6400
rect 353220 4622 353248 241470
rect 354600 4690 354628 244038
rect 354876 241534 354904 244052
rect 355534 244038 356008 244066
rect 355232 242344 355284 242350
rect 355508 242344 355560 242350
rect 355284 242292 355508 242298
rect 355232 242286 355560 242292
rect 355244 242270 355548 242286
rect 354772 241528 354824 241534
rect 354772 241470 354824 241476
rect 354864 241528 354916 241534
rect 354864 241470 354916 241476
rect 355876 241528 355928 241534
rect 355876 241470 355928 241476
rect 354784 241346 354812 241470
rect 354784 241318 354904 241346
rect 354588 4684 354640 4690
rect 354588 4626 354640 4632
rect 353208 4616 353260 4622
rect 353208 4558 353260 4564
rect 351828 4480 351880 4486
rect 351828 4422 351880 4428
rect 351736 4412 351788 4418
rect 351736 4354 351788 4360
rect 352564 3868 352616 3874
rect 352564 3810 352616 3816
rect 350816 604 350868 610
rect 350816 546 350868 552
rect 351368 604 351420 610
rect 351368 546 351420 552
rect 351380 480 351408 546
rect 352576 480 352604 3810
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 353772 480 353800 3334
rect 354876 626 354904 241318
rect 355888 6390 355916 241470
rect 355876 6384 355928 6390
rect 355876 6326 355928 6332
rect 355980 4010 356008 244038
rect 356164 241534 356192 244052
rect 356730 244038 357112 244066
rect 357084 241602 357112 244038
rect 357360 242554 357388 244052
rect 357348 242548 357400 242554
rect 357348 242490 357400 242496
rect 357530 242312 357586 242321
rect 357440 242276 357492 242282
rect 357530 242247 357586 242256
rect 357440 242218 357492 242224
rect 357452 242162 357480 242218
rect 357544 242162 357572 242247
rect 357452 242134 357572 242162
rect 357440 241732 357492 241738
rect 357440 241674 357492 241680
rect 356704 241596 356756 241602
rect 356704 241538 356756 241544
rect 357072 241596 357124 241602
rect 357072 241538 357124 241544
rect 356152 241528 356204 241534
rect 356152 241470 356204 241476
rect 356336 241460 356388 241466
rect 356336 241402 356388 241408
rect 356348 12442 356376 241402
rect 356336 12436 356388 12442
rect 356336 12378 356388 12384
rect 355968 4004 356020 4010
rect 355968 3946 356020 3952
rect 356716 3806 356744 241538
rect 357348 241528 357400 241534
rect 357348 241470 357400 241476
rect 357360 225010 357388 241470
rect 357164 225004 357216 225010
rect 357164 224946 357216 224952
rect 357348 225004 357400 225010
rect 357348 224946 357400 224952
rect 357176 224890 357204 224946
rect 357176 224862 357296 224890
rect 357268 215370 357296 224862
rect 357268 215342 357388 215370
rect 357360 205698 357388 215342
rect 357164 205692 357216 205698
rect 357164 205634 357216 205640
rect 357348 205692 357400 205698
rect 357348 205634 357400 205640
rect 357176 205578 357204 205634
rect 357176 205550 357296 205578
rect 357268 196058 357296 205550
rect 357268 196030 357388 196058
rect 357360 186386 357388 196030
rect 357164 186380 357216 186386
rect 357164 186322 357216 186328
rect 357348 186380 357400 186386
rect 357348 186322 357400 186328
rect 357176 186266 357204 186322
rect 357176 186238 357296 186266
rect 357268 183569 357296 186238
rect 357070 183560 357126 183569
rect 357070 183495 357126 183504
rect 357254 183560 357310 183569
rect 357254 183495 357310 183504
rect 357084 173942 357112 183495
rect 357072 173936 357124 173942
rect 357072 173878 357124 173884
rect 357348 173936 357400 173942
rect 357348 173878 357400 173884
rect 357360 167074 357388 173878
rect 357164 167068 357216 167074
rect 357164 167010 357216 167016
rect 357348 167068 357400 167074
rect 357348 167010 357400 167016
rect 357176 166954 357204 167010
rect 357176 166926 357296 166954
rect 357268 164218 357296 166926
rect 357256 164212 357308 164218
rect 357256 164154 357308 164160
rect 357256 157344 357308 157350
rect 357256 157286 357308 157292
rect 357268 154578 357296 157286
rect 357268 154550 357388 154578
rect 357360 147694 357388 154550
rect 357164 147688 357216 147694
rect 357348 147688 357400 147694
rect 357216 147636 357296 147642
rect 357164 147630 357296 147636
rect 357348 147630 357400 147636
rect 357176 147614 357296 147630
rect 357268 144906 357296 147614
rect 357256 144900 357308 144906
rect 357256 144842 357308 144848
rect 357256 137964 357308 137970
rect 357256 137906 357308 137912
rect 357268 135266 357296 137906
rect 357268 135238 357388 135266
rect 357360 128382 357388 135238
rect 357164 128376 357216 128382
rect 357348 128376 357400 128382
rect 357216 128324 357296 128330
rect 357164 128318 357296 128324
rect 357348 128318 357400 128324
rect 357176 128302 357296 128318
rect 357268 125594 357296 128302
rect 357256 125588 357308 125594
rect 357256 125530 357308 125536
rect 357256 118652 357308 118658
rect 357256 118594 357308 118600
rect 357268 115954 357296 118594
rect 357268 115926 357388 115954
rect 357360 109070 357388 115926
rect 357164 109064 357216 109070
rect 357348 109064 357400 109070
rect 357216 109012 357296 109018
rect 357164 109006 357296 109012
rect 357348 109006 357400 109012
rect 357176 108990 357296 109006
rect 357268 106282 357296 108990
rect 357256 106276 357308 106282
rect 357256 106218 357308 106224
rect 357256 99340 357308 99346
rect 357256 99282 357308 99288
rect 357268 96642 357296 99282
rect 357268 96614 357388 96642
rect 357360 89758 357388 96614
rect 357164 89752 357216 89758
rect 357348 89752 357400 89758
rect 357216 89700 357296 89706
rect 357164 89694 357296 89700
rect 357348 89694 357400 89700
rect 357176 89678 357296 89694
rect 357268 86970 357296 89678
rect 357256 86964 357308 86970
rect 357256 86906 357308 86912
rect 357348 77308 357400 77314
rect 357348 77250 357400 77256
rect 357360 77178 357388 77250
rect 357348 77172 357400 77178
rect 357348 77114 357400 77120
rect 357256 67652 357308 67658
rect 357256 67594 357308 67600
rect 357268 60738 357296 67594
rect 357268 60710 357388 60738
rect 357360 57934 357388 60710
rect 357348 57928 357400 57934
rect 357348 57870 357400 57876
rect 357256 48340 357308 48346
rect 357256 48282 357308 48288
rect 357268 41426 357296 48282
rect 357268 41398 357388 41426
rect 357360 38622 357388 41398
rect 357348 38616 357400 38622
rect 357348 38558 357400 38564
rect 357256 31748 357308 31754
rect 357256 31690 357308 31696
rect 357268 22114 357296 31690
rect 357268 22086 357388 22114
rect 357360 12458 357388 22086
rect 357176 12430 357388 12458
rect 357452 12442 357480 241674
rect 358004 241534 358032 244052
rect 358570 244038 358676 244066
rect 358084 241664 358136 241670
rect 358084 241606 358136 241612
rect 357992 241528 358044 241534
rect 357992 241470 358044 241476
rect 357440 12436 357492 12442
rect 357176 4554 357204 12430
rect 357440 12378 357492 12384
rect 357348 12368 357400 12374
rect 357348 12310 357400 12316
rect 357164 4548 357216 4554
rect 357164 4490 357216 4496
rect 356152 3800 356204 3806
rect 356152 3742 356204 3748
rect 356704 3800 356756 3806
rect 356704 3742 356756 3748
rect 354876 598 354996 626
rect 354968 480 354996 598
rect 356164 480 356192 3742
rect 357360 480 357388 12310
rect 358096 3330 358124 241606
rect 358544 12436 358596 12442
rect 358544 12378 358596 12384
rect 358084 3324 358136 3330
rect 358084 3266 358136 3272
rect 358556 480 358584 12378
rect 358648 6322 358676 244038
rect 359200 241534 359228 244052
rect 359858 244038 360056 244066
rect 359464 242480 359516 242486
rect 359464 242422 359516 242428
rect 358728 241528 358780 241534
rect 358728 241470 358780 241476
rect 359188 241528 359240 241534
rect 359188 241470 359240 241476
rect 358636 6316 358688 6322
rect 358636 6258 358688 6264
rect 358740 4758 358768 241470
rect 358728 4752 358780 4758
rect 358728 4694 358780 4700
rect 359476 3398 359504 242422
rect 359922 40216 359978 40225
rect 359922 40151 359924 40160
rect 359976 40151 359978 40160
rect 359924 40122 359976 40128
rect 359924 16856 359976 16862
rect 359922 16824 359924 16833
rect 359976 16824 359978 16833
rect 359922 16759 359978 16768
rect 360028 5438 360056 244038
rect 360396 241670 360424 244052
rect 361040 242350 361068 244052
rect 361028 242344 361080 242350
rect 361028 242286 361080 242292
rect 360384 241664 360436 241670
rect 360384 241606 360436 241612
rect 361592 241534 361620 244052
rect 362250 244038 362724 244066
rect 361856 242480 361908 242486
rect 361856 242422 361908 242428
rect 360108 241528 360160 241534
rect 360108 241470 360160 241476
rect 361580 241528 361632 241534
rect 361580 241470 361632 241476
rect 360016 5432 360068 5438
rect 360016 5374 360068 5380
rect 360120 3942 360148 241470
rect 360198 40216 360254 40225
rect 360198 40151 360200 40160
rect 360252 40151 360254 40160
rect 360200 40122 360252 40128
rect 360936 4140 360988 4146
rect 360936 4082 360988 4088
rect 360108 3936 360160 3942
rect 360108 3878 360160 3884
rect 359740 3732 359792 3738
rect 359740 3674 359792 3680
rect 359464 3392 359516 3398
rect 359464 3334 359516 3340
rect 359752 480 359780 3674
rect 360948 480 360976 4082
rect 361868 610 361896 242422
rect 362224 16856 362276 16862
rect 362222 16824 362224 16833
rect 362276 16824 362278 16833
rect 362222 16759 362278 16768
rect 362696 6254 362724 244038
rect 362776 241528 362828 241534
rect 362776 241470 362828 241476
rect 362684 6248 362736 6254
rect 362684 6190 362736 6196
rect 362788 5506 362816 241470
rect 362776 5500 362828 5506
rect 362776 5442 362828 5448
rect 362880 3874 362908 244052
rect 363432 241534 363460 244052
rect 364090 244038 364196 244066
rect 363420 241528 363472 241534
rect 363420 241470 363472 241476
rect 364168 6186 364196 244038
rect 364720 242826 364748 244052
rect 365286 244038 365668 244066
rect 364708 242820 364760 242826
rect 364708 242762 364760 242768
rect 364248 241528 364300 241534
rect 364248 241470 364300 241476
rect 364156 6180 364208 6186
rect 364156 6122 364208 6128
rect 364260 5370 364288 241470
rect 364248 5364 364300 5370
rect 364248 5306 364300 5312
rect 365640 5302 365668 244038
rect 365812 241800 365864 241806
rect 365812 241742 365864 241748
rect 365628 5296 365680 5302
rect 365628 5238 365680 5244
rect 362868 3868 362920 3874
rect 362868 3810 362920 3816
rect 364524 3800 364576 3806
rect 364524 3742 364576 3748
rect 363328 3664 363380 3670
rect 363328 3606 363380 3612
rect 361856 604 361908 610
rect 361856 546 361908 552
rect 362132 604 362184 610
rect 362132 546 362184 552
rect 362144 480 362172 546
rect 363340 480 363368 3606
rect 364536 480 364564 3742
rect 365824 626 365852 241742
rect 365916 241534 365944 244052
rect 366574 244038 366956 244066
rect 367126 244038 367416 244066
rect 365904 241528 365956 241534
rect 365904 241470 365956 241476
rect 366928 3738 366956 244038
rect 367098 242720 367154 242729
rect 367098 242655 367100 242664
rect 367152 242655 367154 242664
rect 367100 242626 367152 242632
rect 367098 242584 367154 242593
rect 367098 242519 367100 242528
rect 367152 242519 367154 242528
rect 367100 242490 367152 242496
rect 367190 242448 367246 242457
rect 367020 242392 367190 242400
rect 367020 242383 367246 242392
rect 367020 242372 367232 242383
rect 367020 242321 367048 242372
rect 367006 242312 367062 242321
rect 367006 242247 367062 242256
rect 367388 241806 367416 244038
rect 367756 242962 367784 244052
rect 367744 242956 367796 242962
rect 367744 242898 367796 242904
rect 367652 242684 367704 242690
rect 367652 242626 367704 242632
rect 367466 242584 367522 242593
rect 367466 242519 367468 242528
rect 367520 242519 367522 242528
rect 367468 242490 367520 242496
rect 367376 241800 367428 241806
rect 367664 241777 367692 242626
rect 368400 242282 368428 244052
rect 368952 243098 368980 244052
rect 369610 244038 369716 244066
rect 368940 243092 368992 243098
rect 368940 243034 368992 243040
rect 369582 242448 369638 242457
rect 369582 242383 369584 242392
rect 369636 242383 369638 242392
rect 369584 242354 369636 242360
rect 368388 242276 368440 242282
rect 368388 242218 368440 242224
rect 368480 241868 368532 241874
rect 368480 241810 368532 241816
rect 368388 241800 368440 241806
rect 367376 241742 367428 241748
rect 367650 241768 367706 241777
rect 368388 241742 368440 241748
rect 367650 241703 367706 241712
rect 367008 241528 367060 241534
rect 367008 241470 367060 241476
rect 367020 3806 367048 241470
rect 368400 5234 368428 241742
rect 368388 5228 368440 5234
rect 368388 5170 368440 5176
rect 367008 3800 367060 3806
rect 367008 3742 367060 3748
rect 366916 3732 366968 3738
rect 366916 3674 366968 3680
rect 366916 3596 366968 3602
rect 366916 3538 366968 3544
rect 365732 598 365852 626
rect 365732 480 365760 598
rect 366928 480 366956 3538
rect 368020 3324 368072 3330
rect 368020 3266 368072 3272
rect 368032 480 368060 3266
rect 368492 610 368520 241810
rect 369124 241800 369176 241806
rect 369124 241742 369176 241748
rect 369136 241670 369164 241742
rect 369124 241664 369176 241670
rect 369124 241606 369176 241612
rect 369688 7682 369716 244038
rect 369768 243092 369820 243098
rect 369768 243034 369820 243040
rect 369676 7676 369728 7682
rect 369676 7618 369728 7624
rect 369780 5166 369808 243034
rect 370148 242826 370176 244052
rect 370806 244038 371096 244066
rect 370136 242820 370188 242826
rect 370136 242762 370188 242768
rect 369768 5160 369820 5166
rect 369768 5102 369820 5108
rect 371068 5098 371096 244038
rect 371148 242820 371200 242826
rect 371148 242762 371200 242768
rect 371056 5092 371108 5098
rect 371056 5034 371108 5040
rect 371160 3670 371188 242762
rect 371436 241874 371464 244052
rect 372002 244038 372568 244066
rect 371424 241868 371476 241874
rect 371424 241810 371476 241816
rect 371148 3664 371200 3670
rect 371148 3606 371200 3612
rect 372540 3602 372568 244038
rect 372632 241534 372660 244052
rect 373290 244038 373764 244066
rect 373842 244038 373948 244066
rect 372804 242004 372856 242010
rect 372804 241946 372856 241952
rect 372620 241528 372672 241534
rect 372620 241470 372672 241476
rect 372816 241346 372844 241946
rect 372632 241318 372844 241346
rect 372528 3596 372580 3602
rect 372528 3538 372580 3544
rect 370412 3528 370464 3534
rect 370412 3470 370464 3476
rect 368480 604 368532 610
rect 368480 546 368532 552
rect 369216 604 369268 610
rect 369216 546 369268 552
rect 369228 480 369256 546
rect 370424 480 370452 3470
rect 371608 3392 371660 3398
rect 371608 3334 371660 3340
rect 371620 480 371648 3334
rect 372632 610 372660 241318
rect 373736 7478 373764 244038
rect 373816 241528 373868 241534
rect 373816 241470 373868 241476
rect 373724 7472 373776 7478
rect 373724 7414 373776 7420
rect 373828 5030 373856 241470
rect 373816 5024 373868 5030
rect 373816 4966 373868 4972
rect 373920 3534 373948 244038
rect 374274 242720 374330 242729
rect 374274 242655 374330 242664
rect 374288 242146 374316 242655
rect 374276 242140 374328 242146
rect 374276 242082 374328 242088
rect 374092 242072 374144 242078
rect 374092 242014 374144 242020
rect 373908 3528 373960 3534
rect 373908 3470 373960 3476
rect 374104 1562 374132 242014
rect 374274 241530 374330 241539
rect 374472 241534 374500 244052
rect 375116 242010 375144 244052
rect 375668 242826 375696 244052
rect 376326 244038 376708 244066
rect 375656 242820 375708 242826
rect 375656 242762 375708 242768
rect 376024 242072 376076 242078
rect 376024 242014 376076 242020
rect 375104 242004 375156 242010
rect 375104 241946 375156 241952
rect 375564 241596 375616 241602
rect 375564 241538 375616 241544
rect 374274 241465 374330 241474
rect 374460 241528 374512 241534
rect 374460 241470 374512 241476
rect 375288 241528 375340 241534
rect 375288 241470 375340 241476
rect 374288 240145 374316 241465
rect 374274 240136 374330 240145
rect 374274 240071 374330 240080
rect 374458 240136 374514 240145
rect 374458 240071 374514 240080
rect 374472 230518 374500 240071
rect 374276 230512 374328 230518
rect 374276 230454 374328 230460
rect 374460 230512 374512 230518
rect 374460 230454 374512 230460
rect 374288 220833 374316 230454
rect 374274 220824 374330 220833
rect 374274 220759 374330 220768
rect 374458 220824 374514 220833
rect 374458 220759 374514 220768
rect 374472 211177 374500 220759
rect 374274 211168 374330 211177
rect 374274 211103 374330 211112
rect 374458 211168 374514 211177
rect 374458 211103 374514 211112
rect 374288 201482 374316 211103
rect 374276 201476 374328 201482
rect 374276 201418 374328 201424
rect 374460 201476 374512 201482
rect 374460 201418 374512 201424
rect 374472 191865 374500 201418
rect 374274 191856 374330 191865
rect 374274 191791 374330 191800
rect 374458 191856 374514 191865
rect 374458 191791 374514 191800
rect 374288 182170 374316 191791
rect 374276 182164 374328 182170
rect 374276 182106 374328 182112
rect 374460 182164 374512 182170
rect 374460 182106 374512 182112
rect 374472 172553 374500 182106
rect 374274 172544 374330 172553
rect 374274 172479 374330 172488
rect 374458 172544 374514 172553
rect 374458 172479 374514 172488
rect 374288 162858 374316 172479
rect 374276 162852 374328 162858
rect 374276 162794 374328 162800
rect 374276 153264 374328 153270
rect 374276 153206 374328 153212
rect 374288 143546 374316 153206
rect 374276 143540 374328 143546
rect 374276 143482 374328 143488
rect 374276 133952 374328 133958
rect 374276 133894 374328 133900
rect 374288 124166 374316 133894
rect 374276 124160 374328 124166
rect 374276 124102 374328 124108
rect 374276 114572 374328 114578
rect 374276 114514 374328 114520
rect 374288 104854 374316 114514
rect 374276 104848 374328 104854
rect 374276 104790 374328 104796
rect 374276 95260 374328 95266
rect 374276 95202 374328 95208
rect 374288 85542 374316 95202
rect 374276 85536 374328 85542
rect 374276 85478 374328 85484
rect 374276 75948 374328 75954
rect 374276 75890 374328 75896
rect 374288 66230 374316 75890
rect 374276 66224 374328 66230
rect 374276 66166 374328 66172
rect 374276 56636 374328 56642
rect 374276 56578 374328 56584
rect 374288 46918 374316 56578
rect 374276 46912 374328 46918
rect 374276 46854 374328 46860
rect 374276 37324 374328 37330
rect 374276 37266 374328 37272
rect 374288 27606 374316 37266
rect 374276 27600 374328 27606
rect 374276 27542 374328 27548
rect 374276 18012 374328 18018
rect 374276 17954 374328 17960
rect 374288 12578 374316 17954
rect 374276 12572 374328 12578
rect 374276 12514 374328 12520
rect 374184 9716 374236 9722
rect 374184 9658 374236 9664
rect 374196 9602 374224 9658
rect 374196 9574 374316 9602
rect 374288 2718 374316 9574
rect 375300 4962 375328 241470
rect 375576 12442 375604 241538
rect 375564 12436 375616 12442
rect 375564 12378 375616 12384
rect 375288 4956 375340 4962
rect 375288 4898 375340 4904
rect 376036 4146 376064 242014
rect 376392 12436 376444 12442
rect 376392 12378 376444 12384
rect 376024 4140 376076 4146
rect 376024 4082 376076 4088
rect 374276 2712 374328 2718
rect 374276 2654 374328 2660
rect 374092 1556 374144 1562
rect 374092 1498 374144 1504
rect 375196 1556 375248 1562
rect 375196 1498 375248 1504
rect 372620 604 372672 610
rect 372620 546 372672 552
rect 372804 604 372856 610
rect 372804 546 372856 552
rect 374000 604 374052 610
rect 374000 546 374052 552
rect 372816 480 372844 546
rect 374012 480 374040 546
rect 375208 480 375236 1498
rect 376404 480 376432 12378
rect 376680 4826 376708 244038
rect 376956 242690 376984 244052
rect 377404 242888 377456 242894
rect 377404 242830 377456 242836
rect 376944 242684 376996 242690
rect 376944 242626 376996 242632
rect 376668 4820 376720 4826
rect 376668 4762 376720 4768
rect 377416 3126 377444 242830
rect 377508 241670 377536 244052
rect 378152 242758 378180 244052
rect 378718 244038 379008 244066
rect 378140 242752 378192 242758
rect 378140 242694 378192 242700
rect 377496 241664 377548 241670
rect 377496 241606 377548 241612
rect 378980 235498 379008 244038
rect 379348 242078 379376 244052
rect 379428 242752 379480 242758
rect 379428 242694 379480 242700
rect 379336 242072 379388 242078
rect 379336 242014 379388 242020
rect 378888 235470 379008 235498
rect 378888 230761 378916 235470
rect 378874 230752 378930 230761
rect 378874 230687 378930 230696
rect 379242 230480 379298 230489
rect 379242 230415 379298 230424
rect 379072 220862 379100 220893
rect 379256 220862 379284 230415
rect 379060 220856 379112 220862
rect 379244 220856 379296 220862
rect 379112 220804 379192 220810
rect 379060 220798 379192 220804
rect 379244 220798 379296 220804
rect 379072 220794 379192 220798
rect 379072 220788 379204 220794
rect 379072 220782 379152 220788
rect 379152 220730 379204 220736
rect 379336 220788 379388 220794
rect 379336 220730 379388 220736
rect 379348 211154 379376 220730
rect 379164 211138 379376 211154
rect 379152 211132 379376 211138
rect 379204 211126 379244 211132
rect 379152 211074 379204 211080
rect 379296 211126 379376 211132
rect 379244 211074 379296 211080
rect 379164 211043 379192 211074
rect 379256 201521 379284 211074
rect 379058 201512 379114 201521
rect 379058 201447 379114 201456
rect 379242 201512 379298 201521
rect 379242 201447 379298 201456
rect 379072 193202 379100 201447
rect 378888 193174 379100 193202
rect 378888 183666 378916 193174
rect 378876 183660 378928 183666
rect 378876 183602 378928 183608
rect 379060 183660 379112 183666
rect 379060 183602 379112 183608
rect 379072 182170 379100 183602
rect 379060 182164 379112 182170
rect 379060 182106 379112 182112
rect 379336 182164 379388 182170
rect 379336 182106 379388 182112
rect 379348 164286 379376 182106
rect 379152 164280 379204 164286
rect 379072 164228 379152 164234
rect 379072 164222 379204 164228
rect 379336 164280 379388 164286
rect 379336 164222 379388 164228
rect 379072 164206 379192 164222
rect 379072 162858 379100 164206
rect 379060 162852 379112 162858
rect 379060 162794 379112 162800
rect 379060 157344 379112 157350
rect 379060 157286 379112 157292
rect 379072 153218 379100 157286
rect 379072 153190 379192 153218
rect 379164 144974 379192 153190
rect 379152 144968 379204 144974
rect 379152 144910 379204 144916
rect 379152 144832 379204 144838
rect 379152 144774 379204 144780
rect 379164 142118 379192 144774
rect 379152 142112 379204 142118
rect 379152 142054 379204 142060
rect 379244 132524 379296 132530
rect 379244 132466 379296 132472
rect 379256 132394 379284 132466
rect 379244 132388 379296 132394
rect 379244 132330 379296 132336
rect 379152 122868 379204 122874
rect 379152 122810 379204 122816
rect 379164 100094 379192 122810
rect 379152 100088 379204 100094
rect 379152 100030 379204 100036
rect 379152 89412 379204 89418
rect 379152 89354 379204 89360
rect 379164 66230 379192 89354
rect 379152 66224 379204 66230
rect 379152 66166 379204 66172
rect 379152 56704 379204 56710
rect 379152 56646 379204 56652
rect 379164 56574 379192 56646
rect 379152 56568 379204 56574
rect 379152 56510 379204 56516
rect 379244 46980 379296 46986
rect 379244 46922 379296 46928
rect 379256 37330 379284 46922
rect 379152 37324 379204 37330
rect 379152 37266 379204 37272
rect 379244 37324 379296 37330
rect 379244 37266 379296 37272
rect 379164 37233 379192 37266
rect 379150 37224 379206 37233
rect 379150 37159 379206 37168
rect 379334 37224 379390 37233
rect 379334 37159 379390 37168
rect 379348 31822 379376 37159
rect 379336 31816 379388 31822
rect 379336 31758 379388 31764
rect 379244 31680 379296 31686
rect 379244 31622 379296 31628
rect 379256 27538 379284 31622
rect 379244 27532 379296 27538
rect 379244 27474 379296 27480
rect 379336 22092 379388 22098
rect 379336 22034 379388 22040
rect 379244 16856 379296 16862
rect 379242 16824 379244 16833
rect 379296 16824 379298 16833
rect 379242 16759 379298 16768
rect 379348 14498 379376 22034
rect 379256 14470 379376 14498
rect 379256 7002 379284 14470
rect 379244 6996 379296 7002
rect 379244 6938 379296 6944
rect 379336 5024 379388 5030
rect 379334 4992 379336 5001
rect 379388 4992 379390 5001
rect 379334 4927 379390 4936
rect 379440 4894 379468 242694
rect 379704 242616 379756 242622
rect 379704 242558 379756 242564
rect 379612 16856 379664 16862
rect 379610 16824 379612 16833
rect 379664 16824 379666 16833
rect 379610 16759 379666 16768
rect 379520 5024 379572 5030
rect 379518 4992 379520 5001
rect 379572 4992 379574 5001
rect 379518 4927 379574 4936
rect 379428 4888 379480 4894
rect 379428 4830 379480 4836
rect 377588 4140 377640 4146
rect 377588 4082 377640 4088
rect 377404 3120 377456 3126
rect 377404 3062 377456 3068
rect 377600 480 377628 4082
rect 378784 3460 378836 3466
rect 378784 3402 378836 3408
rect 378796 480 378824 3402
rect 379716 610 379744 242558
rect 379992 241534 380020 244052
rect 380558 244038 380756 244066
rect 380164 241936 380216 241942
rect 380164 241878 380216 241884
rect 379980 241528 380032 241534
rect 379980 241470 380032 241476
rect 380176 3330 380204 241878
rect 380256 241664 380308 241670
rect 380256 241606 380308 241612
rect 380164 3324 380216 3330
rect 380164 3266 380216 3272
rect 380268 3262 380296 241606
rect 380728 9450 380756 244038
rect 381188 241602 381216 244052
rect 381846 244038 382228 244066
rect 381176 241596 381228 241602
rect 381176 241538 381228 241544
rect 380808 241528 380860 241534
rect 380808 241470 380860 241476
rect 380716 9444 380768 9450
rect 380716 9386 380768 9392
rect 380820 4865 380848 241470
rect 380806 4856 380862 4865
rect 380806 4791 380862 4800
rect 382200 4214 382228 244038
rect 382384 241534 382412 244052
rect 382464 242412 382516 242418
rect 382464 242354 382516 242360
rect 382372 241528 382424 241534
rect 382372 241470 382424 241476
rect 381176 4208 381228 4214
rect 381176 4150 381228 4156
rect 382188 4208 382240 4214
rect 382188 4150 382240 4156
rect 380256 3256 380308 3262
rect 380256 3198 380308 3204
rect 379704 604 379756 610
rect 379704 546 379756 552
rect 379980 604 380032 610
rect 379980 546 380032 552
rect 379992 480 380020 546
rect 381188 480 381216 4150
rect 382372 3120 382424 3126
rect 382372 3062 382424 3068
rect 382384 480 382412 3062
rect 382476 610 382504 242354
rect 383028 241670 383056 244052
rect 383016 241664 383068 241670
rect 383016 241606 383068 241612
rect 383672 241534 383700 244052
rect 384238 244038 384620 244066
rect 384304 242140 384356 242146
rect 384304 242082 384356 242088
rect 383568 241528 383620 241534
rect 383568 241470 383620 241476
rect 383660 241528 383712 241534
rect 383660 241470 383712 241476
rect 383580 9518 383608 241470
rect 383568 9512 383620 9518
rect 383568 9454 383620 9460
rect 384316 3194 384344 242082
rect 384488 241800 384540 241806
rect 384488 241742 384540 241748
rect 384396 241596 384448 241602
rect 384396 241538 384448 241544
rect 384408 124166 384436 241538
rect 384500 124166 384528 241742
rect 384592 237266 384620 244038
rect 384868 242146 384896 244052
rect 384856 242140 384908 242146
rect 384856 242082 384908 242088
rect 385420 241534 385448 244052
rect 386078 244038 386276 244066
rect 385684 242684 385736 242690
rect 385684 242626 385736 242632
rect 384948 241528 385000 241534
rect 384948 241470 385000 241476
rect 385408 241528 385460 241534
rect 385408 241470 385460 241476
rect 384592 237238 384712 237266
rect 384684 230489 384712 237238
rect 384670 230480 384726 230489
rect 384670 230415 384726 230424
rect 384854 230480 384910 230489
rect 384854 230415 384910 230424
rect 384592 220862 384620 220893
rect 384868 220862 384896 230415
rect 384580 220856 384632 220862
rect 384856 220856 384908 220862
rect 384632 220804 384712 220810
rect 384580 220798 384712 220804
rect 384856 220798 384908 220804
rect 384592 220782 384712 220798
rect 384684 220674 384712 220782
rect 384592 220646 384712 220674
rect 384592 211154 384620 220646
rect 384592 211138 384712 211154
rect 384592 211132 384724 211138
rect 384592 211126 384672 211132
rect 384672 211074 384724 211080
rect 384684 211043 384712 211074
rect 384672 205624 384724 205630
rect 384672 205566 384724 205572
rect 384684 183666 384712 205566
rect 384580 183660 384632 183666
rect 384580 183602 384632 183608
rect 384672 183660 384724 183666
rect 384672 183602 384724 183608
rect 384592 182170 384620 183602
rect 384580 182164 384632 182170
rect 384580 182106 384632 182112
rect 384580 176656 384632 176662
rect 384580 176598 384632 176604
rect 384592 164370 384620 176598
rect 384592 164342 384712 164370
rect 384684 164234 384712 164342
rect 384592 164206 384712 164234
rect 384592 162858 384620 164206
rect 384580 162852 384632 162858
rect 384580 162794 384632 162800
rect 384580 153264 384632 153270
rect 384580 153206 384632 153212
rect 384592 144838 384620 153206
rect 384580 144832 384632 144838
rect 384580 144774 384632 144780
rect 384856 144832 384908 144838
rect 384856 144774 384908 144780
rect 384868 135289 384896 144774
rect 384670 135280 384726 135289
rect 384670 135215 384726 135224
rect 384854 135280 384910 135289
rect 384854 135215 384910 135224
rect 384684 133890 384712 135215
rect 384672 133884 384724 133890
rect 384672 133826 384724 133832
rect 384672 127832 384724 127838
rect 384672 127774 384724 127780
rect 384396 124160 384448 124166
rect 384396 124102 384448 124108
rect 384488 124160 384540 124166
rect 384488 124102 384540 124108
rect 384488 124024 384540 124030
rect 384488 123966 384540 123972
rect 384396 123956 384448 123962
rect 384396 123898 384448 123904
rect 384304 3188 384356 3194
rect 384304 3130 384356 3136
rect 384408 2990 384436 123898
rect 384500 8378 384528 123966
rect 384684 114578 384712 127774
rect 384580 114572 384632 114578
rect 384580 114514 384632 114520
rect 384672 114572 384724 114578
rect 384672 114514 384724 114520
rect 384592 114442 384620 114514
rect 384580 114436 384632 114442
rect 384580 114378 384632 114384
rect 384856 104916 384908 104922
rect 384856 104858 384908 104864
rect 384868 96665 384896 104858
rect 384670 96656 384726 96665
rect 384670 96591 384672 96600
rect 384724 96591 384726 96600
rect 384854 96656 384910 96665
rect 384854 96591 384856 96600
rect 384672 96562 384724 96568
rect 384908 96591 384910 96600
rect 384856 96562 384908 96568
rect 384868 87009 384896 96562
rect 384670 87000 384726 87009
rect 384670 86935 384726 86944
rect 384854 87000 384910 87009
rect 384854 86935 384910 86944
rect 384684 75886 384712 86935
rect 384672 75880 384724 75886
rect 384672 75822 384724 75828
rect 384764 66292 384816 66298
rect 384764 66234 384816 66240
rect 384776 61418 384804 66234
rect 384776 61390 384896 61418
rect 384868 48346 384896 61390
rect 384764 48340 384816 48346
rect 384764 48282 384816 48288
rect 384856 48340 384908 48346
rect 384856 48282 384908 48288
rect 384776 38690 384804 48282
rect 384672 38684 384724 38690
rect 384672 38626 384724 38632
rect 384764 38684 384816 38690
rect 384764 38626 384816 38632
rect 384684 31754 384712 38626
rect 384672 31748 384724 31754
rect 384672 31690 384724 31696
rect 384856 31748 384908 31754
rect 384856 31690 384908 31696
rect 384868 27606 384896 31690
rect 384856 27600 384908 27606
rect 384856 27542 384908 27548
rect 384580 18012 384632 18018
rect 384580 17954 384632 17960
rect 384592 9722 384620 17954
rect 384580 9716 384632 9722
rect 384580 9658 384632 9664
rect 384856 9716 384908 9722
rect 384856 9658 384908 9664
rect 384868 9382 384896 9658
rect 384856 9376 384908 9382
rect 384856 9318 384908 9324
rect 384500 8350 384896 8378
rect 384672 4276 384724 4282
rect 384672 4218 384724 4224
rect 384396 2984 384448 2990
rect 384396 2926 384448 2932
rect 382464 604 382516 610
rect 382464 546 382516 552
rect 383568 604 383620 610
rect 383568 546 383620 552
rect 383580 480 383608 546
rect 384684 480 384712 4218
rect 384868 4214 384896 8350
rect 384960 5574 384988 241470
rect 384948 5568 385000 5574
rect 384948 5510 385000 5516
rect 384856 4208 384908 4214
rect 384856 4150 384908 4156
rect 385696 4146 385724 242626
rect 386248 9314 386276 244038
rect 386708 241602 386736 244052
rect 387274 244038 387748 244066
rect 386696 241596 386748 241602
rect 386696 241538 386748 241544
rect 386328 241528 386380 241534
rect 386328 241470 386380 241476
rect 386236 9308 386288 9314
rect 386236 9250 386288 9256
rect 386340 5642 386368 241470
rect 387720 5710 387748 244038
rect 387904 241534 387932 244052
rect 388442 242176 388498 242185
rect 388442 242111 388498 242120
rect 387892 241528 387944 241534
rect 387892 241470 387944 241476
rect 387708 5704 387760 5710
rect 387708 5646 387760 5652
rect 386328 5636 386380 5642
rect 386328 5578 386380 5584
rect 388260 4344 388312 4350
rect 388260 4286 388312 4292
rect 385684 4140 385736 4146
rect 385684 4082 385736 4088
rect 387064 4140 387116 4146
rect 387064 4082 387116 4088
rect 385868 4072 385920 4078
rect 385868 4014 385920 4020
rect 385880 480 385908 4014
rect 387076 480 387104 4082
rect 388272 480 388300 4286
rect 388456 3058 388484 242111
rect 388548 241874 388576 244052
rect 388628 242208 388680 242214
rect 388628 242150 388680 242156
rect 388536 241868 388588 241874
rect 388536 241810 388588 241816
rect 388536 241596 388588 241602
rect 388536 241538 388588 241544
rect 388548 3126 388576 241538
rect 388640 4282 388668 242150
rect 388996 241528 389048 241534
rect 388996 241470 389048 241476
rect 389008 9246 389036 241470
rect 388996 9240 389048 9246
rect 388996 9182 389048 9188
rect 389100 5778 389128 244052
rect 389744 242418 389772 244052
rect 389732 242412 389784 242418
rect 389732 242354 389784 242360
rect 390388 241670 390416 244052
rect 390376 241664 390428 241670
rect 390376 241606 390428 241612
rect 390940 241534 390968 244052
rect 391598 244038 391796 244066
rect 391204 242548 391256 242554
rect 391204 242490 391256 242496
rect 390928 241528 390980 241534
rect 390928 241470 390980 241476
rect 389088 5772 389140 5778
rect 389088 5714 389140 5720
rect 390652 4412 390704 4418
rect 390652 4354 390704 4360
rect 388628 4276 388680 4282
rect 388628 4218 388680 4224
rect 389456 3324 389508 3330
rect 389456 3266 389508 3272
rect 388536 3120 388588 3126
rect 388536 3062 388588 3068
rect 388444 3052 388496 3058
rect 388444 2994 388496 3000
rect 389468 480 389496 3266
rect 390664 480 390692 4354
rect 391216 3398 391244 242490
rect 391388 241936 391440 241942
rect 391388 241878 391440 241884
rect 391296 241732 391348 241738
rect 391296 241674 391348 241680
rect 391308 4593 391336 241674
rect 391294 4584 391350 4593
rect 391294 4519 391350 4528
rect 391400 4418 391428 241878
rect 391768 9178 391796 244038
rect 392228 242214 392256 244052
rect 392794 244038 393268 244066
rect 392216 242208 392268 242214
rect 392216 242150 392268 242156
rect 392584 241664 392636 241670
rect 392584 241606 392636 241612
rect 391848 241528 391900 241534
rect 391848 241470 391900 241476
rect 391756 9172 391808 9178
rect 391756 9114 391808 9120
rect 391860 5846 391888 241470
rect 391848 5840 391900 5846
rect 391848 5782 391900 5788
rect 391848 4480 391900 4486
rect 391848 4422 391900 4428
rect 391388 4412 391440 4418
rect 391388 4354 391440 4360
rect 391204 3392 391256 3398
rect 391204 3334 391256 3340
rect 391860 480 391888 4422
rect 392596 3330 392624 241606
rect 393240 5914 393268 244038
rect 393424 241942 393452 244052
rect 393412 241936 393464 241942
rect 393412 241878 393464 241884
rect 393976 241534 394004 244052
rect 394056 242004 394108 242010
rect 394056 241946 394108 241952
rect 393964 241528 394016 241534
rect 393778 241496 393834 241505
rect 394068 241505 394096 241946
rect 393964 241470 394016 241476
rect 394054 241496 394110 241505
rect 393778 241431 393834 241440
rect 394054 241431 394110 241440
rect 393792 231878 393820 241431
rect 393780 231872 393832 231878
rect 393780 231814 393832 231820
rect 393964 231872 394016 231878
rect 393964 231814 394016 231820
rect 393976 31754 394004 231814
rect 393964 31748 394016 31754
rect 393964 31690 394016 31696
rect 394148 31748 394200 31754
rect 394148 31690 394200 31696
rect 394160 28966 394188 31690
rect 394148 28960 394200 28966
rect 394148 28902 394200 28908
rect 394056 19372 394108 19378
rect 394056 19314 394108 19320
rect 394068 12458 394096 19314
rect 394068 12430 394464 12458
rect 393228 5908 393280 5914
rect 393228 5850 393280 5856
rect 394436 4622 394464 12430
rect 394620 5982 394648 244052
rect 395264 242418 395292 244052
rect 395344 242480 395396 242486
rect 395344 242422 395396 242428
rect 395252 242412 395304 242418
rect 395252 242354 395304 242360
rect 395356 8242 395384 242422
rect 395816 242010 395844 244052
rect 395804 242004 395856 242010
rect 395804 241946 395856 241952
rect 396460 241534 396488 244052
rect 397104 242486 397132 244052
rect 397656 242554 397684 244052
rect 398314 244038 398788 244066
rect 398104 242888 398156 242894
rect 398104 242830 398156 242836
rect 397644 242548 397696 242554
rect 397644 242490 397696 242496
rect 397092 242480 397144 242486
rect 397092 242422 397144 242428
rect 395436 241528 395488 241534
rect 395436 241470 395488 241476
rect 396448 241528 396500 241534
rect 396448 241470 396500 241476
rect 397368 241528 397420 241534
rect 397368 241470 397420 241476
rect 395264 8214 395384 8242
rect 394608 5976 394660 5982
rect 394608 5918 394660 5924
rect 394240 4616 394292 4622
rect 394240 4558 394292 4564
rect 394424 4616 394476 4622
rect 394424 4558 394476 4564
rect 394698 4584 394754 4593
rect 392584 3324 392636 3330
rect 392584 3266 392636 3272
rect 393044 3188 393096 3194
rect 393044 3130 393096 3136
rect 393056 480 393084 3130
rect 394252 480 394280 4558
rect 394698 4519 394754 4528
rect 394712 4486 394740 4519
rect 394700 4480 394752 4486
rect 394700 4422 394752 4428
rect 395264 4078 395292 8214
rect 395344 6452 395396 6458
rect 395344 6394 395396 6400
rect 395252 4072 395304 4078
rect 395252 4014 395304 4020
rect 395356 4026 395384 6394
rect 395448 4146 395476 241470
rect 397380 6050 397408 241470
rect 397368 6044 397420 6050
rect 397368 5986 397420 5992
rect 398116 4690 398144 242830
rect 398654 16824 398710 16833
rect 398654 16759 398656 16768
rect 398708 16759 398710 16768
rect 398656 16730 398708 16736
rect 398760 6866 398788 244038
rect 398944 241534 398972 244052
rect 399496 242894 399524 244052
rect 400048 244038 400154 244066
rect 399484 242888 399536 242894
rect 399484 242830 399536 242836
rect 398932 241528 398984 241534
rect 398932 241470 398984 241476
rect 400048 7070 400076 244038
rect 400784 241534 400812 244052
rect 401336 242622 401364 244052
rect 401324 242616 401376 242622
rect 401324 242558 401376 242564
rect 401980 241534 402008 244052
rect 402546 244038 402928 244066
rect 400128 241528 400180 241534
rect 400128 241470 400180 241476
rect 400772 241528 400824 241534
rect 400772 241470 400824 241476
rect 401508 241528 401560 241534
rect 401508 241470 401560 241476
rect 401968 241528 402020 241534
rect 401968 241470 402020 241476
rect 402796 241528 402848 241534
rect 402796 241470 402848 241476
rect 400036 7064 400088 7070
rect 400036 7006 400088 7012
rect 398748 6860 398800 6866
rect 398748 6802 398800 6808
rect 399024 6384 399076 6390
rect 399024 6326 399076 6332
rect 398748 5024 398800 5030
rect 398746 4992 398748 5001
rect 398800 4992 398802 5001
rect 398746 4927 398802 4936
rect 398840 4888 398892 4894
rect 398892 4836 398972 4842
rect 398840 4830 398972 4836
rect 398852 4814 398972 4830
rect 398944 4729 398972 4814
rect 398930 4720 398986 4729
rect 397828 4684 397880 4690
rect 397828 4626 397880 4632
rect 398104 4684 398156 4690
rect 398104 4626 398156 4632
rect 398840 4684 398892 4690
rect 398930 4655 398986 4664
rect 398840 4626 398892 4632
rect 395436 4140 395488 4146
rect 395436 4082 395488 4088
rect 395356 3998 395476 4026
rect 395448 480 395476 3998
rect 396632 3052 396684 3058
rect 396632 2994 396684 3000
rect 396644 480 396672 2994
rect 397840 480 397868 4626
rect 398852 4593 398880 4626
rect 398838 4584 398894 4593
rect 398838 4519 398894 4528
rect 399036 480 399064 6326
rect 400140 6118 400168 241470
rect 400862 16824 400918 16833
rect 400862 16759 400864 16768
rect 400916 16759 400918 16768
rect 400864 16730 400916 16736
rect 401520 6798 401548 241470
rect 402808 7138 402836 241470
rect 402796 7132 402848 7138
rect 402796 7074 402848 7080
rect 401508 6792 401560 6798
rect 401508 6734 401560 6740
rect 402900 6730 402928 244038
rect 403176 242690 403204 244052
rect 403834 244038 404308 244066
rect 403164 242684 403216 242690
rect 403164 242626 403216 242632
rect 403624 242548 403676 242554
rect 403624 242490 403676 242496
rect 403636 234734 403664 242490
rect 403624 234728 403676 234734
rect 403624 234670 403676 234676
rect 403532 234592 403584 234598
rect 403532 234534 403584 234540
rect 403544 231810 403572 234534
rect 403532 231804 403584 231810
rect 403532 231746 403584 231752
rect 403716 222216 403768 222222
rect 403716 222158 403768 222164
rect 403728 215218 403756 222158
rect 403532 215212 403584 215218
rect 403532 215154 403584 215160
rect 403716 215212 403768 215218
rect 403716 215154 403768 215160
rect 403544 205630 403572 215154
rect 403532 205624 403584 205630
rect 403532 205566 403584 205572
rect 403716 205624 403768 205630
rect 403716 205566 403768 205572
rect 403728 202881 403756 205566
rect 403714 202872 403770 202881
rect 403714 202807 403770 202816
rect 403990 202872 404046 202881
rect 403990 202807 404046 202816
rect 404004 193254 404032 202807
rect 403808 193248 403860 193254
rect 403808 193190 403860 193196
rect 403992 193248 404044 193254
rect 403992 193190 404044 193196
rect 403820 186266 403848 193190
rect 403728 186238 403848 186266
rect 403728 183569 403756 186238
rect 403714 183560 403770 183569
rect 403714 183495 403770 183504
rect 403990 183560 404046 183569
rect 403990 183495 404046 183504
rect 404004 173942 404032 183495
rect 403808 173936 403860 173942
rect 403808 173878 403860 173884
rect 403992 173936 404044 173942
rect 403992 173878 404044 173884
rect 403820 166954 403848 173878
rect 403728 166926 403848 166954
rect 403728 164218 403756 166926
rect 403532 164212 403584 164218
rect 403532 164154 403584 164160
rect 403716 164212 403768 164218
rect 403716 164154 403768 164160
rect 403544 154601 403572 164154
rect 403530 154592 403586 154601
rect 403530 154527 403586 154536
rect 403806 154592 403862 154601
rect 403806 154527 403862 154536
rect 403820 147642 403848 154527
rect 403636 147614 403848 147642
rect 403636 138106 403664 147614
rect 403624 138100 403676 138106
rect 403624 138042 403676 138048
rect 403532 137964 403584 137970
rect 403532 137906 403584 137912
rect 403544 135250 403572 137906
rect 403256 135244 403308 135250
rect 403256 135186 403308 135192
rect 403532 135244 403584 135250
rect 403532 135186 403584 135192
rect 403268 125633 403296 135186
rect 403254 125624 403310 125633
rect 403254 125559 403310 125568
rect 403438 125624 403494 125633
rect 403438 125559 403494 125568
rect 403452 118726 403480 125559
rect 403440 118720 403492 118726
rect 403440 118662 403492 118668
rect 403532 118652 403584 118658
rect 403532 118594 403584 118600
rect 403544 115938 403572 118594
rect 403256 115932 403308 115938
rect 403256 115874 403308 115880
rect 403532 115932 403584 115938
rect 403532 115874 403584 115880
rect 403268 106321 403296 115874
rect 403254 106312 403310 106321
rect 403254 106247 403310 106256
rect 403438 106312 403494 106321
rect 403438 106247 403494 106256
rect 403452 99414 403480 106247
rect 403440 99408 403492 99414
rect 403440 99350 403492 99356
rect 403532 99340 403584 99346
rect 403532 99282 403584 99288
rect 403544 96626 403572 99282
rect 403256 96620 403308 96626
rect 403256 96562 403308 96568
rect 403532 96620 403584 96626
rect 403532 96562 403584 96568
rect 403268 87009 403296 96562
rect 403254 87000 403310 87009
rect 403254 86935 403310 86944
rect 403438 87000 403494 87009
rect 403438 86935 403494 86944
rect 403452 80102 403480 86935
rect 403440 80096 403492 80102
rect 403440 80038 403492 80044
rect 403532 79960 403584 79966
rect 403532 79902 403584 79908
rect 403544 62150 403572 79902
rect 403440 62144 403492 62150
rect 403440 62086 403492 62092
rect 403532 62144 403584 62150
rect 403532 62086 403584 62092
rect 403452 60874 403480 62086
rect 403452 60846 403664 60874
rect 403636 52494 403664 60846
rect 403624 52488 403676 52494
rect 403624 52430 403676 52436
rect 403716 52488 403768 52494
rect 403716 52430 403768 52436
rect 403728 48346 403756 52430
rect 403716 48340 403768 48346
rect 403716 48282 403768 48288
rect 403808 48340 403860 48346
rect 403808 48282 403860 48288
rect 403820 48226 403848 48282
rect 403820 48198 403940 48226
rect 403912 38865 403940 48198
rect 403898 38856 403954 38865
rect 403898 38791 403954 38800
rect 403806 38720 403862 38729
rect 403806 38655 403862 38664
rect 403820 38622 403848 38655
rect 403808 38616 403860 38622
rect 403808 38558 403860 38564
rect 403900 29028 403952 29034
rect 403900 28970 403952 28976
rect 403912 22250 403940 28970
rect 403820 22222 403940 22250
rect 403820 19378 403848 22222
rect 403716 19372 403768 19378
rect 403716 19314 403768 19320
rect 403808 19372 403860 19378
rect 403808 19314 403860 19320
rect 403728 12458 403756 19314
rect 403728 12430 403848 12458
rect 402888 6724 402940 6730
rect 402888 6666 402940 6672
rect 400128 6112 400180 6118
rect 400128 6054 400180 6060
rect 403624 5092 403676 5098
rect 403624 5034 403676 5040
rect 403636 5001 403664 5034
rect 403622 4992 403678 5001
rect 403622 4927 403678 4936
rect 403716 4616 403768 4622
rect 401414 4584 401470 4593
rect 401324 4548 401376 4554
rect 403452 4564 403716 4570
rect 403452 4558 403768 4564
rect 403452 4554 403756 4558
rect 401414 4519 401416 4528
rect 401324 4490 401376 4496
rect 401468 4519 401470 4528
rect 403440 4548 403756 4554
rect 401416 4490 401468 4496
rect 403492 4542 403756 4548
rect 403440 4490 403492 4496
rect 400220 4004 400272 4010
rect 400220 3946 400272 3952
rect 400232 480 400260 3946
rect 401336 480 401364 4490
rect 402520 4276 402572 4282
rect 402520 4218 402572 4224
rect 402532 480 402560 4218
rect 403820 3398 403848 12430
rect 404280 7206 404308 244038
rect 404372 241534 404400 244052
rect 405016 242758 405044 244052
rect 405568 244038 405674 244066
rect 405004 242752 405056 242758
rect 405004 242694 405056 242700
rect 404360 241528 404412 241534
rect 404360 241470 404412 241476
rect 405568 7274 405596 244038
rect 406212 241534 406240 244052
rect 406856 242214 406884 244052
rect 406844 242208 406896 242214
rect 406844 242150 406896 242156
rect 407500 241534 407528 244052
rect 408066 244038 408448 244066
rect 405648 241528 405700 241534
rect 405648 241470 405700 241476
rect 406200 241528 406252 241534
rect 406200 241470 406252 241476
rect 407028 241528 407080 241534
rect 407028 241470 407080 241476
rect 407488 241528 407540 241534
rect 407488 241470 407540 241476
rect 408316 241528 408368 241534
rect 408316 241470 408368 241476
rect 405556 7268 405608 7274
rect 405556 7210 405608 7216
rect 404268 7200 404320 7206
rect 404268 7142 404320 7148
rect 405660 6662 405688 241470
rect 405648 6656 405700 6662
rect 405648 6598 405700 6604
rect 407040 6594 407068 241470
rect 408328 7342 408356 241470
rect 408316 7336 408368 7342
rect 408316 7278 408368 7284
rect 407028 6588 407080 6594
rect 407028 6530 407080 6536
rect 408420 6526 408448 244038
rect 408696 242146 408724 244052
rect 409354 244038 409828 244066
rect 409144 242344 409196 242350
rect 409144 242286 409196 242292
rect 408684 242140 408736 242146
rect 408684 242082 408736 242088
rect 408408 6520 408460 6526
rect 408408 6462 408460 6468
rect 406108 6316 406160 6322
rect 406108 6258 406160 6264
rect 404912 4820 404964 4826
rect 404912 4762 404964 4768
rect 405004 4820 405056 4826
rect 405004 4762 405056 4768
rect 403716 3392 403768 3398
rect 403716 3334 403768 3340
rect 403808 3392 403860 3398
rect 403808 3334 403860 3340
rect 403728 480 403756 3334
rect 404924 480 404952 4762
rect 405016 4729 405044 4762
rect 405002 4720 405058 4729
rect 405002 4655 405058 4664
rect 406120 480 406148 6258
rect 408500 5432 408552 5438
rect 408500 5374 408552 5380
rect 407304 3936 407356 3942
rect 407304 3878 407356 3884
rect 407316 480 407344 3878
rect 408512 480 408540 5374
rect 409156 3942 409184 242286
rect 409800 7410 409828 244038
rect 409892 241534 409920 244052
rect 410536 242350 410564 244052
rect 410524 242344 410576 242350
rect 410524 242286 410576 242292
rect 409880 241528 409932 241534
rect 409880 241470 409932 241476
rect 411088 7478 411116 244052
rect 411732 242282 411760 244052
rect 411260 242276 411312 242282
rect 411260 242218 411312 242224
rect 411720 242276 411772 242282
rect 411720 242218 411772 242224
rect 411272 241534 411300 242218
rect 412376 241534 412404 244052
rect 412548 242276 412600 242282
rect 412548 242218 412600 242224
rect 411168 241528 411220 241534
rect 411168 241470 411220 241476
rect 411260 241528 411312 241534
rect 411260 241470 411312 241476
rect 411904 241528 411956 241534
rect 411904 241470 411956 241476
rect 412364 241528 412416 241534
rect 412364 241470 412416 241476
rect 411076 7472 411128 7478
rect 411076 7414 411128 7420
rect 409788 7404 409840 7410
rect 409788 7346 409840 7352
rect 411180 6458 411208 241470
rect 411168 6452 411220 6458
rect 411168 6394 411220 6400
rect 409696 4344 409748 4350
rect 409696 4286 409748 4292
rect 409144 3936 409196 3942
rect 409144 3878 409196 3884
rect 409708 480 409736 4286
rect 410892 4072 410944 4078
rect 410892 4014 410944 4020
rect 410904 480 410932 4014
rect 411916 3058 411944 241470
rect 412560 6390 412588 242218
rect 412928 242146 412956 244052
rect 413586 244038 413876 244066
rect 414230 244038 414520 244066
rect 414782 244038 415348 244066
rect 412916 242140 412968 242146
rect 412916 242082 412968 242088
rect 412548 6384 412600 6390
rect 412548 6326 412600 6332
rect 413848 6322 413876 244038
rect 414492 242962 414520 244038
rect 414480 242956 414532 242962
rect 414480 242898 414532 242904
rect 413928 242140 413980 242146
rect 413928 242082 413980 242088
rect 413836 6316 413888 6322
rect 413836 6258 413888 6264
rect 413284 6248 413336 6254
rect 413284 6190 413336 6196
rect 412088 5500 412140 5506
rect 412088 5442 412140 5448
rect 411904 3052 411956 3058
rect 411904 2994 411956 3000
rect 412100 480 412128 5442
rect 413296 480 413324 6190
rect 413940 4282 413968 242082
rect 415320 4350 415348 244038
rect 415412 242146 415440 244052
rect 416056 242350 416084 244052
rect 416044 242344 416096 242350
rect 416044 242286 416096 242292
rect 415400 242140 415452 242146
rect 415400 242082 415452 242088
rect 416504 242140 416556 242146
rect 416504 242082 416556 242088
rect 416516 6254 416544 242082
rect 416504 6248 416556 6254
rect 416504 6190 416556 6196
rect 416608 5506 416636 244052
rect 416688 242344 416740 242350
rect 416688 242286 416740 242292
rect 416596 5500 416648 5506
rect 416596 5442 416648 5448
rect 415676 5364 415728 5370
rect 415676 5306 415728 5312
rect 415308 4344 415360 4350
rect 415308 4286 415360 4292
rect 413928 4276 413980 4282
rect 413928 4218 413980 4224
rect 414480 3868 414532 3874
rect 414480 3810 414532 3816
rect 414492 480 414520 3810
rect 415688 480 415716 5306
rect 416700 4010 416728 242286
rect 417252 242146 417280 244052
rect 417804 242185 417832 244052
rect 417790 242176 417846 242185
rect 417240 242140 417292 242146
rect 417790 242111 417846 242120
rect 418068 242140 418120 242146
rect 417240 242082 417292 242088
rect 418068 242082 418120 242088
rect 417974 16824 418030 16833
rect 417974 16759 417976 16768
rect 418028 16759 418030 16768
rect 417976 16730 418028 16736
rect 418080 6186 418108 242082
rect 418448 241534 418476 244052
rect 419106 244038 419396 244066
rect 418436 241528 418488 241534
rect 418436 241470 418488 241476
rect 418250 16824 418306 16833
rect 418250 16759 418252 16768
rect 418304 16759 418306 16768
rect 418252 16730 418304 16736
rect 419368 7546 419396 244038
rect 419644 242146 419672 244052
rect 420302 244038 420868 244066
rect 420184 242412 420236 242418
rect 420184 242354 420236 242360
rect 419632 242140 419684 242146
rect 419632 242082 419684 242088
rect 419448 241528 419500 241534
rect 419448 241470 419500 241476
rect 419356 7540 419408 7546
rect 419356 7482 419408 7488
rect 416872 6180 416924 6186
rect 416872 6122 416924 6128
rect 418068 6180 418120 6186
rect 418068 6122 418120 6128
rect 416688 4004 416740 4010
rect 416688 3946 416740 3952
rect 416884 480 416912 6122
rect 419460 5506 419488 241470
rect 419448 5500 419500 5506
rect 419448 5442 419500 5448
rect 419172 5296 419224 5302
rect 419172 5238 419224 5244
rect 420090 5264 420146 5273
rect 417976 3936 418028 3942
rect 417976 3878 418028 3884
rect 417988 480 418016 3878
rect 419184 480 419212 5238
rect 420090 5199 420146 5208
rect 420104 5098 420132 5199
rect 420092 5092 420144 5098
rect 420092 5034 420144 5040
rect 420196 2922 420224 242354
rect 420840 8158 420868 244038
rect 420932 241534 420960 244052
rect 421484 242418 421512 244052
rect 422142 244038 422248 244066
rect 421564 242480 421616 242486
rect 421564 242422 421616 242428
rect 421472 242412 421524 242418
rect 421472 242354 421524 242360
rect 420920 241528 420972 241534
rect 420920 241470 420972 241476
rect 420828 8152 420880 8158
rect 420828 8094 420880 8100
rect 421576 7698 421604 242422
rect 421656 242140 421708 242146
rect 421656 242082 421708 242088
rect 421484 7670 421604 7698
rect 420368 3800 420420 3806
rect 420368 3742 420420 3748
rect 420184 2916 420236 2922
rect 420184 2858 420236 2864
rect 420380 480 420408 3742
rect 421484 2990 421512 7670
rect 421668 3942 421696 242082
rect 422116 241528 422168 241534
rect 422116 241470 422168 241476
rect 422128 8294 422156 241470
rect 422116 8288 422168 8294
rect 422116 8230 422168 8236
rect 422220 4758 422248 244038
rect 422944 242276 422996 242282
rect 422944 242218 422996 242224
rect 422956 8242 422984 242218
rect 423232 241466 423260 244174
rect 423338 244038 423628 244066
rect 423220 241460 423272 241466
rect 423220 241402 423272 241408
rect 423312 239284 423364 239290
rect 423312 239226 423364 239232
rect 423324 231826 423352 239226
rect 423232 231798 423352 231826
rect 423232 225010 423260 231798
rect 423220 225004 423272 225010
rect 423220 224946 423272 224952
rect 423220 222216 423272 222222
rect 423220 222158 423272 222164
rect 423232 215422 423260 222158
rect 423220 215416 423272 215422
rect 423220 215358 423272 215364
rect 423220 215280 423272 215286
rect 423220 215222 423272 215228
rect 423232 205698 423260 215222
rect 423220 205692 423272 205698
rect 423220 205634 423272 205640
rect 423220 202904 423272 202910
rect 423220 202846 423272 202852
rect 423232 202774 423260 202846
rect 423220 202768 423272 202774
rect 423220 202710 423272 202716
rect 423312 193316 423364 193322
rect 423312 193258 423364 193264
rect 423324 193202 423352 193258
rect 423232 193174 423352 193202
rect 423232 186386 423260 193174
rect 423220 186380 423272 186386
rect 423220 186322 423272 186328
rect 423128 183592 423180 183598
rect 423128 183534 423180 183540
rect 423140 182170 423168 183534
rect 423128 182164 423180 182170
rect 423128 182106 423180 182112
rect 423220 182164 423272 182170
rect 423220 182106 423272 182112
rect 423232 173754 423260 182106
rect 423232 173726 423352 173754
rect 423324 172514 423352 173726
rect 423312 172508 423364 172514
rect 423312 172450 423364 172456
rect 423220 162920 423272 162926
rect 423220 162862 423272 162868
rect 423232 157418 423260 162862
rect 423220 157412 423272 157418
rect 423220 157354 423272 157360
rect 423312 157276 423364 157282
rect 423312 157218 423364 157224
rect 423324 153202 423352 157218
rect 423312 153196 423364 153202
rect 423312 153138 423364 153144
rect 423220 143608 423272 143614
rect 423220 143550 423272 143556
rect 423232 138038 423260 143550
rect 423220 138032 423272 138038
rect 423220 137974 423272 137980
rect 423312 137964 423364 137970
rect 423312 137906 423364 137912
rect 423324 129062 423352 137906
rect 423312 129056 423364 129062
rect 423312 128998 423364 129004
rect 423496 129056 423548 129062
rect 423496 128998 423548 129004
rect 423508 124273 423536 128998
rect 423310 124264 423366 124273
rect 423232 124222 423310 124250
rect 423232 122806 423260 124222
rect 423310 124199 423366 124208
rect 423494 124264 423550 124273
rect 423494 124199 423550 124208
rect 423220 122800 423272 122806
rect 423220 122742 423272 122748
rect 423312 113212 423364 113218
rect 423312 113154 423364 113160
rect 423324 109750 423352 113154
rect 423312 109744 423364 109750
rect 423312 109686 423364 109692
rect 423036 104916 423088 104922
rect 423036 104858 423088 104864
rect 423048 96626 423076 104858
rect 423036 96620 423088 96626
rect 423036 96562 423088 96568
rect 423128 96620 423180 96626
rect 423128 96562 423180 96568
rect 423140 86986 423168 96562
rect 423140 86970 423260 86986
rect 423140 86964 423272 86970
rect 423140 86958 423220 86964
rect 423220 86906 423272 86912
rect 423404 86964 423456 86970
rect 423404 86906 423456 86912
rect 423416 79914 423444 86906
rect 423324 79886 423444 79914
rect 423324 67658 423352 79886
rect 423220 67652 423272 67658
rect 423220 67594 423272 67600
rect 423312 67652 423364 67658
rect 423312 67594 423364 67600
rect 423232 58070 423260 67594
rect 423220 58064 423272 58070
rect 423220 58006 423272 58012
rect 423496 58064 423548 58070
rect 423496 58006 423548 58012
rect 423508 38758 423536 58006
rect 423312 38752 423364 38758
rect 423312 38694 423364 38700
rect 423496 38752 423548 38758
rect 423496 38694 423548 38700
rect 423324 31822 423352 38694
rect 423312 31816 423364 31822
rect 423312 31758 423364 31764
rect 423404 31680 423456 31686
rect 423404 31622 423456 31628
rect 423416 28914 423444 31622
rect 423416 28886 423536 28914
rect 423508 12458 423536 28886
rect 423416 12430 423536 12458
rect 422956 8214 423260 8242
rect 423416 8226 423444 12430
rect 422760 5228 422812 5234
rect 422760 5170 422812 5176
rect 422208 4752 422260 4758
rect 422208 4694 422260 4700
rect 421656 3936 421708 3942
rect 421656 3878 421708 3884
rect 421564 3732 421616 3738
rect 421564 3674 421616 3680
rect 421472 2984 421524 2990
rect 421472 2926 421524 2932
rect 421576 480 421604 3674
rect 422772 480 422800 5170
rect 423232 4078 423260 8214
rect 423404 8220 423456 8226
rect 423404 8162 423456 8168
rect 423220 4072 423272 4078
rect 423220 4014 423272 4020
rect 423600 3874 423628 244038
rect 423968 241534 423996 244052
rect 424626 244038 424916 244066
rect 423864 241528 423916 241534
rect 423864 241470 423916 241476
rect 423956 241528 424008 241534
rect 423956 241470 424008 241476
rect 424784 241528 424836 241534
rect 424784 241470 424836 241476
rect 423876 238626 423904 241470
rect 423876 238598 424364 238626
rect 424140 5432 424192 5438
rect 424140 5374 424192 5380
rect 424152 5273 424180 5374
rect 424138 5264 424194 5273
rect 424138 5199 424194 5208
rect 423956 4480 424008 4486
rect 423956 4422 424008 4428
rect 423588 3868 423640 3874
rect 423588 3810 423640 3816
rect 423968 480 423996 4422
rect 424336 3330 424364 238598
rect 424796 222290 424824 241470
rect 424692 222284 424744 222290
rect 424692 222226 424744 222232
rect 424784 222284 424836 222290
rect 424784 222226 424836 222232
rect 424704 222154 424732 222226
rect 424692 222148 424744 222154
rect 424692 222090 424744 222096
rect 424784 212560 424836 212566
rect 424598 212528 424654 212537
rect 424598 212463 424654 212472
rect 424782 212528 424784 212537
rect 424836 212528 424838 212537
rect 424782 212463 424838 212472
rect 424612 202910 424640 212463
rect 424600 202904 424652 202910
rect 424506 202872 424562 202881
rect 424692 202904 424744 202910
rect 424600 202846 424652 202852
rect 424690 202872 424692 202881
rect 424744 202872 424746 202881
rect 424506 202807 424562 202816
rect 424690 202807 424746 202816
rect 424520 193254 424548 202807
rect 424508 193248 424560 193254
rect 424784 193248 424836 193254
rect 424508 193190 424560 193196
rect 424598 193216 424654 193225
rect 424598 193151 424654 193160
rect 424782 193216 424784 193225
rect 424836 193216 424838 193225
rect 424782 193151 424838 193160
rect 424612 183598 424640 193151
rect 424600 183592 424652 183598
rect 424506 183560 424562 183569
rect 424692 183592 424744 183598
rect 424600 183534 424652 183540
rect 424690 183560 424692 183569
rect 424744 183560 424746 183569
rect 424506 183495 424562 183504
rect 424690 183495 424746 183504
rect 424520 182170 424548 183495
rect 424508 182164 424560 182170
rect 424508 182106 424560 182112
rect 424692 173868 424744 173874
rect 424692 173810 424744 173816
rect 424704 172514 424732 173810
rect 424692 172508 424744 172514
rect 424692 172450 424744 172456
rect 424782 162888 424838 162897
rect 424704 162858 424782 162874
rect 424692 162852 424782 162858
rect 424744 162846 424782 162852
rect 424782 162823 424838 162832
rect 424692 162794 424744 162800
rect 424692 157344 424744 157350
rect 424692 157286 424744 157292
rect 424704 153218 424732 157286
rect 424704 153202 424824 153218
rect 424692 153196 424836 153202
rect 424744 153190 424784 153196
rect 424692 153138 424744 153144
rect 424784 153138 424836 153144
rect 424704 143546 424732 153138
rect 424796 153107 424824 153138
rect 424692 143540 424744 143546
rect 424692 143482 424744 143488
rect 424692 137964 424744 137970
rect 424692 137906 424744 137912
rect 424704 133906 424732 137906
rect 424704 133890 424824 133906
rect 424704 133884 424836 133890
rect 424704 133878 424784 133884
rect 424784 133826 424836 133832
rect 424796 133795 424824 133826
rect 424692 124296 424744 124302
rect 424692 124238 424744 124244
rect 424704 124166 424732 124238
rect 424692 124160 424744 124166
rect 424692 124102 424744 124108
rect 424784 114572 424836 114578
rect 424784 114514 424836 114520
rect 424796 107098 424824 114514
rect 424784 107092 424836 107098
rect 424784 107034 424836 107040
rect 424692 99340 424744 99346
rect 424692 99282 424744 99288
rect 424704 96642 424732 99282
rect 424704 96614 424824 96642
rect 424796 86986 424824 96614
rect 424704 86970 424824 86986
rect 424692 86964 424824 86970
rect 424744 86958 424824 86964
rect 424692 86906 424744 86912
rect 424784 77308 424836 77314
rect 424784 77250 424836 77256
rect 424796 67833 424824 77250
rect 424782 67824 424838 67833
rect 424782 67759 424838 67768
rect 424690 67688 424746 67697
rect 424690 67623 424746 67632
rect 424704 67590 424732 67623
rect 424692 67584 424744 67590
rect 424692 67526 424744 67532
rect 424784 57996 424836 58002
rect 424784 57938 424836 57944
rect 424796 53122 424824 57938
rect 424704 53094 424824 53122
rect 424704 48278 424732 53094
rect 424692 48272 424744 48278
rect 424692 48214 424744 48220
rect 424784 38684 424836 38690
rect 424784 38626 424836 38632
rect 424796 31822 424824 38626
rect 424784 31816 424836 31822
rect 424784 31758 424836 31764
rect 424784 12504 424836 12510
rect 424784 12446 424836 12452
rect 424796 4690 424824 12446
rect 424888 8158 424916 244038
rect 425164 242622 425192 244052
rect 425152 242616 425204 242622
rect 425152 242558 425204 242564
rect 425808 241534 425836 244052
rect 426268 244038 426374 244066
rect 425796 241528 425848 241534
rect 425796 241470 425848 241476
rect 424968 172508 425020 172514
rect 424968 172450 425020 172456
rect 424980 162897 425008 172450
rect 424966 162888 425022 162897
rect 424966 162823 425022 162832
rect 424968 31816 425020 31822
rect 424968 31758 425020 31764
rect 424980 12510 425008 31758
rect 424968 12504 425020 12510
rect 424968 12446 425020 12452
rect 424876 8152 424928 8158
rect 424876 8094 424928 8100
rect 426268 8090 426296 244038
rect 427004 241534 427032 244052
rect 426348 241528 426400 241534
rect 426348 241470 426400 241476
rect 426992 241528 427044 241534
rect 426992 241470 427044 241476
rect 426256 8084 426308 8090
rect 426256 8026 426308 8032
rect 426360 5234 426388 241470
rect 427544 7676 427596 7682
rect 427544 7618 427596 7624
rect 426348 5228 426400 5234
rect 426348 5170 426400 5176
rect 424784 4684 424836 4690
rect 424784 4626 424836 4632
rect 426348 4548 426400 4554
rect 426348 4490 426400 4496
rect 424324 3324 424376 3330
rect 424324 3266 424376 3272
rect 425152 3052 425204 3058
rect 425152 2994 425204 3000
rect 425164 480 425192 2994
rect 426360 480 426388 4490
rect 427556 480 427584 7618
rect 427648 5166 427676 244052
rect 428200 241534 428228 244052
rect 428844 242282 428872 244052
rect 428832 242276 428884 242282
rect 428832 242218 428884 242224
rect 429488 241534 429516 244052
rect 430054 244038 430436 244066
rect 427728 241528 427780 241534
rect 427728 241470 427780 241476
rect 428188 241528 428240 241534
rect 428188 241470 428240 241476
rect 429108 241528 429160 241534
rect 429108 241470 429160 241476
rect 429476 241528 429528 241534
rect 429476 241470 429528 241476
rect 427636 5160 427688 5166
rect 427636 5102 427688 5108
rect 427636 4820 427688 4826
rect 427636 4762 427688 4768
rect 427648 4457 427676 4762
rect 427634 4448 427690 4457
rect 427634 4383 427690 4392
rect 427740 3806 427768 241470
rect 429120 8022 429148 241470
rect 429108 8016 429160 8022
rect 429108 7958 429160 7964
rect 430408 7954 430436 244038
rect 430684 241534 430712 244052
rect 431342 244038 431816 244066
rect 431224 242480 431276 242486
rect 431224 242422 431276 242428
rect 430488 241528 430540 241534
rect 430488 241470 430540 241476
rect 430672 241528 430724 241534
rect 430672 241470 430724 241476
rect 430396 7948 430448 7954
rect 430396 7890 430448 7896
rect 429936 5432 429988 5438
rect 429936 5374 429988 5380
rect 427910 4448 427966 4457
rect 427910 4383 427912 4392
rect 427964 4383 427966 4392
rect 427912 4354 427964 4360
rect 427728 3800 427780 3806
rect 427728 3742 427780 3748
rect 428740 3664 428792 3670
rect 428740 3606 428792 3612
rect 428752 480 428780 3606
rect 429948 480 429976 5374
rect 430500 5370 430528 241470
rect 430488 5364 430540 5370
rect 430488 5306 430540 5312
rect 431132 4820 431184 4826
rect 431132 4762 431184 4768
rect 431144 480 431172 4762
rect 431236 2854 431264 242422
rect 431684 241528 431736 241534
rect 431684 241470 431736 241476
rect 431696 7886 431724 241470
rect 431684 7880 431736 7886
rect 431684 7822 431736 7828
rect 431788 5438 431816 244038
rect 431880 241534 431908 244052
rect 432524 242622 432552 244052
rect 433182 244038 433288 244066
rect 432512 242616 432564 242622
rect 432512 242558 432564 242564
rect 431868 241528 431920 241534
rect 431868 241470 431920 241476
rect 431868 241392 431920 241398
rect 431868 241334 431920 241340
rect 431776 5432 431828 5438
rect 431776 5374 431828 5380
rect 431880 3738 431908 241334
rect 432604 5500 432656 5506
rect 432604 5442 432656 5448
rect 432616 5166 432644 5442
rect 432788 5432 432840 5438
rect 432788 5374 432840 5380
rect 432604 5160 432656 5166
rect 432604 5102 432656 5108
rect 432800 5098 432828 5374
rect 433260 5370 433288 244038
rect 433720 241534 433748 244052
rect 434378 244038 434668 244066
rect 433708 241528 433760 241534
rect 433708 241470 433760 241476
rect 434536 241528 434588 241534
rect 434536 241470 434588 241476
rect 434548 7818 434576 241470
rect 434536 7812 434588 7818
rect 434536 7754 434588 7760
rect 434536 7608 434588 7614
rect 434536 7550 434588 7556
rect 433248 5364 433300 5370
rect 433248 5306 433300 5312
rect 433524 5160 433576 5166
rect 433524 5102 433576 5108
rect 432788 5092 432840 5098
rect 432788 5034 432840 5040
rect 432696 5024 432748 5030
rect 432432 4972 432696 4978
rect 432432 4966 432748 4972
rect 432432 4950 432736 4966
rect 432432 4894 432460 4950
rect 432420 4888 432472 4894
rect 432420 4830 432472 4836
rect 431868 3732 431920 3738
rect 431868 3674 431920 3680
rect 432328 3596 432380 3602
rect 432328 3538 432380 3544
rect 431224 2848 431276 2854
rect 431224 2790 431276 2796
rect 432340 480 432368 3538
rect 433536 480 433564 5102
rect 434548 1714 434576 7550
rect 434640 3670 434668 244038
rect 434916 241534 434944 244052
rect 435574 244038 435956 244066
rect 435364 242752 435416 242758
rect 435364 242694 435416 242700
rect 434904 241528 434956 241534
rect 434904 241470 434956 241476
rect 434628 3664 434680 3670
rect 434628 3606 434680 3612
rect 435376 3058 435404 242694
rect 435928 7750 435956 244038
rect 436204 242758 436232 244052
rect 436192 242752 436244 242758
rect 436192 242694 436244 242700
rect 436756 241534 436784 244052
rect 437308 244038 437414 244066
rect 436008 241528 436060 241534
rect 436008 241470 436060 241476
rect 436744 241528 436796 241534
rect 436744 241470 436796 241476
rect 435916 7744 435968 7750
rect 435916 7686 435968 7692
rect 436020 5166 436048 241470
rect 437202 40216 437258 40225
rect 437202 40151 437258 40160
rect 437216 39817 437244 40151
rect 437202 39808 437258 39817
rect 437202 39743 437258 39752
rect 437202 16824 437258 16833
rect 437202 16759 437258 16768
rect 437216 16425 437244 16759
rect 437202 16416 437258 16425
rect 437202 16351 437258 16360
rect 437308 7682 437336 244038
rect 438044 241534 438072 244052
rect 438610 244038 438716 244066
rect 437388 241528 437440 241534
rect 437388 241470 437440 241476
rect 438032 241528 438084 241534
rect 438032 241470 438084 241476
rect 437296 7676 437348 7682
rect 437296 7618 437348 7624
rect 437400 5234 437428 241470
rect 437388 5228 437440 5234
rect 437388 5170 437440 5176
rect 436008 5160 436060 5166
rect 436008 5102 436060 5108
rect 438688 5030 438716 244038
rect 439044 242820 439096 242826
rect 439044 242762 439096 242768
rect 438768 241528 438820 241534
rect 438768 241470 438820 241476
rect 437020 5024 437072 5030
rect 437020 4966 437072 4972
rect 438676 5024 438728 5030
rect 438676 4966 438728 4972
rect 435824 3528 435876 3534
rect 435824 3470 435876 3476
rect 435364 3052 435416 3058
rect 435364 2994 435416 3000
rect 434548 1686 434668 1714
rect 434640 480 434668 1686
rect 435836 480 435864 3470
rect 437032 480 437060 4966
rect 438216 4888 438268 4894
rect 438216 4830 438268 4836
rect 438228 480 438256 4830
rect 438780 3602 438808 241470
rect 438768 3596 438820 3602
rect 438768 3538 438820 3544
rect 439056 610 439084 242762
rect 439240 241534 439268 244052
rect 439898 244038 440188 244066
rect 440160 241618 440188 244038
rect 440436 242146 440464 244052
rect 441094 244038 441476 244066
rect 440424 242140 440476 242146
rect 440424 242082 440476 242088
rect 440160 241590 440280 241618
rect 440252 241534 440280 241590
rect 439228 241528 439280 241534
rect 439228 241470 439280 241476
rect 440148 241528 440200 241534
rect 440148 241470 440200 241476
rect 440240 241528 440292 241534
rect 440240 241470 440292 241476
rect 440160 6225 440188 241470
rect 441448 7614 441476 244038
rect 441724 242146 441752 244052
rect 442290 244038 442856 244066
rect 441528 242140 441580 242146
rect 441528 242082 441580 242088
rect 441712 242140 441764 242146
rect 441712 242082 441764 242088
rect 441436 7608 441488 7614
rect 441436 7550 441488 7556
rect 440146 6216 440202 6225
rect 440146 6151 440202 6160
rect 441540 5166 441568 242082
rect 442724 242072 442776 242078
rect 442724 242014 442776 242020
rect 442736 7585 442764 242014
rect 442722 7576 442778 7585
rect 442722 7511 442778 7520
rect 441528 5160 441580 5166
rect 441528 5102 441580 5108
rect 440608 4956 440660 4962
rect 440608 4898 440660 4904
rect 439044 604 439096 610
rect 439044 546 439096 552
rect 439412 604 439464 610
rect 439412 546 439464 552
rect 439424 480 439452 546
rect 440620 480 440648 4898
rect 442828 4826 442856 244038
rect 442920 242078 442948 244052
rect 443472 242826 443500 244052
rect 444130 244038 444328 244066
rect 443460 242820 443512 242826
rect 443460 242762 443512 242768
rect 443000 242140 443052 242146
rect 443000 242082 443052 242088
rect 442908 242072 442960 242078
rect 442908 242014 442960 242020
rect 443012 241890 443040 242082
rect 442920 241862 443040 241890
rect 441804 4820 441856 4826
rect 441804 4762 441856 4768
rect 442816 4820 442868 4826
rect 442816 4762 442868 4768
rect 441816 480 441844 4762
rect 442920 3534 442948 241862
rect 444300 4894 444328 244038
rect 444760 242078 444788 244052
rect 445326 244038 445708 244066
rect 444748 242072 444800 242078
rect 444748 242014 444800 242020
rect 445576 242072 445628 242078
rect 445576 242014 445628 242020
rect 444380 40112 444432 40118
rect 444378 40080 444380 40089
rect 444432 40080 444434 40089
rect 444378 40015 444434 40024
rect 444380 16720 444432 16726
rect 444378 16688 444380 16697
rect 444432 16688 444434 16697
rect 444378 16623 444434 16632
rect 445588 9110 445616 242014
rect 445576 9104 445628 9110
rect 445576 9046 445628 9052
rect 445392 6996 445444 7002
rect 445392 6938 445444 6944
rect 444196 4888 444248 4894
rect 444196 4830 444248 4836
rect 444288 4888 444340 4894
rect 444288 4830 444340 4836
rect 442908 3528 442960 3534
rect 442908 3470 442960 3476
rect 443000 3460 443052 3466
rect 443000 3402 443052 3408
rect 443012 480 443040 3402
rect 444208 480 444236 4830
rect 445404 480 445432 6938
rect 445680 3466 445708 244038
rect 445760 242140 445812 242146
rect 445760 242082 445812 242088
rect 445668 3460 445720 3466
rect 445668 3402 445720 3408
rect 445772 610 445800 242082
rect 445956 242078 445984 244052
rect 446614 244038 446996 244066
rect 445944 242072 445996 242078
rect 445944 242014 445996 242020
rect 446968 9042 446996 244038
rect 447152 242146 447180 244052
rect 447140 242140 447192 242146
rect 447140 242082 447192 242088
rect 447796 242078 447824 244052
rect 448348 244038 448454 244066
rect 447048 242072 447100 242078
rect 447048 242014 447100 242020
rect 447784 242072 447836 242078
rect 447784 242014 447836 242020
rect 446956 9036 447008 9042
rect 446956 8978 447008 8984
rect 447060 4826 447088 242014
rect 447230 40352 447286 40361
rect 447230 40287 447286 40296
rect 447244 40118 447272 40287
rect 447232 40112 447284 40118
rect 447232 40054 447284 40060
rect 447230 16960 447286 16969
rect 447230 16895 447286 16904
rect 447244 16726 447272 16895
rect 447232 16720 447284 16726
rect 447232 16662 447284 16668
rect 448348 8974 448376 244038
rect 448992 242078 449020 244052
rect 448428 242072 448480 242078
rect 448428 242014 448480 242020
rect 448980 242072 449032 242078
rect 448980 242014 449032 242020
rect 448336 8968 448388 8974
rect 448336 8910 448388 8916
rect 448440 4865 448468 242014
rect 449176 182170 449204 545362
rect 449268 229090 449296 545430
rect 449360 405686 449388 549034
rect 449440 544808 449492 544814
rect 449440 544750 449492 544756
rect 449452 416770 449480 544750
rect 449544 452606 449572 549170
rect 449624 549160 449676 549166
rect 449624 549102 449676 549108
rect 449636 463690 449664 549102
rect 449716 544876 449768 544882
rect 449716 544818 449768 544824
rect 449728 487150 449756 544818
rect 449806 542872 449862 542881
rect 449806 542807 449862 542816
rect 449820 510610 449848 542807
rect 449808 510604 449860 510610
rect 449808 510546 449860 510552
rect 449716 487144 449768 487150
rect 449716 487086 449768 487092
rect 449624 463684 449676 463690
rect 449624 463626 449676 463632
rect 449532 452600 449584 452606
rect 449532 452542 449584 452548
rect 449440 416764 449492 416770
rect 449440 416706 449492 416712
rect 449348 405680 449400 405686
rect 449348 405622 449400 405628
rect 485780 242888 485832 242894
rect 485780 242830 485832 242836
rect 449808 242072 449860 242078
rect 449808 242014 449860 242020
rect 449256 229084 449308 229090
rect 449256 229026 449308 229032
rect 449164 182164 449216 182170
rect 449164 182106 449216 182112
rect 448980 9444 449032 9450
rect 448980 9386 449032 9392
rect 447782 4856 447838 4865
rect 447048 4820 447100 4826
rect 447782 4791 447838 4800
rect 448426 4856 448482 4865
rect 448426 4791 448482 4800
rect 447048 4762 447100 4768
rect 445760 604 445812 610
rect 445760 546 445812 552
rect 446588 604 446640 610
rect 446588 546 446640 552
rect 446600 480 446628 546
rect 447796 480 447824 4791
rect 448992 480 449020 9386
rect 449820 3369 449848 242014
rect 477592 242004 477644 242010
rect 477592 241946 477644 241952
rect 473360 241936 473412 241942
rect 473360 241878 473412 241884
rect 470600 241868 470652 241874
rect 470600 241810 470652 241816
rect 466460 241800 466512 241806
rect 466460 241742 466512 241748
rect 463700 241732 463752 241738
rect 463700 241674 463752 241680
rect 456800 241664 456852 241670
rect 456800 241606 456852 241612
rect 452660 241596 452712 241602
rect 452660 241538 452712 241544
rect 452476 9512 452528 9518
rect 452476 9454 452528 9460
rect 451280 4208 451332 4214
rect 451280 4150 451332 4156
rect 449806 3360 449862 3369
rect 449806 3295 449862 3304
rect 450176 3120 450228 3126
rect 450176 3062 450228 3068
rect 450188 480 450216 3062
rect 451292 480 451320 4150
rect 452488 480 452516 9454
rect 452672 3346 452700 241538
rect 456064 9376 456116 9382
rect 456064 9318 456116 9324
rect 454868 5568 454920 5574
rect 454868 5510 454920 5516
rect 452672 3318 453712 3346
rect 453684 480 453712 3318
rect 454880 480 454908 5510
rect 456076 480 456104 9318
rect 456812 3346 456840 241606
rect 459652 9308 459704 9314
rect 459652 9250 459704 9256
rect 458456 5636 458508 5642
rect 458456 5578 458508 5584
rect 456812 3318 457300 3346
rect 457272 480 457300 3318
rect 458468 480 458496 5578
rect 459664 480 459692 9250
rect 463240 9240 463292 9246
rect 463240 9182 463292 9188
rect 462044 5704 462096 5710
rect 462044 5646 462096 5652
rect 460848 3188 460900 3194
rect 460848 3130 460900 3136
rect 460860 480 460888 3130
rect 462056 480 462084 5646
rect 463252 480 463280 9182
rect 463712 3346 463740 241674
rect 465632 5772 465684 5778
rect 465632 5714 465684 5720
rect 463712 3318 464476 3346
rect 464448 480 464476 3318
rect 465644 480 465672 5714
rect 466472 3346 466500 241742
rect 470324 9172 470376 9178
rect 470324 9114 470376 9120
rect 469128 5840 469180 5846
rect 469128 5782 469180 5788
rect 466472 3318 466868 3346
rect 466840 480 466868 3318
rect 467932 3256 467984 3262
rect 467932 3198 467984 3204
rect 467944 480 467972 3198
rect 469140 480 469168 5782
rect 470336 480 470364 9114
rect 470612 610 470640 241810
rect 471886 40488 471942 40497
rect 471886 40423 471942 40432
rect 471900 40089 471928 40423
rect 471886 40080 471942 40089
rect 471886 40015 471942 40024
rect 471886 17096 471942 17105
rect 471886 17031 471942 17040
rect 471900 16697 471928 17031
rect 471886 16688 471942 16697
rect 471886 16623 471942 16632
rect 472716 5908 472768 5914
rect 472716 5850 472768 5856
rect 470600 604 470652 610
rect 470600 546 470652 552
rect 471520 604 471572 610
rect 471520 546 471572 552
rect 471532 480 471560 546
rect 472728 480 472756 5850
rect 473372 610 473400 241878
rect 476028 40112 476080 40118
rect 476026 40080 476028 40089
rect 476080 40080 476082 40089
rect 476026 40015 476082 40024
rect 476028 16720 476080 16726
rect 476026 16688 476028 16697
rect 476080 16688 476082 16697
rect 476026 16623 476082 16632
rect 476304 5976 476356 5982
rect 476304 5918 476356 5924
rect 475108 4140 475160 4146
rect 475108 4082 475160 4088
rect 473360 604 473412 610
rect 473360 546 473412 552
rect 473912 604 473964 610
rect 473912 546 473964 552
rect 473924 480 473952 546
rect 475120 480 475148 4082
rect 476316 480 476344 5918
rect 477500 2916 477552 2922
rect 477500 2858 477552 2864
rect 477512 480 477540 2858
rect 477604 610 477632 241946
rect 482926 40352 482982 40361
rect 482926 40287 482982 40296
rect 482940 40118 482968 40287
rect 482928 40112 482980 40118
rect 482928 40054 482980 40060
rect 482926 16960 482982 16969
rect 482926 16895 482982 16904
rect 482940 16726 482968 16895
rect 482928 16720 482980 16726
rect 482928 16662 482980 16668
rect 483480 6860 483532 6866
rect 483480 6802 483532 6808
rect 479892 6044 479944 6050
rect 479892 5986 479944 5992
rect 477592 604 477644 610
rect 477592 546 477644 552
rect 478696 604 478748 610
rect 478696 546 478748 552
rect 478708 480 478736 546
rect 479904 480 479932 5986
rect 482284 3392 482336 3398
rect 482284 3334 482336 3340
rect 481088 2984 481140 2990
rect 481088 2926 481140 2932
rect 481100 480 481128 2926
rect 482296 480 482324 3334
rect 483492 480 483520 6802
rect 484584 6112 484636 6118
rect 484584 6054 484636 6060
rect 484596 480 484624 6054
rect 485792 480 485820 242830
rect 525064 242752 525116 242758
rect 525064 242694 525116 242700
rect 492680 242684 492732 242690
rect 492680 242626 492732 242632
rect 490564 7132 490616 7138
rect 490564 7074 490616 7080
rect 486976 7064 487028 7070
rect 486976 7006 487028 7012
rect 486988 480 487016 7006
rect 488172 6792 488224 6798
rect 488172 6734 488224 6740
rect 488184 480 488212 6734
rect 489368 2848 489420 2854
rect 489368 2790 489420 2796
rect 489380 480 489408 2790
rect 490576 480 490604 7074
rect 491760 6724 491812 6730
rect 491760 6666 491812 6672
rect 491772 480 491800 6666
rect 492692 626 492720 242626
rect 523684 242616 523736 242622
rect 523684 242558 523736 242564
rect 502984 242548 503036 242554
rect 502984 242490 503036 242496
rect 499580 242208 499632 242214
rect 499580 242150 499632 242156
rect 497740 7268 497792 7274
rect 497740 7210 497792 7216
rect 494152 7200 494204 7206
rect 494152 7142 494204 7148
rect 492692 598 492904 626
rect 492876 592 492904 598
rect 492876 564 492996 592
rect 492968 480 492996 564
rect 494164 480 494192 7142
rect 495348 6656 495400 6662
rect 495348 6598 495400 6604
rect 495360 480 495388 6598
rect 496544 3052 496596 3058
rect 496544 2994 496596 3000
rect 496556 480 496584 2994
rect 497752 480 497780 7210
rect 498936 6588 498988 6594
rect 498936 6530 498988 6536
rect 498948 480 498976 6530
rect 499592 610 499620 242150
rect 501236 7336 501288 7342
rect 501236 7278 501288 7284
rect 499580 604 499632 610
rect 499580 546 499632 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500144 480 500172 546
rect 501248 480 501276 7278
rect 502432 6520 502484 6526
rect 502432 6462 502484 6468
rect 502444 480 502472 6462
rect 502996 3058 503024 242490
rect 518164 242480 518216 242486
rect 518164 242422 518216 242428
rect 514024 242412 514076 242418
rect 514024 242354 514076 242360
rect 507124 242344 507176 242350
rect 507124 242286 507176 242292
rect 504824 7404 504876 7410
rect 504824 7346 504876 7352
rect 503628 3324 503680 3330
rect 503628 3266 503680 3272
rect 502984 3052 503036 3058
rect 502984 2994 503036 3000
rect 503640 480 503668 3266
rect 504836 480 504864 7346
rect 506020 6452 506072 6458
rect 506020 6394 506072 6400
rect 506032 480 506060 6394
rect 507136 4146 507164 242286
rect 511262 242176 511318 242185
rect 511262 242111 511318 242120
rect 508412 7472 508464 7478
rect 508412 7414 508464 7420
rect 507124 4140 507176 4146
rect 507124 4082 507176 4088
rect 507216 3052 507268 3058
rect 507216 2994 507268 3000
rect 507228 480 507256 2994
rect 508424 480 508452 7414
rect 509608 6384 509660 6390
rect 509608 6326 509660 6332
rect 509620 480 509648 6326
rect 511276 4078 511304 242111
rect 513196 6316 513248 6322
rect 513196 6258 513248 6264
rect 512000 4276 512052 4282
rect 512000 4218 512052 4224
rect 510804 4072 510856 4078
rect 510804 4014 510856 4020
rect 511264 4072 511316 4078
rect 511264 4014 511316 4020
rect 510816 480 510844 4014
rect 512012 480 512040 4218
rect 513208 480 513236 6258
rect 514036 3194 514064 242354
rect 516784 6248 516836 6254
rect 516784 6190 516836 6196
rect 515588 4344 515640 4350
rect 515588 4286 515640 4292
rect 514392 4140 514444 4146
rect 514392 4082 514444 4088
rect 514024 3188 514076 3194
rect 514024 3130 514076 3136
rect 514404 480 514432 4082
rect 515600 480 515628 4286
rect 516796 480 516824 6190
rect 517888 4004 517940 4010
rect 517888 3946 517940 3952
rect 517900 480 517928 3946
rect 518176 3262 518204 242422
rect 520924 242276 520976 242282
rect 520924 242218 520976 242224
rect 520280 6180 520332 6186
rect 520280 6122 520332 6128
rect 519084 4480 519136 4486
rect 519084 4422 519136 4428
rect 518164 3256 518216 3262
rect 518164 3198 518216 3204
rect 519096 480 519124 4422
rect 520292 480 520320 6122
rect 520936 3330 520964 242218
rect 522672 4412 522724 4418
rect 522672 4354 522724 4360
rect 521476 4072 521528 4078
rect 521476 4014 521528 4020
rect 520924 3324 520976 3330
rect 520924 3266 520976 3272
rect 521488 480 521516 4014
rect 522684 480 522712 4354
rect 523696 3398 523724 242558
rect 523868 7540 523920 7546
rect 523868 7482 523920 7488
rect 523684 3392 523736 3398
rect 523684 3334 523736 3340
rect 523880 480 523908 7482
rect 525076 4146 525104 242694
rect 529204 242140 529256 242146
rect 529204 242082 529256 242088
rect 527824 241528 527876 241534
rect 527824 241470 527876 241476
rect 527456 8288 527508 8294
rect 527456 8230 527508 8236
rect 526260 4548 526312 4554
rect 526260 4490 526312 4496
rect 525064 4140 525116 4146
rect 525064 4082 525116 4088
rect 525064 3936 525116 3942
rect 525064 3878 525116 3884
rect 525076 480 525104 3878
rect 526272 480 526300 4490
rect 527468 480 527496 8230
rect 527836 4078 527864 241470
rect 527824 4072 527876 4078
rect 527824 4014 527876 4020
rect 529216 4010 529244 242082
rect 530584 242072 530636 242078
rect 530584 242014 530636 242020
rect 529848 4616 529900 4622
rect 529848 4558 529900 4564
rect 529204 4004 529256 4010
rect 529204 3946 529256 3952
rect 528652 3188 528704 3194
rect 528652 3130 528704 3136
rect 528664 480 528692 3130
rect 529860 480 529888 4558
rect 530596 3942 530624 242014
rect 577516 30326 577544 552026
rect 577778 548448 577834 548457
rect 577778 548383 577834 548392
rect 577594 548176 577650 548185
rect 577594 548111 577650 548120
rect 577608 64734 577636 548111
rect 577688 543992 577740 543998
rect 577688 543934 577740 543940
rect 577700 77246 577728 543934
rect 577792 111790 577820 548383
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545358 580212 545527
rect 580172 545352 580224 545358
rect 580172 545294 580224 545300
rect 580724 545216 580776 545222
rect 580724 545158 580776 545164
rect 580540 545148 580592 545154
rect 580540 545090 580592 545096
rect 580080 544740 580132 544746
rect 580080 544682 580132 544688
rect 578056 544468 578108 544474
rect 578056 544410 578108 544416
rect 577964 544332 578016 544338
rect 577964 544274 578016 544280
rect 577872 544128 577924 544134
rect 577872 544070 577924 544076
rect 577884 135250 577912 544070
rect 577976 158710 578004 544274
rect 578068 205630 578096 544410
rect 579618 543688 579674 543697
rect 579618 543623 579674 543632
rect 579632 439929 579660 543623
rect 579802 543552 579858 543561
rect 579802 543487 579858 543496
rect 579618 439920 579674 439929
rect 579618 439855 579674 439864
rect 579816 393009 579844 543487
rect 579986 543416 580042 543425
rect 579986 543351 580042 543360
rect 579896 534064 579948 534070
rect 579896 534006 579948 534012
rect 579908 533905 579936 534006
rect 579894 533896 579950 533905
rect 579894 533831 579950 533840
rect 579896 510604 579948 510610
rect 579896 510546 579948 510552
rect 579908 510377 579936 510546
rect 579894 510368 579950 510377
rect 579894 510303 579950 510312
rect 579802 393000 579858 393009
rect 579802 392935 579858 392944
rect 580000 369617 580028 543351
rect 580092 498681 580120 544682
rect 580448 544400 580500 544406
rect 580448 544342 580500 544348
rect 580356 544196 580408 544202
rect 580356 544138 580408 544144
rect 580170 543280 580226 543289
rect 580170 543215 580226 543224
rect 580078 498672 580134 498681
rect 580078 498607 580134 498616
rect 580080 487144 580132 487150
rect 580080 487086 580132 487092
rect 580092 486849 580120 487086
rect 580078 486840 580134 486849
rect 580078 486775 580134 486784
rect 580080 463684 580132 463690
rect 580080 463626 580132 463632
rect 580092 463457 580120 463626
rect 580078 463448 580134 463457
rect 580078 463383 580134 463392
rect 580080 452600 580132 452606
rect 580080 452542 580132 452548
rect 580092 451761 580120 452542
rect 580078 451752 580134 451761
rect 580078 451687 580134 451696
rect 580080 416764 580132 416770
rect 580080 416706 580132 416712
rect 580092 416537 580120 416706
rect 580078 416528 580134 416537
rect 580078 416463 580134 416472
rect 580080 405680 580132 405686
rect 580080 405622 580132 405628
rect 580092 404841 580120 405622
rect 580078 404832 580134 404841
rect 580078 404767 580134 404776
rect 579986 369608 580042 369617
rect 579986 369543 580042 369552
rect 580184 346089 580212 543215
rect 580264 542904 580316 542910
rect 580264 542846 580316 542852
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 578056 205624 578108 205630
rect 578056 205566 578108 205572
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 577964 158704 578016 158710
rect 577964 158646 578016 158652
rect 580080 158704 580132 158710
rect 580080 158646 580132 158652
rect 580092 158409 580120 158646
rect 580078 158400 580134 158409
rect 580078 158335 580134 158344
rect 577872 135244 577924 135250
rect 577872 135186 577924 135192
rect 577780 111784 577832 111790
rect 577780 111726 577832 111732
rect 580276 87961 580304 542846
rect 580368 123185 580396 544138
rect 580460 170105 580488 544342
rect 580552 217025 580580 545090
rect 580632 544536 580684 544542
rect 580632 544478 580684 544484
rect 580644 263945 580672 544478
rect 580736 275777 580764 545158
rect 580908 544604 580960 544610
rect 580908 544546 580960 544552
rect 580814 543144 580870 543153
rect 580814 543079 580870 543088
rect 580828 310865 580856 543079
rect 580920 322697 580948 544546
rect 580906 322688 580962 322697
rect 580906 322623 580962 322632
rect 580814 310856 580870 310865
rect 580814 310791 580870 310800
rect 580722 275768 580778 275777
rect 580722 275703 580778 275712
rect 580630 263936 580686 263945
rect 580630 263871 580686 263880
rect 580538 217016 580594 217025
rect 580538 216951 580594 216960
rect 580816 205624 580868 205630
rect 580816 205566 580868 205572
rect 580828 205329 580856 205566
rect 580814 205320 580870 205329
rect 580814 205255 580870 205264
rect 580446 170096 580502 170105
rect 580446 170031 580502 170040
rect 580632 135244 580684 135250
rect 580632 135186 580684 135192
rect 580644 134881 580672 135186
rect 580630 134872 580686 134881
rect 580630 134807 580686 134816
rect 580354 123176 580410 123185
rect 580354 123111 580410 123120
rect 580632 111784 580684 111790
rect 580632 111726 580684 111732
rect 580644 111489 580672 111726
rect 580630 111480 580686 111489
rect 580630 111415 580686 111424
rect 580262 87952 580318 87961
rect 580262 87887 580318 87896
rect 577688 77240 577740 77246
rect 577688 77182 577740 77188
rect 579620 77240 579672 77246
rect 579620 77182 579672 77188
rect 579632 76265 579660 77182
rect 579618 76256 579674 76265
rect 579618 76191 579674 76200
rect 577596 64728 577648 64734
rect 577596 64670 577648 64676
rect 580356 64728 580408 64734
rect 580356 64670 580408 64676
rect 580368 64569 580396 64670
rect 580354 64560 580410 64569
rect 580354 64495 580410 64504
rect 577504 30320 577556 30326
rect 577504 30262 577556 30268
rect 579620 30320 579672 30326
rect 579620 30262 579672 30268
rect 579632 29345 579660 30262
rect 579618 29336 579674 29345
rect 579618 29271 579674 29280
rect 573824 9104 573876 9110
rect 573824 9046 573876 9052
rect 531044 8220 531096 8226
rect 531044 8162 531096 8168
rect 530584 3936 530636 3942
rect 530584 3878 530636 3884
rect 531056 480 531084 8162
rect 534540 8152 534592 8158
rect 534540 8094 534592 8100
rect 533436 4684 533488 4690
rect 533436 4626 533488 4632
rect 532240 3868 532292 3874
rect 532240 3810 532292 3816
rect 532252 480 532280 3810
rect 533448 480 533476 4626
rect 534552 480 534580 8094
rect 538128 8084 538180 8090
rect 538128 8026 538180 8032
rect 536932 4752 536984 4758
rect 536932 4694 536984 4700
rect 535736 3256 535788 3262
rect 535736 3198 535788 3204
rect 535748 480 535776 3198
rect 536944 480 536972 4694
rect 538140 480 538168 8026
rect 541716 8016 541768 8022
rect 541716 7958 541768 7964
rect 540520 5500 540572 5506
rect 540520 5442 540572 5448
rect 539324 3800 539376 3806
rect 539324 3742 539376 3748
rect 539336 480 539364 3742
rect 540532 480 540560 5442
rect 541728 480 541756 7958
rect 545304 7948 545356 7954
rect 545304 7890 545356 7896
rect 544108 5432 544160 5438
rect 544108 5374 544160 5380
rect 542912 3324 542964 3330
rect 542912 3266 542964 3272
rect 542924 480 542952 3266
rect 544120 480 544148 5374
rect 545316 480 545344 7890
rect 548892 7880 548944 7886
rect 548892 7822 548944 7828
rect 547696 5364 547748 5370
rect 547696 5306 547748 5312
rect 546500 3732 546552 3738
rect 546500 3674 546552 3680
rect 546512 480 546540 3674
rect 547708 480 547736 5306
rect 548904 480 548932 7822
rect 552388 7812 552440 7818
rect 552388 7754 552440 7760
rect 551192 5296 551244 5302
rect 551192 5238 551244 5244
rect 550088 3392 550140 3398
rect 550088 3334 550140 3340
rect 550100 480 550128 3334
rect 551204 480 551232 5238
rect 552400 480 552428 7754
rect 555976 7744 556028 7750
rect 555976 7686 556028 7692
rect 554780 5228 554832 5234
rect 554780 5170 554832 5176
rect 553584 3664 553636 3670
rect 553584 3606 553636 3612
rect 553596 480 553624 3606
rect 554792 480 554820 5170
rect 555988 480 556016 7686
rect 559564 7676 559616 7682
rect 559564 7618 559616 7624
rect 558368 5160 558420 5166
rect 558368 5102 558420 5108
rect 557172 4140 557224 4146
rect 557172 4082 557224 4088
rect 557184 480 557212 4082
rect 558380 480 558408 5102
rect 559576 480 559604 7618
rect 566740 7608 566792 7614
rect 566740 7550 566792 7556
rect 570234 7576 570290 7585
rect 563150 6216 563206 6225
rect 563150 6151 563206 6160
rect 561956 5024 562008 5030
rect 561956 4966 562008 4972
rect 560760 3596 560812 3602
rect 560760 3538 560812 3544
rect 560772 480 560800 3538
rect 561968 480 561996 4966
rect 563164 480 563192 6151
rect 565544 5092 565596 5098
rect 565544 5034 565596 5040
rect 564348 4072 564400 4078
rect 564348 4014 564400 4020
rect 564360 480 564388 4014
rect 565556 480 565584 5034
rect 566752 480 566780 7550
rect 570234 7511 570290 7520
rect 569040 4956 569092 4962
rect 569040 4898 569092 4904
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 567856 480 567884 3470
rect 569052 480 569080 4898
rect 570248 480 570276 7511
rect 572628 4888 572680 4894
rect 572628 4830 572680 4836
rect 571432 4004 571484 4010
rect 571432 3946 571484 3952
rect 571444 480 571472 3946
rect 572640 480 572668 4830
rect 573836 480 573864 9046
rect 577412 9036 577464 9042
rect 577412 8978 577464 8984
rect 576216 4820 576268 4826
rect 576216 4762 576268 4768
rect 575020 3460 575072 3466
rect 575020 3402 575072 3408
rect 575032 480 575060 3402
rect 576228 480 576256 4762
rect 577424 480 577452 8978
rect 581000 8968 581052 8974
rect 581000 8910 581052 8916
rect 579802 4856 579858 4865
rect 579802 4791 579858 4800
rect 578608 3936 578660 3942
rect 578608 3878 578660 3884
rect 578620 480 578648 3878
rect 579816 480 579844 4791
rect 581012 480 581040 8910
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 582208 480 582236 3295
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 3422 567296 3478 567352
rect 3422 553016 3478 553072
rect 4802 549208 4858 549264
rect 2962 538600 3018 538656
rect 2962 509940 2964 509960
rect 2964 509940 3016 509960
rect 3016 509940 3018 509960
rect 2962 509904 3018 509940
rect 2778 495524 2780 495544
rect 2780 495524 2832 495544
rect 2832 495524 2834 495544
rect 2778 495488 2834 495524
rect 2778 481108 2780 481128
rect 2780 481108 2832 481128
rect 2832 481108 2834 481128
rect 2778 481072 2834 481108
rect 3054 452376 3110 452432
rect 2778 437960 2834 438016
rect 2778 423680 2834 423736
rect 3146 394984 3202 395040
rect 2962 380604 2964 380624
rect 2964 380604 3016 380624
rect 3016 380604 3018 380624
rect 2962 380568 3018 380604
rect 2778 366152 2834 366208
rect 3698 547984 3754 548040
rect 3330 542952 3386 543008
rect 3238 337456 3294 337512
rect 3146 323040 3202 323096
rect 3330 308760 3386 308816
rect 3146 280100 3148 280120
rect 3148 280100 3200 280120
rect 3200 280100 3202 280120
rect 3146 280064 3202 280100
rect 2778 265648 2834 265704
rect 3054 236952 3110 237008
rect 3330 222536 3386 222592
rect 2778 193876 2780 193896
rect 2780 193876 2832 193896
rect 2832 193876 2834 193896
rect 2778 193840 2834 193876
rect 2778 179460 2780 179480
rect 2780 179460 2832 179480
rect 2832 179460 2834 179480
rect 2778 179424 2834 179460
rect 3330 150728 3386 150784
rect 2962 122712 3018 122768
rect 2962 122032 3018 122088
rect 3330 80008 3386 80064
rect 3330 78920 3386 78976
rect 3330 64504 3386 64560
rect 4066 294344 4122 294400
rect 3974 251232 4030 251288
rect 3882 136312 3938 136368
rect 3790 107616 3846 107672
rect 3698 93200 3754 93256
rect 3606 50088 3662 50144
rect 3514 35808 3570 35864
rect 3422 21392 3478 21448
rect 21362 548256 21418 548312
rect 13082 242120 13138 242176
rect 2778 7112 2834 7168
rect 5262 3304 5318 3360
rect 12438 4800 12494 4856
rect 210698 549072 210754 549128
rect 197818 548936 197874 548992
rect 189998 548664 190054 548720
rect 166722 548392 166778 548448
rect 158994 548120 159050 548176
rect 299570 560496 299626 560552
rect 299570 560360 299626 560416
rect 331310 700304 331366 700360
rect 365074 686024 365130 686080
rect 364522 685888 364578 685944
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 364154 579672 364210 579728
rect 364338 579672 364394 579728
rect 493874 579672 493930 579728
rect 494058 579672 494114 579728
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 440882 549208 440938 549264
rect 407302 548800 407358 548856
rect 415030 548528 415086 548584
rect 435730 548256 435786 548312
rect 425334 547984 425390 548040
rect 27894 8880 27950 8936
rect 37370 6160 37426 6216
rect 70674 7520 70730 7576
rect 44546 6296 44602 6352
rect 93858 5364 93914 5400
rect 93858 5344 93860 5364
rect 93860 5344 93912 5364
rect 93912 5344 93914 5364
rect 103426 5364 103482 5400
rect 103426 5344 103428 5364
rect 103428 5344 103480 5364
rect 103480 5344 103482 5364
rect 113178 5364 113234 5400
rect 113178 5344 113180 5364
rect 113180 5344 113232 5364
rect 113232 5344 113234 5364
rect 122654 5364 122710 5400
rect 122654 5344 122656 5364
rect 122656 5344 122708 5364
rect 122708 5344 122710 5364
rect 132498 5364 132554 5400
rect 132498 5344 132500 5364
rect 132500 5344 132552 5364
rect 132552 5344 132554 5364
rect 141974 5364 142030 5400
rect 141974 5344 141976 5364
rect 141976 5344 142028 5364
rect 142028 5344 142030 5364
rect 142158 4972 142160 4992
rect 142160 4972 142212 4992
rect 142212 4972 142214 4992
rect 142158 4936 142214 4972
rect 422482 545264 422538 545320
rect 430486 545128 430542 545184
rect 151542 544584 151598 544640
rect 154026 544584 154082 544640
rect 203154 544584 203210 544640
rect 205454 544584 205510 544640
rect 208030 544584 208086 544640
rect 213458 544584 213514 544640
rect 221278 544584 221334 544640
rect 231582 544584 231638 544640
rect 386510 544584 386566 544640
rect 151726 237088 151782 237144
rect 151726 221040 151782 221096
rect 151634 206216 151690 206272
rect 151634 193160 151690 193216
rect 151818 193160 151874 193216
rect 151450 177248 151506 177304
rect 151450 165416 151506 165472
rect 150714 164328 150770 164384
rect 150806 164192 150862 164248
rect 151542 112920 151598 112976
rect 151542 104216 151598 104272
rect 151082 92792 151138 92848
rect 150990 92656 151046 92712
rect 150714 92520 150770 92576
rect 151082 91296 151138 91352
rect 151358 81368 151414 81424
rect 151358 71848 151414 71904
rect 150530 51040 150586 51096
rect 150714 51040 150770 51096
rect 150530 33088 150586 33144
rect 150714 33088 150770 33144
rect 153290 242120 153346 242176
rect 152002 201320 152058 201376
rect 152002 196560 152058 196616
rect 152738 215192 152794 215248
rect 152738 208256 152794 208312
rect 152002 193160 152058 193216
rect 152094 15136 152150 15192
rect 152278 15136 152334 15192
rect 152002 5616 152058 5672
rect 152278 5616 152334 5672
rect 150898 4956 150954 4992
rect 150898 4936 150900 4956
rect 150900 4936 150952 4956
rect 150952 4936 150954 4956
rect 152002 3304 152058 3360
rect 153382 220768 153438 220824
rect 153566 220768 153622 220824
rect 153382 133884 153438 133920
rect 153382 133864 153384 133884
rect 153384 133864 153436 133884
rect 153436 133864 153438 133884
rect 153566 133864 153622 133920
rect 154762 183504 154818 183560
rect 154946 183504 155002 183560
rect 154854 173848 154910 173904
rect 155038 173848 155094 173904
rect 154854 164192 154910 164248
rect 155038 164192 155094 164248
rect 154762 86944 154818 87000
rect 154946 86944 155002 87000
rect 156142 133884 156198 133920
rect 156142 133864 156144 133884
rect 156144 133864 156196 133884
rect 156196 133864 156198 133884
rect 156326 133864 156382 133920
rect 155958 4800 156014 4856
rect 162858 87080 162914 87136
rect 162950 86944 163006 87000
rect 164422 8880 164478 8936
rect 168562 202816 168618 202872
rect 168838 202816 168894 202872
rect 169758 202816 169814 202872
rect 169942 202816 169998 202872
rect 168562 183504 168618 183560
rect 168838 183504 168894 183560
rect 169758 183504 169814 183560
rect 169942 183504 169998 183560
rect 168470 143520 168526 143576
rect 168838 143520 168894 143576
rect 169758 135224 169814 135280
rect 170034 135224 170090 135280
rect 169758 115912 169814 115968
rect 170034 115912 170090 115968
rect 169758 96600 169814 96656
rect 170034 96600 170090 96656
rect 168654 67768 168710 67824
rect 168562 67598 168618 67654
rect 168470 6160 168526 6216
rect 173990 183504 174046 183560
rect 174266 183504 174322 183560
rect 173898 16668 173900 16688
rect 173900 16668 173952 16688
rect 173952 16668 173954 16688
rect 173898 16632 173954 16668
rect 172610 6296 172666 6352
rect 176382 40296 176438 40352
rect 176566 40296 176622 40352
rect 177946 57976 178002 58032
rect 179694 241440 179750 241496
rect 179878 241440 179934 241496
rect 179602 231820 179604 231840
rect 179604 231820 179656 231840
rect 179656 231820 179658 231840
rect 179602 231784 179658 231820
rect 179786 231784 179842 231840
rect 178222 202816 178278 202872
rect 178406 202816 178462 202872
rect 178222 183504 178278 183560
rect 178406 183504 178462 183560
rect 178222 154536 178278 154592
rect 178406 154536 178462 154592
rect 178222 135224 178278 135280
rect 178406 135224 178462 135280
rect 178130 57976 178186 58032
rect 178682 5344 178738 5400
rect 183466 16668 183468 16688
rect 183468 16668 183520 16688
rect 183520 16668 183522 16688
rect 183466 16632 183522 16668
rect 183466 5344 183522 5400
rect 185214 241440 185270 241496
rect 185398 241440 185454 241496
rect 185122 231820 185124 231840
rect 185124 231820 185176 231840
rect 185176 231820 185178 231840
rect 185122 231784 185178 231820
rect 185306 231784 185362 231840
rect 185030 7520 185086 7576
rect 188986 95240 189042 95296
rect 190458 212472 190514 212528
rect 190458 202852 190460 202872
rect 190460 202852 190512 202872
rect 190512 202852 190514 202872
rect 190458 202816 190514 202852
rect 190458 153176 190514 153232
rect 189262 145016 189318 145072
rect 189262 144880 189318 144936
rect 190366 133864 190422 133920
rect 189262 125704 189318 125760
rect 189262 125568 189318 125624
rect 190458 124208 190514 124264
rect 189170 104760 189226 104816
rect 189170 85448 189226 85504
rect 189262 85312 189318 85368
rect 189262 27784 189318 27840
rect 189170 27648 189226 27704
rect 190734 222128 190790 222184
rect 190918 222128 190974 222184
rect 190734 212508 190736 212528
rect 190736 212508 190788 212528
rect 190788 212508 190790 212528
rect 190734 212472 190790 212508
rect 190642 202852 190644 202872
rect 190644 202852 190696 202872
rect 190696 202852 190698 202872
rect 190642 202816 190698 202852
rect 190734 193196 190736 193216
rect 190736 193196 190788 193216
rect 190788 193196 190790 193216
rect 190734 193160 190790 193196
rect 190918 193160 190974 193216
rect 190734 153176 190790 153232
rect 190642 133884 190698 133920
rect 190642 133864 190644 133884
rect 190644 133864 190696 133884
rect 190696 133864 190698 133884
rect 190642 124208 190698 124264
rect 190642 106276 190698 106312
rect 190642 106256 190644 106276
rect 190644 106256 190696 106276
rect 190696 106256 190698 106276
rect 190826 106256 190882 106312
rect 190642 86964 190698 87000
rect 190642 86944 190644 86964
rect 190644 86944 190696 86964
rect 190696 86944 190698 86964
rect 190826 86944 190882 87000
rect 191746 222128 191802 222184
rect 191930 222164 191932 222184
rect 191932 222164 191984 222184
rect 191984 222164 191986 222184
rect 191930 222128 191986 222164
rect 192022 202952 192078 203008
rect 191838 202816 191894 202872
rect 192022 193196 192024 193216
rect 192024 193196 192076 193216
rect 192076 193196 192078 193216
rect 192022 193160 192078 193196
rect 192206 193160 192262 193216
rect 192022 162832 192078 162888
rect 192114 162696 192170 162752
rect 191930 144900 191986 144936
rect 191930 144880 191932 144900
rect 191932 144880 191984 144900
rect 191984 144880 191986 144900
rect 192114 144880 192170 144936
rect 191838 135224 191894 135280
rect 192022 135224 192078 135280
rect 191746 111696 191802 111752
rect 191930 111696 191986 111752
rect 191930 44104 191986 44160
rect 192114 44104 192170 44160
rect 191746 26152 191802 26208
rect 191930 26152 191986 26208
rect 194506 198736 194562 198792
rect 194506 44104 194562 44160
rect 195978 198736 196034 198792
rect 194782 198464 194838 198520
rect 194782 44104 194838 44160
rect 196346 198464 196402 198520
rect 196162 140664 196218 140720
rect 196254 140528 196310 140584
rect 198186 211132 198242 211168
rect 198186 211112 198188 211132
rect 198188 211112 198240 211132
rect 198240 211112 198242 211132
rect 198370 211132 198426 211168
rect 198370 211112 198372 211132
rect 198372 211112 198424 211132
rect 198424 211112 198426 211132
rect 201498 40180 201554 40216
rect 201498 40160 201500 40180
rect 201500 40160 201552 40180
rect 201552 40160 201554 40180
rect 206926 220768 206982 220824
rect 207110 220768 207166 220824
rect 206926 211112 206982 211168
rect 207110 211112 207166 211168
rect 205914 201476 205970 201512
rect 205914 201456 205916 201476
rect 205916 201456 205968 201476
rect 205968 201456 205970 201476
rect 206098 201456 206154 201512
rect 207018 135224 207074 135280
rect 207202 135224 207258 135280
rect 207110 116048 207166 116104
rect 207018 115912 207074 115968
rect 208398 191800 208454 191856
rect 208582 191800 208638 191856
rect 208582 85584 208638 85640
rect 208766 85584 208822 85640
rect 213826 242120 213882 242176
rect 216586 183504 216642 183560
rect 216770 183504 216826 183560
rect 216862 162968 216918 163024
rect 216770 162832 216826 162888
rect 217966 151816 218022 151872
rect 217966 151680 218022 151736
rect 218426 229064 218482 229120
rect 218978 229064 219034 229120
rect 218334 162968 218390 163024
rect 218242 162832 218298 162888
rect 219346 40024 219402 40080
rect 219530 230424 219586 230480
rect 219714 230424 219770 230480
rect 219530 211132 219586 211168
rect 219530 211112 219532 211132
rect 219532 211112 219584 211132
rect 219584 211112 219586 211132
rect 219714 211112 219770 211168
rect 222474 135224 222530 135280
rect 222658 135224 222714 135280
rect 223762 231784 223818 231840
rect 223946 231784 224002 231840
rect 223762 211112 223818 211168
rect 223946 211112 224002 211168
rect 223854 182144 223910 182200
rect 224038 182144 224094 182200
rect 223762 135224 223818 135280
rect 223946 135224 224002 135280
rect 224038 87080 224094 87136
rect 223854 86964 223910 87000
rect 223854 86944 223856 86964
rect 223856 86944 223908 86964
rect 223908 86944 223910 86964
rect 225050 231820 225052 231840
rect 225052 231820 225104 231840
rect 225104 231820 225106 231840
rect 225050 231784 225106 231820
rect 225234 231784 225290 231840
rect 225142 220804 225144 220824
rect 225144 220804 225196 220824
rect 225196 220804 225198 220824
rect 225142 220768 225198 220804
rect 225326 220768 225382 220824
rect 226706 190576 226762 190632
rect 226430 190460 226486 190496
rect 226430 190440 226432 190460
rect 226432 190440 226484 190460
rect 226484 190440 226486 190460
rect 226614 180784 226670 180840
rect 226798 180784 226854 180840
rect 226522 154672 226578 154728
rect 226522 154556 226578 154592
rect 226522 154536 226524 154556
rect 226524 154536 226576 154556
rect 226576 154536 226578 154556
rect 226522 135224 226578 135280
rect 226706 135224 226762 135280
rect 229006 40296 229062 40352
rect 229006 39752 229062 39808
rect 229282 135224 229338 135280
rect 229466 135224 229522 135280
rect 231214 3612 231216 3632
rect 231216 3612 231268 3632
rect 231268 3612 231270 3632
rect 231214 3576 231270 3612
rect 232502 3576 232558 3632
rect 234802 193196 234804 193216
rect 234804 193196 234856 193216
rect 234856 193196 234858 193216
rect 234802 193160 234858 193196
rect 234986 193160 235042 193216
rect 234802 162832 234858 162888
rect 234986 162832 235042 162888
rect 234802 135244 234858 135280
rect 234802 135224 234804 135244
rect 234804 135224 234856 135244
rect 234856 135224 234858 135244
rect 234986 135244 235042 135280
rect 234986 135224 234988 135244
rect 234988 135224 235040 135244
rect 235040 135224 235042 135244
rect 234802 87080 234858 87136
rect 234710 86944 234766 87000
rect 236366 116048 236422 116104
rect 236274 115932 236330 115968
rect 236274 115912 236276 115932
rect 236276 115912 236328 115932
rect 236328 115912 236330 115932
rect 238482 240080 238538 240136
rect 238666 240080 238722 240136
rect 238482 220768 238538 220824
rect 238666 220768 238722 220824
rect 238482 211112 238538 211168
rect 238666 211112 238722 211168
rect 238482 201476 238538 201512
rect 238482 201456 238484 201476
rect 238484 201456 238536 201476
rect 238536 201456 238538 201476
rect 238666 201476 238722 201512
rect 238666 201456 238668 201476
rect 238668 201456 238720 201476
rect 238720 201456 238722 201476
rect 238390 153176 238446 153232
rect 238574 153176 238630 153232
rect 237654 116048 237710 116104
rect 237562 115932 237618 115968
rect 237562 115912 237564 115932
rect 237564 115912 237616 115932
rect 237616 115912 237618 115932
rect 237562 87080 237618 87136
rect 237470 86944 237526 87000
rect 238666 40568 238722 40624
rect 238666 40024 238722 40080
rect 239034 193196 239036 193216
rect 239036 193196 239088 193216
rect 239088 193196 239090 193216
rect 239034 193160 239090 193196
rect 239218 193196 239220 193216
rect 239220 193196 239272 193216
rect 239272 193196 239274 193216
rect 239218 193160 239274 193196
rect 240046 40568 240102 40624
rect 240046 40296 240102 40352
rect 247958 230424 248014 230480
rect 248142 230460 248144 230480
rect 248144 230460 248196 230480
rect 248196 230460 248198 230480
rect 248142 230424 248198 230460
rect 245842 202816 245898 202872
rect 246118 202816 246174 202872
rect 247038 202816 247094 202872
rect 247222 202816 247278 202872
rect 245842 183504 245898 183560
rect 246118 183504 246174 183560
rect 247038 183504 247094 183560
rect 247222 183504 247278 183560
rect 248142 172488 248198 172544
rect 248326 172488 248382 172544
rect 247038 154536 247094 154592
rect 247314 154536 247370 154592
rect 245750 114688 245806 114744
rect 245934 114552 245990 114608
rect 245750 95376 245806 95432
rect 245934 95240 245990 95296
rect 252558 183504 252614 183560
rect 252742 183504 252798 183560
rect 258078 202816 258134 202872
rect 258262 202816 258318 202872
rect 258078 183504 258134 183560
rect 258262 183504 258318 183560
rect 258078 154536 258134 154592
rect 258354 154536 258410 154592
rect 258078 135224 258134 135280
rect 258354 135224 258410 135280
rect 258078 115912 258134 115968
rect 258354 115912 258410 115968
rect 258078 96600 258134 96656
rect 258354 96600 258410 96656
rect 259550 242120 259606 242176
rect 265162 231784 265218 231840
rect 265346 231784 265402 231840
rect 263598 202816 263654 202872
rect 263782 202816 263838 202872
rect 263598 183504 263654 183560
rect 263782 183504 263838 183560
rect 265070 144880 265126 144936
rect 265254 144880 265310 144936
rect 263782 143656 263838 143712
rect 263782 143520 263838 143576
rect 265070 135224 265126 135280
rect 265254 135224 265310 135280
rect 263782 67768 263838 67824
rect 263782 67632 263838 67688
rect 263690 48184 263746 48240
rect 263782 48048 263838 48104
rect 268474 241576 268530 241632
rect 270590 241576 270646 241632
rect 270498 231784 270554 231840
rect 270682 231784 270738 231840
rect 270498 144880 270554 144936
rect 270774 144880 270830 144936
rect 271878 202816 271934 202872
rect 272062 202816 272118 202872
rect 271878 183504 271934 183560
rect 272062 183504 272118 183560
rect 271878 144880 271934 144936
rect 272062 144880 272118 144936
rect 271878 125568 271934 125624
rect 272062 125568 272118 125624
rect 284390 183504 284446 183560
rect 284666 183504 284722 183560
rect 302146 40160 302202 40216
rect 302330 40160 302386 40216
rect 302146 16768 302202 16824
rect 302330 16768 302386 16824
rect 303618 96620 303674 96656
rect 303618 96600 303620 96620
rect 303620 96600 303672 96620
rect 303672 96600 303674 96620
rect 303986 96600 304042 96656
rect 307666 57976 307722 58032
rect 307942 183504 307998 183560
rect 308218 183504 308274 183560
rect 307850 57976 307906 58032
rect 307942 48184 307998 48240
rect 308034 38664 308090 38720
rect 318798 16788 318854 16824
rect 318798 16768 318800 16788
rect 318800 16768 318852 16788
rect 318852 16768 318854 16788
rect 321282 40180 321338 40216
rect 321282 40160 321284 40180
rect 321284 40160 321336 40180
rect 321336 40160 321338 40180
rect 321558 40180 321614 40216
rect 321558 40160 321560 40180
rect 321560 40160 321612 40180
rect 321612 40160 321614 40180
rect 321558 16788 321614 16824
rect 321558 16768 321560 16788
rect 321560 16768 321612 16788
rect 321612 16768 321614 16788
rect 338210 16804 338212 16824
rect 338212 16804 338264 16824
rect 338264 16804 338266 16824
rect 338210 16768 338266 16804
rect 340694 40196 340696 40216
rect 340696 40196 340748 40216
rect 340748 40196 340750 40216
rect 340694 40160 340750 40196
rect 340970 40196 340972 40216
rect 340972 40196 341024 40216
rect 341024 40196 341026 40216
rect 340970 40160 341026 40196
rect 342626 16804 342628 16824
rect 342628 16804 342680 16824
rect 342680 16804 342682 16824
rect 342626 16768 342682 16804
rect 346030 183504 346086 183560
rect 346214 183504 346270 183560
rect 346122 77152 346178 77208
rect 346306 77152 346362 77208
rect 353666 242120 353722 242176
rect 357530 242256 357586 242312
rect 357070 183504 357126 183560
rect 357254 183504 357310 183560
rect 359922 40180 359978 40216
rect 359922 40160 359924 40180
rect 359924 40160 359976 40180
rect 359976 40160 359978 40180
rect 359922 16804 359924 16824
rect 359924 16804 359976 16824
rect 359976 16804 359978 16824
rect 359922 16768 359978 16804
rect 360198 40180 360254 40216
rect 360198 40160 360200 40180
rect 360200 40160 360252 40180
rect 360252 40160 360254 40180
rect 362222 16804 362224 16824
rect 362224 16804 362276 16824
rect 362276 16804 362278 16824
rect 362222 16768 362278 16804
rect 367098 242684 367154 242720
rect 367098 242664 367100 242684
rect 367100 242664 367152 242684
rect 367152 242664 367154 242684
rect 367098 242548 367154 242584
rect 367098 242528 367100 242548
rect 367100 242528 367152 242548
rect 367152 242528 367154 242548
rect 367190 242392 367246 242448
rect 367006 242256 367062 242312
rect 367466 242548 367522 242584
rect 367466 242528 367468 242548
rect 367468 242528 367520 242548
rect 367520 242528 367522 242548
rect 369582 242412 369638 242448
rect 369582 242392 369584 242412
rect 369584 242392 369636 242412
rect 369636 242392 369638 242412
rect 367650 241712 367706 241768
rect 374274 242664 374330 242720
rect 374274 241474 374330 241530
rect 374274 240080 374330 240136
rect 374458 240080 374514 240136
rect 374274 220768 374330 220824
rect 374458 220768 374514 220824
rect 374274 211112 374330 211168
rect 374458 211112 374514 211168
rect 374274 191800 374330 191856
rect 374458 191800 374514 191856
rect 374274 172488 374330 172544
rect 374458 172488 374514 172544
rect 378874 230696 378930 230752
rect 379242 230424 379298 230480
rect 379058 201456 379114 201512
rect 379242 201456 379298 201512
rect 379150 37168 379206 37224
rect 379334 37168 379390 37224
rect 379242 16804 379244 16824
rect 379244 16804 379296 16824
rect 379296 16804 379298 16824
rect 379242 16768 379298 16804
rect 379334 4972 379336 4992
rect 379336 4972 379388 4992
rect 379388 4972 379390 4992
rect 379334 4936 379390 4972
rect 379610 16804 379612 16824
rect 379612 16804 379664 16824
rect 379664 16804 379666 16824
rect 379610 16768 379666 16804
rect 379518 4972 379520 4992
rect 379520 4972 379572 4992
rect 379572 4972 379574 4992
rect 379518 4936 379574 4972
rect 380806 4800 380862 4856
rect 384670 230424 384726 230480
rect 384854 230424 384910 230480
rect 384670 135224 384726 135280
rect 384854 135224 384910 135280
rect 384670 96620 384726 96656
rect 384670 96600 384672 96620
rect 384672 96600 384724 96620
rect 384724 96600 384726 96620
rect 384854 96620 384910 96656
rect 384854 96600 384856 96620
rect 384856 96600 384908 96620
rect 384908 96600 384910 96620
rect 384670 86944 384726 87000
rect 384854 86944 384910 87000
rect 388442 242120 388498 242176
rect 391294 4528 391350 4584
rect 393778 241440 393834 241496
rect 394054 241440 394110 241496
rect 394698 4528 394754 4584
rect 398654 16788 398710 16824
rect 398654 16768 398656 16788
rect 398656 16768 398708 16788
rect 398708 16768 398710 16788
rect 398746 4972 398748 4992
rect 398748 4972 398800 4992
rect 398800 4972 398802 4992
rect 398746 4936 398802 4972
rect 398930 4664 398986 4720
rect 398838 4528 398894 4584
rect 400862 16788 400918 16824
rect 400862 16768 400864 16788
rect 400864 16768 400916 16788
rect 400916 16768 400918 16788
rect 403714 202816 403770 202872
rect 403990 202816 404046 202872
rect 403714 183504 403770 183560
rect 403990 183504 404046 183560
rect 403530 154536 403586 154592
rect 403806 154536 403862 154592
rect 403254 125568 403310 125624
rect 403438 125568 403494 125624
rect 403254 106256 403310 106312
rect 403438 106256 403494 106312
rect 403254 86944 403310 87000
rect 403438 86944 403494 87000
rect 403898 38800 403954 38856
rect 403806 38664 403862 38720
rect 403622 4936 403678 4992
rect 401414 4548 401470 4584
rect 401414 4528 401416 4548
rect 401416 4528 401468 4548
rect 401468 4528 401470 4548
rect 405002 4664 405058 4720
rect 417790 242120 417846 242176
rect 417974 16788 418030 16824
rect 417974 16768 417976 16788
rect 417976 16768 418028 16788
rect 418028 16768 418030 16788
rect 418250 16788 418306 16824
rect 418250 16768 418252 16788
rect 418252 16768 418304 16788
rect 418304 16768 418306 16788
rect 420090 5208 420146 5264
rect 423310 124208 423366 124264
rect 423494 124208 423550 124264
rect 424138 5208 424194 5264
rect 424598 212472 424654 212528
rect 424782 212508 424784 212528
rect 424784 212508 424836 212528
rect 424836 212508 424838 212528
rect 424782 212472 424838 212508
rect 424506 202816 424562 202872
rect 424690 202852 424692 202872
rect 424692 202852 424744 202872
rect 424744 202852 424746 202872
rect 424690 202816 424746 202852
rect 424598 193160 424654 193216
rect 424782 193196 424784 193216
rect 424784 193196 424836 193216
rect 424836 193196 424838 193216
rect 424782 193160 424838 193196
rect 424506 183504 424562 183560
rect 424690 183540 424692 183560
rect 424692 183540 424744 183560
rect 424744 183540 424746 183560
rect 424690 183504 424746 183540
rect 424782 162832 424838 162888
rect 424782 67768 424838 67824
rect 424690 67632 424746 67688
rect 424966 162832 425022 162888
rect 427634 4392 427690 4448
rect 427910 4412 427966 4448
rect 427910 4392 427912 4412
rect 427912 4392 427964 4412
rect 427964 4392 427966 4412
rect 437202 40160 437258 40216
rect 437202 39752 437258 39808
rect 437202 16768 437258 16824
rect 437202 16360 437258 16416
rect 440146 6160 440202 6216
rect 442722 7520 442778 7576
rect 444378 40060 444380 40080
rect 444380 40060 444432 40080
rect 444432 40060 444434 40080
rect 444378 40024 444434 40060
rect 444378 16668 444380 16688
rect 444380 16668 444432 16688
rect 444432 16668 444434 16688
rect 444378 16632 444434 16668
rect 447230 40296 447286 40352
rect 447230 16904 447286 16960
rect 449806 542816 449862 542872
rect 447782 4800 447838 4856
rect 448426 4800 448482 4856
rect 449806 3304 449862 3360
rect 471886 40432 471942 40488
rect 471886 40024 471942 40080
rect 471886 17040 471942 17096
rect 471886 16632 471942 16688
rect 476026 40060 476028 40080
rect 476028 40060 476080 40080
rect 476080 40060 476082 40080
rect 476026 40024 476082 40060
rect 476026 16668 476028 16688
rect 476028 16668 476080 16688
rect 476080 16668 476082 16688
rect 476026 16632 476082 16668
rect 482926 40296 482982 40352
rect 482926 16904 482982 16960
rect 511262 242120 511318 242176
rect 577778 548392 577834 548448
rect 577594 548120 577650 548176
rect 580170 545536 580226 545592
rect 579618 543632 579674 543688
rect 579802 543496 579858 543552
rect 579618 439864 579674 439920
rect 579986 543360 580042 543416
rect 579894 533840 579950 533896
rect 579894 510312 579950 510368
rect 579802 392944 579858 393000
rect 580170 543224 580226 543280
rect 580078 498616 580134 498672
rect 580078 486784 580134 486840
rect 580078 463392 580134 463448
rect 580078 451696 580134 451752
rect 580078 416472 580134 416528
rect 580078 404776 580134 404832
rect 579986 369552 580042 369608
rect 580170 346024 580226 346080
rect 580170 228792 580226 228848
rect 580170 181872 580226 181928
rect 580078 158344 580134 158400
rect 580814 543088 580870 543144
rect 580906 322632 580962 322688
rect 580814 310800 580870 310856
rect 580722 275712 580778 275768
rect 580630 263880 580686 263936
rect 580538 216960 580594 217016
rect 580814 205264 580870 205320
rect 580446 170040 580502 170096
rect 580630 134816 580686 134872
rect 580354 123120 580410 123176
rect 580630 111424 580686 111480
rect 580262 87896 580318 87952
rect 579618 76200 579674 76256
rect 580354 64504 580410 64560
rect 579618 29280 579674 29336
rect 563150 6160 563206 6216
rect 570234 7520 570290 7576
rect 579802 4800 579858 4856
rect 582194 3304 582250 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 331305 700362 331371 700365
rect 8109 700360 331371 700362
rect 8109 700304 8114 700360
rect 8170 700304 331310 700360
rect 331366 700304 331371 700360
rect 8109 700302 331371 700304
rect 8109 700299 8175 700302
rect 331305 700299 331371 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 365069 686082 365135 686085
rect 494881 686082 494947 686085
rect 364382 686080 365135 686082
rect 364382 686024 365074 686080
rect 365130 686024 365135 686080
rect 364382 686022 365135 686024
rect 364382 685946 364442 686022
rect 365069 686019 365135 686022
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 364517 685946 364583 685949
rect 364382 685944 364583 685946
rect 364382 685888 364522 685944
rect 364578 685888 364583 685944
rect 364382 685886 364583 685888
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 364517 685883 364583 685886
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 364149 579730 364215 579733
rect 364333 579730 364399 579733
rect 364149 579728 364399 579730
rect 364149 579672 364154 579728
rect 364210 579672 364338 579728
rect 364394 579672 364399 579728
rect 364149 579670 364399 579672
rect 364149 579667 364215 579670
rect 364333 579667 364399 579670
rect 493869 579730 493935 579733
rect 494053 579730 494119 579733
rect 493869 579728 494119 579730
rect 493869 579672 493874 579728
rect 493930 579672 494058 579728
rect 494114 579672 494119 579728
rect 493869 579670 494119 579672
rect 493869 579667 493935 579670
rect 494053 579667 494119 579670
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 299565 560554 299631 560557
rect 299430 560552 299631 560554
rect 299430 560496 299570 560552
rect 299626 560496 299631 560552
rect 299430 560494 299631 560496
rect 299430 560418 299490 560494
rect 299565 560491 299631 560494
rect 299565 560418 299631 560421
rect 299430 560416 299631 560418
rect 299430 560360 299570 560416
rect 299626 560360 299631 560416
rect 299430 560358 299631 560360
rect 299565 560355 299631 560358
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3417 553074 3483 553077
rect -960 553072 3483 553074
rect -960 553016 3422 553072
rect 3478 553016 3483 553072
rect -960 553014 3483 553016
rect -960 552924 480 553014
rect 3417 553011 3483 553014
rect 4797 549266 4863 549269
rect 440877 549266 440943 549269
rect 4797 549264 440943 549266
rect 4797 549208 4802 549264
rect 4858 549208 440882 549264
rect 440938 549208 440943 549264
rect 4797 549206 440943 549208
rect 4797 549203 4863 549206
rect 440877 549203 440943 549206
rect 210693 549130 210759 549133
rect 447726 549130 447732 549132
rect 210693 549128 447732 549130
rect 210693 549072 210698 549128
rect 210754 549072 447732 549128
rect 210693 549070 447732 549072
rect 210693 549067 210759 549070
rect 447726 549068 447732 549070
rect 447796 549068 447802 549132
rect 197813 548994 197879 548997
rect 446622 548994 446628 548996
rect 197813 548992 446628 548994
rect 197813 548936 197818 548992
rect 197874 548936 446628 548992
rect 197813 548934 446628 548936
rect 197813 548931 197879 548934
rect 446622 548932 446628 548934
rect 446692 548932 446698 548996
rect 152774 548796 152780 548860
rect 152844 548858 152850 548860
rect 407297 548858 407363 548861
rect 152844 548856 407363 548858
rect 152844 548800 407302 548856
rect 407358 548800 407363 548856
rect 152844 548798 407363 548800
rect 152844 548796 152850 548798
rect 407297 548795 407363 548798
rect 189993 548722 190059 548725
rect 446438 548722 446444 548724
rect 189993 548720 446444 548722
rect 189993 548664 189998 548720
rect 190054 548664 446444 548720
rect 189993 548662 446444 548664
rect 189993 548659 190059 548662
rect 446438 548660 446444 548662
rect 446508 548660 446514 548724
rect 151854 548524 151860 548588
rect 151924 548586 151930 548588
rect 415025 548586 415091 548589
rect 151924 548584 415091 548586
rect 151924 548528 415030 548584
rect 415086 548528 415091 548584
rect 151924 548526 415091 548528
rect 151924 548524 151930 548526
rect 415025 548523 415091 548526
rect 166717 548450 166783 548453
rect 577773 548450 577839 548453
rect 166717 548448 577839 548450
rect 166717 548392 166722 548448
rect 166778 548392 577778 548448
rect 577834 548392 577839 548448
rect 166717 548390 577839 548392
rect 166717 548387 166783 548390
rect 577773 548387 577839 548390
rect 21357 548314 21423 548317
rect 435725 548314 435791 548317
rect 21357 548312 435791 548314
rect 21357 548256 21362 548312
rect 21418 548256 435730 548312
rect 435786 548256 435791 548312
rect 21357 548254 435791 548256
rect 21357 548251 21423 548254
rect 435725 548251 435791 548254
rect 158989 548178 159055 548181
rect 577589 548178 577655 548181
rect 158989 548176 577655 548178
rect 158989 548120 158994 548176
rect 159050 548120 577594 548176
rect 577650 548120 577655 548176
rect 158989 548118 577655 548120
rect 158989 548115 159055 548118
rect 577589 548115 577655 548118
rect 3693 548042 3759 548045
rect 425329 548042 425395 548045
rect 3693 548040 425395 548042
rect 3693 547984 3698 548040
rect 3754 547984 425334 548040
rect 425390 547984 425395 548040
rect 3693 547982 425395 547984
rect 3693 547979 3759 547982
rect 425329 547979 425395 547982
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 152222 545260 152228 545324
rect 152292 545322 152298 545324
rect 422477 545322 422543 545325
rect 152292 545320 422543 545322
rect 152292 545264 422482 545320
rect 422538 545264 422543 545320
rect 152292 545262 422543 545264
rect 152292 545260 152298 545262
rect 422477 545259 422543 545262
rect 152958 545124 152964 545188
rect 153028 545186 153034 545188
rect 430481 545186 430547 545189
rect 153028 545184 430547 545186
rect 153028 545128 430486 545184
rect 430542 545128 430547 545184
rect 153028 545126 430547 545128
rect 153028 545124 153034 545126
rect 430481 545123 430547 545126
rect 151537 544642 151603 544645
rect 154021 544644 154087 544645
rect 203149 544644 203215 544645
rect 205449 544644 205515 544645
rect 151670 544642 151676 544644
rect 151537 544640 151676 544642
rect 151537 544584 151542 544640
rect 151598 544584 151676 544640
rect 151537 544582 151676 544584
rect 151537 544579 151603 544582
rect 151670 544580 151676 544582
rect 151740 544580 151746 544644
rect 154021 544640 154068 544644
rect 154132 544642 154138 544644
rect 154021 544584 154026 544640
rect 154021 544580 154068 544584
rect 154132 544582 154178 544642
rect 203149 544640 203196 544644
rect 203260 544642 203266 544644
rect 205398 544642 205404 544644
rect 203149 544584 203154 544640
rect 154132 544580 154138 544582
rect 203149 544580 203196 544584
rect 203260 544582 203306 544642
rect 205358 544582 205404 544642
rect 205468 544640 205515 544644
rect 205510 544584 205515 544640
rect 203260 544580 203266 544582
rect 205398 544580 205404 544582
rect 205468 544580 205515 544584
rect 154021 544579 154087 544580
rect 203149 544579 203215 544580
rect 205449 544579 205515 544580
rect 208025 544642 208091 544645
rect 213453 544644 213519 544645
rect 208158 544642 208164 544644
rect 208025 544640 208164 544642
rect 208025 544584 208030 544640
rect 208086 544584 208164 544640
rect 208025 544582 208164 544584
rect 208025 544579 208091 544582
rect 208158 544580 208164 544582
rect 208228 544580 208234 544644
rect 213453 544640 213500 544644
rect 213564 544642 213570 544644
rect 221273 544642 221339 544645
rect 231577 544644 231643 544645
rect 386505 544644 386571 544645
rect 221406 544642 221412 544644
rect 213453 544584 213458 544640
rect 213453 544580 213500 544584
rect 213564 544582 213610 544642
rect 221273 544640 221412 544642
rect 221273 544584 221278 544640
rect 221334 544584 221412 544640
rect 221273 544582 221412 544584
rect 213564 544580 213570 544582
rect 213453 544579 213519 544580
rect 221273 544579 221339 544582
rect 221406 544580 221412 544582
rect 221476 544580 221482 544644
rect 231526 544642 231532 544644
rect 231486 544582 231532 544642
rect 231596 544640 231643 544644
rect 386454 544642 386460 544644
rect 231638 544584 231643 544640
rect 231526 544580 231532 544582
rect 231596 544580 231643 544584
rect 386414 544582 386460 544642
rect 386524 544640 386571 544644
rect 386566 544584 386571 544640
rect 386454 544580 386460 544582
rect 386524 544580 386571 544584
rect 231577 544579 231643 544580
rect 386505 544579 386571 544580
rect 226926 543900 226932 543964
rect 226996 543962 227002 543964
rect 231710 543962 231716 543964
rect 226996 543902 231716 543962
rect 226996 543900 227002 543902
rect 231710 543900 231716 543902
rect 231780 543900 231786 543964
rect 221406 543628 221412 543692
rect 221476 543690 221482 543692
rect 579613 543690 579679 543693
rect 221476 543688 579679 543690
rect 221476 543632 579618 543688
rect 579674 543632 579679 543688
rect 221476 543630 579679 543632
rect 221476 543628 221482 543630
rect 579613 543627 579679 543630
rect 213494 543492 213500 543556
rect 213564 543554 213570 543556
rect 579797 543554 579863 543557
rect 213564 543552 579863 543554
rect 213564 543496 579802 543552
rect 579858 543496 579863 543552
rect 213564 543494 579863 543496
rect 213564 543492 213570 543494
rect 579797 543491 579863 543494
rect 208158 543356 208164 543420
rect 208228 543418 208234 543420
rect 579981 543418 580047 543421
rect 208228 543416 580047 543418
rect 208228 543360 579986 543416
rect 580042 543360 580047 543416
rect 208228 543358 580047 543360
rect 208228 543356 208234 543358
rect 579981 543355 580047 543358
rect 205398 543220 205404 543284
rect 205468 543282 205474 543284
rect 226926 543282 226932 543284
rect 205468 543222 226932 543282
rect 205468 543220 205474 543222
rect 226926 543220 226932 543222
rect 226996 543220 227002 543284
rect 231526 543220 231532 543284
rect 231596 543220 231602 543284
rect 231710 543220 231716 543284
rect 231780 543282 231786 543284
rect 580165 543282 580231 543285
rect 231780 543280 580231 543282
rect 231780 543224 580170 543280
rect 580226 543224 580231 543280
rect 231780 543222 580231 543224
rect 231780 543220 231786 543222
rect 203190 543084 203196 543148
rect 203260 543146 203266 543148
rect 231158 543146 231164 543148
rect 203260 543086 231164 543146
rect 203260 543084 203266 543086
rect 231158 543084 231164 543086
rect 231228 543084 231234 543148
rect 3325 543010 3391 543013
rect 231342 543010 231348 543012
rect 3325 543008 231348 543010
rect 3325 542952 3330 543008
rect 3386 542952 231348 543008
rect 3325 542950 231348 542952
rect 3325 542947 3391 542950
rect 231342 542948 231348 542950
rect 231412 542948 231418 543012
rect 231534 542874 231594 543220
rect 580165 543219 580231 543222
rect 231894 543084 231900 543148
rect 231964 543146 231970 543148
rect 580809 543146 580875 543149
rect 231964 543144 580875 543146
rect 231964 543088 580814 543144
rect 580870 543088 580875 543144
rect 231964 543086 580875 543088
rect 231964 543084 231970 543086
rect 580809 543083 580875 543086
rect 231710 542948 231716 543012
rect 231780 543010 231786 543012
rect 386454 543010 386460 543012
rect 231780 542950 386460 543010
rect 231780 542948 231786 542950
rect 386454 542948 386460 542950
rect 386524 542948 386530 543012
rect 449801 542874 449867 542877
rect 231534 542872 449867 542874
rect 231534 542816 449806 542872
rect 449862 542816 449867 542872
rect 231534 542814 449867 542816
rect 449801 542811 449867 542814
rect -960 538658 480 538748
rect 2957 538658 3023 538661
rect -960 538656 3023 538658
rect -960 538600 2962 538656
rect 3018 538600 3023 538656
rect -960 538598 3023 538600
rect -960 538508 480 538598
rect 2957 538595 3023 538598
rect 152222 536148 152228 536212
rect 152292 536210 152298 536212
rect 152958 536210 152964 536212
rect 152292 536150 152964 536210
rect 152292 536148 152298 536150
rect 152958 536148 152964 536150
rect 153028 536148 153034 536212
rect 579889 533898 579955 533901
rect 583520 533898 584960 533988
rect 579889 533896 584960 533898
rect 579889 533840 579894 533896
rect 579950 533840 584960 533896
rect 579889 533838 584960 533840
rect 579889 533835 579955 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 152774 521658 152780 521660
rect 152598 521598 152780 521658
rect 152598 520300 152658 521598
rect 152774 521596 152780 521598
rect 152844 521596 152850 521660
rect 152590 520236 152596 520300
rect 152660 520236 152666 520300
rect 152038 520100 152044 520164
rect 152108 520162 152114 520164
rect 152590 520162 152596 520164
rect 152108 520102 152596 520162
rect 152108 520100 152114 520102
rect 152590 520100 152596 520102
rect 152660 520100 152666 520164
rect 150750 511940 150756 512004
rect 150820 512002 150826 512004
rect 151486 512002 151492 512004
rect 150820 511942 151492 512002
rect 150820 511940 150826 511942
rect 151486 511940 151492 511942
rect 151556 511940 151562 512004
rect 152038 510580 152044 510644
rect 152108 510642 152114 510644
rect 152774 510642 152780 510644
rect 152108 510582 152780 510642
rect 152108 510580 152114 510582
rect 152774 510580 152780 510582
rect 152844 510580 152850 510644
rect 152958 510506 152964 510508
rect 152782 510446 152964 510506
rect 152782 510098 152842 510446
rect 152958 510444 152964 510446
rect 153028 510444 153034 510508
rect 579889 510370 579955 510373
rect 583520 510370 584960 510460
rect 579889 510368 584960 510370
rect 579889 510312 579894 510368
rect 579950 510312 584960 510368
rect 579889 510310 584960 510312
rect 579889 510307 579955 510310
rect 583520 510220 584960 510310
rect 152958 510098 152964 510100
rect -960 509962 480 510052
rect 152782 510038 152964 510098
rect 152958 510036 152964 510038
rect 153028 510036 153034 510100
rect 2957 509962 3023 509965
rect -960 509960 3023 509962
rect -960 509904 2962 509960
rect 3018 509904 3023 509960
rect -960 509902 3023 509904
rect -960 509812 480 509902
rect 2957 509899 3023 509902
rect 150750 502556 150756 502620
rect 150820 502618 150826 502620
rect 150820 502558 151186 502618
rect 150820 502556 150826 502558
rect 151126 502484 151186 502558
rect 151118 502420 151124 502484
rect 151188 502420 151194 502484
rect 580073 498674 580139 498677
rect 583520 498674 584960 498764
rect 580073 498672 584960 498674
rect 580073 498616 580078 498672
rect 580134 498616 584960 498672
rect 580073 498614 584960 498616
rect 580073 498611 580139 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2773 495546 2839 495549
rect -960 495544 2839 495546
rect -960 495488 2778 495544
rect 2834 495488 2839 495544
rect -960 495486 2839 495488
rect -960 495396 480 495486
rect 2773 495483 2839 495486
rect 152590 491404 152596 491468
rect 152660 491466 152666 491468
rect 152660 491406 152842 491466
rect 152660 491404 152666 491406
rect 152782 491332 152842 491406
rect 152774 491268 152780 491332
rect 152844 491268 152850 491332
rect 152774 491132 152780 491196
rect 152844 491194 152850 491196
rect 152844 491134 153026 491194
rect 152844 491132 152850 491134
rect 152038 490860 152044 490924
rect 152108 490922 152114 490924
rect 152966 490922 153026 491134
rect 152108 490862 153026 490922
rect 152108 490860 152114 490862
rect 580073 486842 580139 486845
rect 583520 486842 584960 486932
rect 580073 486840 584960 486842
rect 580073 486784 580078 486840
rect 580134 486784 584960 486840
rect 580073 486782 584960 486784
rect 580073 486779 580139 486782
rect 583520 486692 584960 486782
rect 152038 481612 152044 481676
rect 152108 481674 152114 481676
rect 152774 481674 152780 481676
rect 152108 481614 152780 481674
rect 152108 481612 152114 481614
rect 152774 481612 152780 481614
rect 152844 481612 152850 481676
rect 152222 481476 152228 481540
rect 152292 481538 152298 481540
rect 152774 481538 152780 481540
rect 152292 481478 152780 481538
rect 152292 481476 152298 481478
rect 152774 481476 152780 481478
rect 152844 481476 152850 481540
rect -960 481130 480 481220
rect 2773 481130 2839 481133
rect -960 481128 2839 481130
rect -960 481072 2778 481128
rect 2834 481072 2839 481128
rect -960 481070 2839 481072
rect -960 480980 480 481070
rect 2773 481067 2839 481070
rect 583520 474996 584960 475236
rect 152222 471956 152228 472020
rect 152292 472018 152298 472020
rect 152774 472018 152780 472020
rect 152292 471958 152780 472018
rect 152292 471956 152298 471958
rect 152774 471956 152780 471958
rect 152844 471956 152850 472020
rect -960 466700 480 466940
rect 152774 463524 152780 463588
rect 152844 463586 152850 463588
rect 153142 463586 153148 463588
rect 152844 463526 153148 463586
rect 152844 463524 152850 463526
rect 153142 463524 153148 463526
rect 153212 463524 153218 463588
rect 580073 463450 580139 463453
rect 583520 463450 584960 463540
rect 580073 463448 584960 463450
rect 580073 463392 580078 463448
rect 580134 463392 584960 463448
rect 580073 463390 584960 463392
rect 580073 463387 580139 463390
rect 583520 463300 584960 463390
rect 151486 456922 151492 456924
rect 151310 456862 151492 456922
rect 151310 456652 151370 456862
rect 151486 456860 151492 456862
rect 151556 456860 151562 456924
rect 151302 456588 151308 456652
rect 151372 456588 151378 456652
rect 152774 454140 152780 454204
rect 152844 454202 152850 454204
rect 153142 454202 153148 454204
rect 152844 454142 153148 454202
rect 152844 454140 152850 454142
rect 153142 454140 153148 454142
rect 153212 454140 153218 454204
rect -960 452434 480 452524
rect 152222 452508 152228 452572
rect 152292 452570 152298 452572
rect 152774 452570 152780 452572
rect 152292 452510 152780 452570
rect 152292 452508 152298 452510
rect 152774 452508 152780 452510
rect 152844 452508 152850 452572
rect 3049 452434 3115 452437
rect -960 452432 3115 452434
rect -960 452376 3054 452432
rect 3110 452376 3115 452432
rect -960 452374 3115 452376
rect -960 452284 480 452374
rect 3049 452371 3115 452374
rect 580073 451754 580139 451757
rect 583520 451754 584960 451844
rect 580073 451752 584960 451754
rect 580073 451696 580078 451752
rect 580134 451696 584960 451752
rect 580073 451694 584960 451696
rect 580073 451691 580139 451694
rect 583520 451604 584960 451694
rect 151302 447204 151308 447268
rect 151372 447204 151378 447268
rect 151310 446994 151370 447204
rect 151486 446994 151492 446996
rect 151310 446934 151492 446994
rect 151486 446932 151492 446934
rect 151556 446932 151562 446996
rect 152222 443124 152228 443188
rect 152292 443186 152298 443188
rect 152292 443126 152658 443186
rect 152292 443124 152298 443126
rect 152598 443052 152658 443126
rect 152590 442988 152596 443052
rect 152660 442988 152666 443052
rect 151486 441492 151492 441556
rect 151556 441492 151562 441556
rect 150934 441356 150940 441420
rect 151004 441418 151010 441420
rect 151494 441418 151554 441492
rect 151004 441358 151554 441418
rect 151004 441356 151010 441358
rect 579613 439922 579679 439925
rect 583520 439922 584960 440012
rect 579613 439920 584960 439922
rect 579613 439864 579618 439920
rect 579674 439864 584960 439920
rect 579613 439862 584960 439864
rect 579613 439859 579679 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 2773 438018 2839 438021
rect -960 438016 2839 438018
rect -960 437960 2778 438016
rect 2834 437960 2839 438016
rect -960 437958 2839 437960
rect -960 437868 480 437958
rect 2773 437955 2839 437958
rect 150934 431972 150940 432036
rect 151004 432034 151010 432036
rect 151670 432034 151676 432036
rect 151004 431974 151676 432034
rect 151004 431972 151010 431974
rect 151670 431972 151676 431974
rect 151740 431972 151746 432036
rect 583520 428076 584960 428316
rect 151670 427892 151676 427956
rect 151740 427892 151746 427956
rect 151678 427820 151738 427892
rect 151670 427756 151676 427820
rect 151740 427756 151746 427820
rect -960 423738 480 423828
rect 2773 423738 2839 423741
rect -960 423736 2839 423738
rect -960 423680 2778 423736
rect 2834 423680 2839 423736
rect -960 423678 2839 423680
rect -960 423588 480 423678
rect 2773 423675 2839 423678
rect 151670 423676 151676 423740
rect 151740 423676 151746 423740
rect 151678 423604 151738 423676
rect 151670 423540 151676 423604
rect 151740 423540 151746 423604
rect 152222 423540 152228 423604
rect 152292 423602 152298 423604
rect 152774 423602 152780 423604
rect 152292 423542 152780 423602
rect 152292 423540 152298 423542
rect 152774 423540 152780 423542
rect 152844 423540 152850 423604
rect 580073 416530 580139 416533
rect 583520 416530 584960 416620
rect 580073 416528 584960 416530
rect 580073 416472 580078 416528
rect 580134 416472 584960 416528
rect 580073 416470 584960 416472
rect 580073 416467 580139 416470
rect 583520 416380 584960 416470
rect 152222 414156 152228 414220
rect 152292 414218 152298 414220
rect 152292 414158 152842 414218
rect 152292 414156 152298 414158
rect 152782 414084 152842 414158
rect 152774 414020 152780 414084
rect 152844 414020 152850 414084
rect 151302 412524 151308 412588
rect 151372 412524 151378 412588
rect 151310 412450 151370 412524
rect 151486 412450 151492 412452
rect 151310 412390 151492 412450
rect 151486 412388 151492 412390
rect 151556 412388 151562 412452
rect -960 409172 480 409412
rect 580073 404834 580139 404837
rect 583520 404834 584960 404924
rect 580073 404832 584960 404834
rect 580073 404776 580078 404832
rect 580134 404776 584960 404832
rect 580073 404774 584960 404776
rect 580073 404771 580139 404774
rect 583520 404684 584960 404774
rect 152222 404228 152228 404292
rect 152292 404290 152298 404292
rect 152774 404290 152780 404292
rect 152292 404230 152780 404290
rect 152292 404228 152298 404230
rect 152774 404228 152780 404230
rect 152844 404228 152850 404292
rect 151486 402868 151492 402932
rect 151556 402868 151562 402932
rect 151118 402732 151124 402796
rect 151188 402794 151194 402796
rect 151494 402794 151554 402868
rect 151188 402734 151554 402794
rect 151188 402732 151194 402734
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 152222 394844 152228 394908
rect 152292 394906 152298 394908
rect 152292 394846 152842 394906
rect 152292 394844 152298 394846
rect 152782 394772 152842 394846
rect 152774 394708 152780 394772
rect 152844 394708 152850 394772
rect 151118 393348 151124 393412
rect 151188 393410 151194 393412
rect 151670 393410 151676 393412
rect 151188 393350 151676 393410
rect 151188 393348 151194 393350
rect 151670 393348 151676 393350
rect 151740 393348 151746 393412
rect 579797 393002 579863 393005
rect 583520 393002 584960 393092
rect 579797 393000 584960 393002
rect 579797 392944 579802 393000
rect 579858 392944 584960 393000
rect 579797 392942 584960 392944
rect 579797 392939 579863 392942
rect 583520 392852 584960 392942
rect 151670 389330 151676 389332
rect 151494 389270 151676 389330
rect 151494 389060 151554 389270
rect 151670 389268 151676 389270
rect 151740 389268 151746 389332
rect 151486 388996 151492 389060
rect 151556 388996 151562 389060
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 2957 380626 3023 380629
rect -960 380624 3023 380626
rect -960 380568 2962 380624
rect 3018 380568 3023 380624
rect -960 380566 3023 380568
rect -960 380476 480 380566
rect 2957 380563 3023 380566
rect 579981 369610 580047 369613
rect 583520 369610 584960 369700
rect 579981 369608 584960 369610
rect 579981 369552 579986 369608
rect 580042 369552 584960 369608
rect 579981 369550 584960 369552
rect 579981 369547 580047 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 2773 366210 2839 366213
rect -960 366208 2839 366210
rect -960 366152 2778 366208
rect 2834 366152 2839 366208
rect -960 366150 2839 366152
rect -960 366060 480 366150
rect 2773 366147 2839 366150
rect 152222 365604 152228 365668
rect 152292 365666 152298 365668
rect 152774 365666 152780 365668
rect 152292 365606 152780 365666
rect 152292 365604 152298 365606
rect 152774 365604 152780 365606
rect 152844 365604 152850 365668
rect 151486 364380 151492 364444
rect 151556 364442 151562 364444
rect 151670 364442 151676 364444
rect 151556 364382 151676 364442
rect 151556 364380 151562 364382
rect 151670 364380 151676 364382
rect 151740 364380 151746 364444
rect 583520 357914 584960 358004
rect 583342 357854 584960 357914
rect 447726 357716 447732 357780
rect 447796 357778 447802 357780
rect 447796 357718 451290 357778
rect 447796 357716 447802 357718
rect 451230 357642 451290 357718
rect 460982 357718 470610 357778
rect 451230 357582 460858 357642
rect 460798 357506 460858 357582
rect 460982 357506 461042 357718
rect 470550 357642 470610 357718
rect 480302 357718 489930 357778
rect 470550 357582 480178 357642
rect 460798 357446 461042 357506
rect 480118 357506 480178 357582
rect 480302 357506 480362 357718
rect 489870 357642 489930 357718
rect 499622 357718 509250 357778
rect 489870 357582 499498 357642
rect 480118 357446 480362 357506
rect 499438 357506 499498 357582
rect 499622 357506 499682 357718
rect 509190 357642 509250 357718
rect 518942 357718 528570 357778
rect 509190 357582 518818 357642
rect 499438 357446 499682 357506
rect 518758 357506 518818 357582
rect 518942 357506 519002 357718
rect 528510 357642 528570 357718
rect 538262 357718 547890 357778
rect 528510 357582 538138 357642
rect 518758 357446 519002 357506
rect 538078 357506 538138 357582
rect 538262 357506 538322 357718
rect 547830 357642 547890 357718
rect 557582 357718 567210 357778
rect 547830 357582 557458 357642
rect 538078 357446 538322 357506
rect 557398 357506 557458 357582
rect 557582 357506 557642 357718
rect 567150 357642 567210 357718
rect 583342 357642 583402 357854
rect 583520 357764 584960 357854
rect 567150 357582 576778 357642
rect 557398 357446 557642 357506
rect 576718 357506 576778 357582
rect 576902 357582 583402 357642
rect 576902 357506 576962 357582
rect 576718 357446 576962 357506
rect 151670 356282 151676 356284
rect 151494 356222 151676 356282
rect 151494 356148 151554 356222
rect 151670 356220 151676 356222
rect 151740 356220 151746 356284
rect 152222 356220 152228 356284
rect 152292 356282 152298 356284
rect 152292 356222 152842 356282
rect 152292 356220 152298 356222
rect 152782 356148 152842 356222
rect 151486 356084 151492 356148
rect 151556 356084 151562 356148
rect 152774 356084 152780 356148
rect 152844 356084 152850 356148
rect -960 351780 480 352020
rect 151486 348468 151492 348532
rect 151556 348530 151562 348532
rect 152222 348530 152228 348532
rect 151556 348470 152228 348530
rect 151556 348468 151562 348470
rect 152222 348468 152228 348470
rect 152292 348468 152298 348532
rect 151854 346564 151860 346628
rect 151924 346564 151930 346628
rect 151862 346220 151922 346564
rect 151854 346156 151860 346220
rect 151924 346156 151930 346220
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 3233 337514 3299 337517
rect -960 337512 3299 337514
rect -960 337456 3238 337512
rect 3294 337456 3299 337512
rect -960 337454 3299 337456
rect -960 337364 480 337454
rect 3233 337451 3299 337454
rect 152038 335412 152044 335476
rect 152108 335474 152114 335476
rect 152222 335474 152228 335476
rect 152108 335414 152228 335474
rect 152108 335412 152114 335414
rect 152222 335412 152228 335414
rect 152292 335412 152298 335476
rect 151854 335276 151860 335340
rect 151924 335338 151930 335340
rect 151924 335278 152290 335338
rect 151924 335276 151930 335278
rect 152230 335204 152290 335278
rect 152038 335140 152044 335204
rect 152108 335140 152114 335204
rect 152222 335140 152228 335204
rect 152292 335140 152298 335204
rect 151854 334052 151860 334116
rect 151924 334114 151930 334116
rect 152046 334114 152106 335140
rect 583520 334236 584960 334476
rect 151924 334054 152106 334114
rect 151924 334052 151930 334054
rect 152774 327524 152780 327588
rect 152844 327524 152850 327588
rect 152958 327524 152964 327588
rect 153028 327524 153034 327588
rect 151854 327450 151860 327452
rect 151494 327390 151860 327450
rect 151494 327180 151554 327390
rect 151854 327388 151860 327390
rect 151924 327388 151930 327452
rect 152782 327180 152842 327524
rect 152966 327180 153026 327524
rect 151486 327116 151492 327180
rect 151556 327116 151562 327180
rect 152774 327116 152780 327180
rect 152844 327116 152850 327180
rect 152958 327116 152964 327180
rect 153028 327116 153034 327180
rect 152222 326980 152228 327044
rect 152292 327042 152298 327044
rect 152774 327042 152780 327044
rect 152292 326982 152780 327042
rect 152292 326980 152298 326982
rect 152774 326980 152780 326982
rect 152844 326980 152850 327044
rect 150750 325620 150756 325684
rect 150820 325682 150826 325684
rect 151486 325682 151492 325684
rect 150820 325622 151492 325682
rect 150820 325620 150826 325622
rect 151486 325620 151492 325622
rect 151556 325620 151562 325684
rect -960 323098 480 323188
rect 3141 323098 3207 323101
rect -960 323096 3207 323098
rect -960 323040 3146 323096
rect 3202 323040 3207 323096
rect -960 323038 3207 323040
rect -960 322948 480 323038
rect 3141 323035 3207 323038
rect 580901 322690 580967 322693
rect 583520 322690 584960 322780
rect 580901 322688 584960 322690
rect 580901 322632 580906 322688
rect 580962 322632 584960 322688
rect 580901 322630 584960 322632
rect 580901 322627 580967 322630
rect 583520 322540 584960 322630
rect 152222 317596 152228 317660
rect 152292 317658 152298 317660
rect 152292 317598 152842 317658
rect 152292 317596 152298 317598
rect 152782 317524 152842 317598
rect 152774 317460 152780 317524
rect 152844 317460 152850 317524
rect 150750 316236 150756 316300
rect 150820 316298 150826 316300
rect 151302 316298 151308 316300
rect 150820 316238 151308 316298
rect 150820 316236 150826 316238
rect 151302 316236 151308 316238
rect 151372 316236 151378 316300
rect 151302 315964 151308 316028
rect 151372 316026 151378 316028
rect 151486 316026 151492 316028
rect 151372 315966 151492 316026
rect 151372 315964 151378 315966
rect 151486 315964 151492 315966
rect 151556 315964 151562 316028
rect 151302 314604 151308 314668
rect 151372 314666 151378 314668
rect 151486 314666 151492 314668
rect 151372 314606 151492 314666
rect 151372 314604 151378 314606
rect 151486 314604 151492 314606
rect 151556 314604 151562 314668
rect 580809 310858 580875 310861
rect 583520 310858 584960 310948
rect 580809 310856 584960 310858
rect 580809 310800 580814 310856
rect 580870 310800 584960 310856
rect 580809 310798 584960 310800
rect 580809 310795 580875 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 152222 307668 152228 307732
rect 152292 307730 152298 307732
rect 152774 307730 152780 307732
rect 152292 307670 152780 307730
rect 152292 307668 152298 307670
rect 152774 307668 152780 307670
rect 152844 307668 152850 307732
rect 151118 304948 151124 305012
rect 151188 305010 151194 305012
rect 151302 305010 151308 305012
rect 151188 304950 151308 305010
rect 151188 304948 151194 304950
rect 151302 304948 151308 304950
rect 151372 304948 151378 305012
rect 583520 299162 584960 299252
rect 583342 299102 584960 299162
rect 446622 298420 446628 298484
rect 446692 298482 446698 298484
rect 446692 298422 451290 298482
rect 446692 298420 446698 298422
rect 152222 298284 152228 298348
rect 152292 298346 152298 298348
rect 451230 298346 451290 298422
rect 460982 298422 470610 298482
rect 152292 298286 152842 298346
rect 451230 298286 460858 298346
rect 152292 298284 152298 298286
rect 152782 298212 152842 298286
rect 152774 298148 152780 298212
rect 152844 298148 152850 298212
rect 460798 298210 460858 298286
rect 460982 298210 461042 298422
rect 470550 298346 470610 298422
rect 480302 298422 489930 298482
rect 470550 298286 480178 298346
rect 460798 298150 461042 298210
rect 480118 298210 480178 298286
rect 480302 298210 480362 298422
rect 489870 298346 489930 298422
rect 499622 298422 509250 298482
rect 489870 298286 499498 298346
rect 480118 298150 480362 298210
rect 499438 298210 499498 298286
rect 499622 298210 499682 298422
rect 509190 298346 509250 298422
rect 518942 298422 528570 298482
rect 509190 298286 518818 298346
rect 499438 298150 499682 298210
rect 518758 298210 518818 298286
rect 518942 298210 519002 298422
rect 528510 298346 528570 298422
rect 538262 298422 547890 298482
rect 528510 298286 538138 298346
rect 518758 298150 519002 298210
rect 538078 298210 538138 298286
rect 538262 298210 538322 298422
rect 547830 298346 547890 298422
rect 557582 298422 567210 298482
rect 547830 298286 557458 298346
rect 538078 298150 538322 298210
rect 557398 298210 557458 298286
rect 557582 298210 557642 298422
rect 567150 298346 567210 298422
rect 583342 298346 583402 299102
rect 583520 299012 584960 299102
rect 567150 298286 576778 298346
rect 557398 298150 557642 298210
rect 576718 298210 576778 298286
rect 576902 298286 583402 298346
rect 576902 298210 576962 298286
rect 576718 298150 576962 298210
rect 151118 296788 151124 296852
rect 151188 296850 151194 296852
rect 151670 296850 151676 296852
rect 151188 296790 151676 296850
rect 151188 296788 151194 296790
rect 151670 296788 151676 296790
rect 151740 296788 151746 296852
rect -960 294402 480 294492
rect 4061 294402 4127 294405
rect -960 294400 4127 294402
rect -960 294344 4066 294400
rect 4122 294344 4127 294400
rect -960 294342 4127 294344
rect -960 294252 480 294342
rect 4061 294339 4127 294342
rect 151670 292770 151676 292772
rect 151494 292710 151676 292770
rect 151494 292500 151554 292710
rect 151670 292708 151676 292710
rect 151740 292708 151746 292772
rect 151486 292436 151492 292500
rect 151556 292436 151562 292500
rect 152222 288356 152228 288420
rect 152292 288418 152298 288420
rect 152774 288418 152780 288420
rect 152292 288358 152780 288418
rect 152292 288356 152298 288358
rect 152774 288356 152780 288358
rect 152844 288356 152850 288420
rect 583520 287316 584960 287556
rect 151118 280740 151124 280804
rect 151188 280802 151194 280804
rect 151486 280802 151492 280804
rect 151188 280742 151492 280802
rect 151188 280740 151194 280742
rect 151486 280740 151492 280742
rect 151556 280740 151562 280804
rect -960 280122 480 280212
rect 3141 280122 3207 280125
rect -960 280120 3207 280122
rect -960 280064 3146 280120
rect 3202 280064 3207 280120
rect -960 280062 3207 280064
rect -960 279972 480 280062
rect 3141 280059 3207 280062
rect 152222 278972 152228 279036
rect 152292 279034 152298 279036
rect 152292 278974 152842 279034
rect 152292 278972 152298 278974
rect 152782 278900 152842 278974
rect 152774 278836 152780 278900
rect 152844 278836 152850 278900
rect 151118 275980 151124 276044
rect 151188 276042 151194 276044
rect 151486 276042 151492 276044
rect 151188 275982 151492 276042
rect 151188 275980 151194 275982
rect 151486 275980 151492 275982
rect 151556 275980 151562 276044
rect 580717 275770 580783 275773
rect 583520 275770 584960 275860
rect 580717 275768 584960 275770
rect 580717 275712 580722 275768
rect 580778 275712 584960 275768
rect 580717 275710 584960 275712
rect 580717 275707 580783 275710
rect 583520 275620 584960 275710
rect 151118 266188 151124 266252
rect 151188 266250 151194 266252
rect 151486 266250 151492 266252
rect 151188 266190 151492 266250
rect 151188 266188 151194 266190
rect 151486 266188 151492 266190
rect 151556 266188 151562 266252
rect -960 265706 480 265796
rect 2773 265706 2839 265709
rect -960 265704 2839 265706
rect -960 265648 2778 265704
rect 2834 265648 2839 265704
rect -960 265646 2839 265648
rect -960 265556 480 265646
rect 2773 265643 2839 265646
rect 580625 263938 580691 263941
rect 583520 263938 584960 264028
rect 580625 263936 584960 263938
rect 580625 263880 580630 263936
rect 580686 263880 584960 263936
rect 580625 263878 584960 263880
rect 580625 263875 580691 263878
rect 583520 263788 584960 263878
rect 152774 259388 152780 259452
rect 152844 259388 152850 259452
rect 152590 259252 152596 259316
rect 152660 259314 152666 259316
rect 152782 259314 152842 259388
rect 152660 259254 152842 259314
rect 152660 259252 152666 259254
rect 151118 256668 151124 256732
rect 151188 256730 151194 256732
rect 151486 256730 151492 256732
rect 151188 256670 151492 256730
rect 151188 256668 151194 256670
rect 151486 256668 151492 256670
rect 151556 256668 151562 256732
rect 583520 252242 584960 252332
rect 583342 252182 584960 252242
rect 446806 251500 446812 251564
rect 446876 251562 446882 251564
rect 446876 251502 451290 251562
rect 446876 251500 446882 251502
rect 451230 251426 451290 251502
rect 460982 251502 470610 251562
rect -960 251290 480 251380
rect 451230 251366 460858 251426
rect 3969 251290 4035 251293
rect -960 251288 4035 251290
rect -960 251232 3974 251288
rect 4030 251232 4035 251288
rect -960 251230 4035 251232
rect 460798 251290 460858 251366
rect 460982 251290 461042 251502
rect 470550 251426 470610 251502
rect 480302 251502 489930 251562
rect 470550 251366 480178 251426
rect 460798 251230 461042 251290
rect 480118 251290 480178 251366
rect 480302 251290 480362 251502
rect 489870 251426 489930 251502
rect 499622 251502 509250 251562
rect 489870 251366 499498 251426
rect 480118 251230 480362 251290
rect 499438 251290 499498 251366
rect 499622 251290 499682 251502
rect 509190 251426 509250 251502
rect 518942 251502 528570 251562
rect 509190 251366 518818 251426
rect 499438 251230 499682 251290
rect 518758 251290 518818 251366
rect 518942 251290 519002 251502
rect 528510 251426 528570 251502
rect 538262 251502 547890 251562
rect 528510 251366 538138 251426
rect 518758 251230 519002 251290
rect 538078 251290 538138 251366
rect 538262 251290 538322 251502
rect 547830 251426 547890 251502
rect 557582 251502 567210 251562
rect 547830 251366 557458 251426
rect 538078 251230 538322 251290
rect 557398 251290 557458 251366
rect 557582 251290 557642 251502
rect 567150 251426 567210 251502
rect 583342 251426 583402 252182
rect 583520 252092 584960 252182
rect 567150 251366 576778 251426
rect 557398 251230 557642 251290
rect 576718 251290 576778 251366
rect 576902 251366 583402 251426
rect 576902 251290 576962 251366
rect 576718 251230 576962 251290
rect -960 251140 480 251230
rect 3969 251227 4035 251230
rect 152590 248508 152596 248572
rect 152660 248508 152666 248572
rect 152598 248434 152658 248508
rect 152774 248434 152780 248436
rect 152598 248374 152780 248434
rect 152774 248372 152780 248374
rect 152844 248372 152850 248436
rect 152774 248236 152780 248300
rect 152844 248298 152850 248300
rect 153510 248298 153516 248300
rect 152844 248238 153516 248298
rect 152844 248236 152850 248238
rect 153510 248236 153516 248238
rect 153580 248236 153586 248300
rect 151118 246876 151124 246940
rect 151188 246938 151194 246940
rect 151486 246938 151492 246940
rect 151188 246878 151492 246938
rect 151188 246876 151194 246878
rect 151486 246876 151492 246878
rect 151556 246876 151562 246940
rect 152958 244428 152964 244492
rect 153028 244428 153034 244492
rect 152966 244220 153026 244428
rect 152958 244156 152964 244220
rect 153028 244156 153034 244220
rect 367093 242722 367159 242725
rect 374269 242722 374335 242725
rect 367093 242720 374335 242722
rect 367093 242664 367098 242720
rect 367154 242664 374274 242720
rect 374330 242664 374335 242720
rect 367093 242662 374335 242664
rect 367093 242659 367159 242662
rect 374269 242659 374335 242662
rect 367093 242586 367159 242589
rect 367461 242586 367527 242589
rect 367093 242584 367527 242586
rect 367093 242528 367098 242584
rect 367154 242528 367466 242584
rect 367522 242528 367527 242584
rect 367093 242526 367527 242528
rect 367093 242523 367159 242526
rect 367461 242523 367527 242526
rect 367185 242450 367251 242453
rect 369577 242450 369643 242453
rect 367185 242448 369643 242450
rect 367185 242392 367190 242448
rect 367246 242392 369582 242448
rect 369638 242392 369643 242448
rect 367185 242390 369643 242392
rect 367185 242387 367251 242390
rect 369577 242387 369643 242390
rect 357525 242314 357591 242317
rect 367001 242314 367067 242317
rect 357525 242312 367067 242314
rect 357525 242256 357530 242312
rect 357586 242256 367006 242312
rect 367062 242256 367067 242312
rect 357525 242254 367067 242256
rect 357525 242251 357591 242254
rect 367001 242251 367067 242254
rect 13077 242178 13143 242181
rect 153285 242178 153351 242181
rect 13077 242176 153351 242178
rect 13077 242120 13082 242176
rect 13138 242120 153290 242176
rect 153346 242120 153351 242176
rect 13077 242118 153351 242120
rect 13077 242115 13143 242118
rect 153285 242115 153351 242118
rect 213821 242178 213887 242181
rect 259545 242178 259611 242181
rect 213821 242176 259611 242178
rect 213821 242120 213826 242176
rect 213882 242120 259550 242176
rect 259606 242120 259611 242176
rect 213821 242118 259611 242120
rect 213821 242115 213887 242118
rect 259545 242115 259611 242118
rect 353661 242178 353727 242181
rect 388437 242178 388503 242181
rect 353661 242176 388503 242178
rect 353661 242120 353666 242176
rect 353722 242120 388442 242176
rect 388498 242120 388503 242176
rect 353661 242118 388503 242120
rect 353661 242115 353727 242118
rect 388437 242115 388503 242118
rect 417785 242178 417851 242181
rect 511257 242178 511323 242181
rect 417785 242176 511323 242178
rect 417785 242120 417790 242176
rect 417846 242120 511262 242176
rect 511318 242120 511323 242176
rect 417785 242118 511323 242120
rect 417785 242115 417851 242118
rect 511257 242115 511323 242118
rect 367645 241770 367711 241773
rect 367645 241768 374194 241770
rect 367645 241712 367650 241768
rect 367706 241712 374194 241768
rect 367645 241710 374194 241712
rect 367645 241707 367711 241710
rect 268469 241634 268535 241637
rect 270585 241634 270651 241637
rect 268469 241632 270651 241634
rect 268469 241576 268474 241632
rect 268530 241576 270590 241632
rect 270646 241576 270651 241632
rect 268469 241574 270651 241576
rect 268469 241571 268535 241574
rect 270585 241571 270651 241574
rect 374134 241532 374194 241710
rect 374269 241532 374335 241535
rect 374134 241530 374335 241532
rect 179689 241498 179755 241501
rect 179873 241498 179939 241501
rect 179689 241496 179939 241498
rect 179689 241440 179694 241496
rect 179750 241440 179878 241496
rect 179934 241440 179939 241496
rect 179689 241438 179939 241440
rect 179689 241435 179755 241438
rect 179873 241435 179939 241438
rect 185209 241498 185275 241501
rect 185393 241498 185459 241501
rect 185209 241496 185459 241498
rect 185209 241440 185214 241496
rect 185270 241440 185398 241496
rect 185454 241440 185459 241496
rect 374134 241474 374274 241530
rect 374330 241474 374335 241530
rect 374134 241472 374335 241474
rect 374269 241469 374335 241472
rect 393773 241498 393839 241501
rect 394049 241498 394115 241501
rect 393773 241496 394115 241498
rect 185209 241438 185459 241440
rect 185209 241435 185275 241438
rect 185393 241435 185459 241438
rect 393773 241440 393778 241496
rect 393834 241440 394054 241496
rect 394110 241440 394115 241496
rect 393773 241438 394115 241440
rect 393773 241435 393839 241438
rect 394049 241435 394115 241438
rect 583520 240396 584960 240636
rect 238477 240138 238543 240141
rect 238661 240138 238727 240141
rect 238477 240136 238727 240138
rect 238477 240080 238482 240136
rect 238538 240080 238666 240136
rect 238722 240080 238727 240136
rect 238477 240078 238727 240080
rect 238477 240075 238543 240078
rect 238661 240075 238727 240078
rect 374269 240138 374335 240141
rect 374453 240138 374519 240141
rect 374269 240136 374519 240138
rect 374269 240080 374274 240136
rect 374330 240080 374458 240136
rect 374514 240080 374519 240136
rect 374269 240078 374519 240080
rect 374269 240075 374335 240078
rect 374453 240075 374519 240078
rect 153142 238716 153148 238780
rect 153212 238778 153218 238780
rect 153510 238778 153516 238780
rect 153212 238718 153516 238778
rect 153212 238716 153218 238718
rect 153510 238716 153516 238718
rect 153580 238716 153586 238780
rect 151118 237356 151124 237420
rect 151188 237418 151194 237420
rect 151486 237418 151492 237420
rect 151188 237358 151492 237418
rect 151188 237356 151194 237358
rect 151486 237356 151492 237358
rect 151556 237356 151562 237420
rect 151486 237220 151492 237284
rect 151556 237220 151562 237284
rect 151494 237146 151554 237220
rect 151721 237146 151787 237149
rect 151494 237144 151787 237146
rect -960 237010 480 237100
rect 151494 237088 151726 237144
rect 151782 237088 151787 237144
rect 151494 237086 151787 237088
rect 151721 237083 151787 237086
rect 3049 237010 3115 237013
rect -960 237008 3115 237010
rect -960 236952 3054 237008
rect 3110 236952 3115 237008
rect -960 236950 3115 236952
rect -960 236860 480 236950
rect 3049 236947 3115 236950
rect 179597 231842 179663 231845
rect 179781 231842 179847 231845
rect 179597 231840 179847 231842
rect 179597 231784 179602 231840
rect 179658 231784 179786 231840
rect 179842 231784 179847 231840
rect 179597 231782 179847 231784
rect 179597 231779 179663 231782
rect 179781 231779 179847 231782
rect 185117 231842 185183 231845
rect 185301 231842 185367 231845
rect 185117 231840 185367 231842
rect 185117 231784 185122 231840
rect 185178 231784 185306 231840
rect 185362 231784 185367 231840
rect 185117 231782 185367 231784
rect 185117 231779 185183 231782
rect 185301 231779 185367 231782
rect 223757 231842 223823 231845
rect 223941 231842 224007 231845
rect 223757 231840 224007 231842
rect 223757 231784 223762 231840
rect 223818 231784 223946 231840
rect 224002 231784 224007 231840
rect 223757 231782 224007 231784
rect 223757 231779 223823 231782
rect 223941 231779 224007 231782
rect 225045 231842 225111 231845
rect 225229 231842 225295 231845
rect 225045 231840 225295 231842
rect 225045 231784 225050 231840
rect 225106 231784 225234 231840
rect 225290 231784 225295 231840
rect 225045 231782 225295 231784
rect 225045 231779 225111 231782
rect 225229 231779 225295 231782
rect 265157 231842 265223 231845
rect 265341 231842 265407 231845
rect 265157 231840 265407 231842
rect 265157 231784 265162 231840
rect 265218 231784 265346 231840
rect 265402 231784 265407 231840
rect 265157 231782 265407 231784
rect 265157 231779 265223 231782
rect 265341 231779 265407 231782
rect 270493 231842 270559 231845
rect 270677 231842 270743 231845
rect 270493 231840 270743 231842
rect 270493 231784 270498 231840
rect 270554 231784 270682 231840
rect 270738 231784 270743 231840
rect 270493 231782 270743 231784
rect 270493 231779 270559 231782
rect 270677 231779 270743 231782
rect 378869 230754 378935 230757
rect 378869 230752 379346 230754
rect 378869 230696 378874 230752
rect 378930 230696 379346 230752
rect 378869 230694 379346 230696
rect 378869 230691 378935 230694
rect 379286 230485 379346 230694
rect 219525 230482 219591 230485
rect 219709 230482 219775 230485
rect 219525 230480 219775 230482
rect 219525 230424 219530 230480
rect 219586 230424 219714 230480
rect 219770 230424 219775 230480
rect 219525 230422 219775 230424
rect 219525 230419 219591 230422
rect 219709 230419 219775 230422
rect 247953 230482 248019 230485
rect 248137 230482 248203 230485
rect 247953 230480 248203 230482
rect 247953 230424 247958 230480
rect 248014 230424 248142 230480
rect 248198 230424 248203 230480
rect 247953 230422 248203 230424
rect 247953 230419 248019 230422
rect 248137 230419 248203 230422
rect 379237 230480 379346 230485
rect 379237 230424 379242 230480
rect 379298 230424 379346 230480
rect 379237 230422 379346 230424
rect 384665 230482 384731 230485
rect 384849 230482 384915 230485
rect 384665 230480 384915 230482
rect 384665 230424 384670 230480
rect 384726 230424 384854 230480
rect 384910 230424 384915 230480
rect 384665 230422 384915 230424
rect 379237 230419 379303 230422
rect 384665 230419 384731 230422
rect 384849 230419 384915 230422
rect 218421 229122 218487 229125
rect 218973 229122 219039 229125
rect 218421 229120 219039 229122
rect 218421 229064 218426 229120
rect 218482 229064 218978 229120
rect 219034 229064 219039 229120
rect 218421 229062 219039 229064
rect 218421 229059 218487 229062
rect 218973 229059 219039 229062
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3325 222594 3391 222597
rect -960 222592 3391 222594
rect -960 222536 3330 222592
rect 3386 222536 3391 222592
rect -960 222534 3391 222536
rect -960 222444 480 222534
rect 3325 222531 3391 222534
rect 153142 222260 153148 222324
rect 153212 222260 153218 222324
rect 153150 222050 153210 222260
rect 190729 222186 190795 222189
rect 190913 222186 190979 222189
rect 190729 222184 190979 222186
rect 190729 222128 190734 222184
rect 190790 222128 190918 222184
rect 190974 222128 190979 222184
rect 190729 222126 190979 222128
rect 190729 222123 190795 222126
rect 190913 222123 190979 222126
rect 191741 222186 191807 222189
rect 191925 222186 191991 222189
rect 191741 222184 191991 222186
rect 191741 222128 191746 222184
rect 191802 222128 191930 222184
rect 191986 222128 191991 222184
rect 191741 222126 191991 222128
rect 191741 222123 191807 222126
rect 191925 222123 191991 222126
rect 153326 222050 153332 222052
rect 153150 221990 153332 222050
rect 153326 221988 153332 221990
rect 153396 221988 153402 222052
rect 151721 221098 151787 221101
rect 151494 221096 151787 221098
rect 151494 221040 151726 221096
rect 151782 221040 151787 221096
rect 151494 221038 151787 221040
rect 151494 220964 151554 221038
rect 151721 221035 151787 221038
rect 151486 220900 151492 220964
rect 151556 220900 151562 220964
rect 153377 220826 153443 220829
rect 153561 220826 153627 220829
rect 153377 220824 153627 220826
rect 153377 220768 153382 220824
rect 153438 220768 153566 220824
rect 153622 220768 153627 220824
rect 153377 220766 153627 220768
rect 153377 220763 153443 220766
rect 153561 220763 153627 220766
rect 206921 220826 206987 220829
rect 207105 220826 207171 220829
rect 206921 220824 207171 220826
rect 206921 220768 206926 220824
rect 206982 220768 207110 220824
rect 207166 220768 207171 220824
rect 206921 220766 207171 220768
rect 206921 220763 206987 220766
rect 207105 220763 207171 220766
rect 225137 220826 225203 220829
rect 225321 220826 225387 220829
rect 225137 220824 225387 220826
rect 225137 220768 225142 220824
rect 225198 220768 225326 220824
rect 225382 220768 225387 220824
rect 225137 220766 225387 220768
rect 225137 220763 225203 220766
rect 225321 220763 225387 220766
rect 238477 220826 238543 220829
rect 238661 220826 238727 220829
rect 238477 220824 238727 220826
rect 238477 220768 238482 220824
rect 238538 220768 238666 220824
rect 238722 220768 238727 220824
rect 238477 220766 238727 220768
rect 238477 220763 238543 220766
rect 238661 220763 238727 220766
rect 374269 220826 374335 220829
rect 374453 220826 374519 220829
rect 374269 220824 374519 220826
rect 374269 220768 374274 220824
rect 374330 220768 374458 220824
rect 374514 220768 374519 220824
rect 374269 220766 374519 220768
rect 374269 220763 374335 220766
rect 374453 220763 374519 220766
rect 580533 217018 580599 217021
rect 583520 217018 584960 217108
rect 580533 217016 584960 217018
rect 580533 216960 580538 217016
rect 580594 216960 584960 217016
rect 580533 216958 584960 216960
rect 580533 216955 580599 216958
rect 583520 216868 584960 216958
rect 152733 215252 152799 215253
rect 152733 215250 152780 215252
rect 152688 215248 152780 215250
rect 152688 215192 152738 215248
rect 152688 215190 152780 215192
rect 152733 215188 152780 215190
rect 152844 215188 152850 215252
rect 152733 215187 152799 215188
rect 152774 215052 152780 215116
rect 152844 215114 152850 215116
rect 153142 215114 153148 215116
rect 152844 215054 153148 215114
rect 152844 215052 152850 215054
rect 153142 215052 153148 215054
rect 153212 215052 153218 215116
rect 151486 212468 151492 212532
rect 151556 212468 151562 212532
rect 190453 212530 190519 212533
rect 190729 212530 190795 212533
rect 190453 212528 190795 212530
rect 190453 212472 190458 212528
rect 190514 212472 190734 212528
rect 190790 212472 190795 212528
rect 190453 212470 190795 212472
rect 151302 212332 151308 212396
rect 151372 212394 151378 212396
rect 151494 212394 151554 212468
rect 190453 212467 190519 212470
rect 190729 212467 190795 212470
rect 424593 212530 424659 212533
rect 424777 212530 424843 212533
rect 424593 212528 424843 212530
rect 424593 212472 424598 212528
rect 424654 212472 424782 212528
rect 424838 212472 424843 212528
rect 424593 212470 424843 212472
rect 424593 212467 424659 212470
rect 424777 212467 424843 212470
rect 151372 212334 151554 212394
rect 151372 212332 151378 212334
rect 198181 211170 198247 211173
rect 198365 211170 198431 211173
rect 198181 211168 198431 211170
rect 198181 211112 198186 211168
rect 198242 211112 198370 211168
rect 198426 211112 198431 211168
rect 198181 211110 198431 211112
rect 198181 211107 198247 211110
rect 198365 211107 198431 211110
rect 206921 211170 206987 211173
rect 207105 211170 207171 211173
rect 206921 211168 207171 211170
rect 206921 211112 206926 211168
rect 206982 211112 207110 211168
rect 207166 211112 207171 211168
rect 206921 211110 207171 211112
rect 206921 211107 206987 211110
rect 207105 211107 207171 211110
rect 219525 211170 219591 211173
rect 219709 211170 219775 211173
rect 219525 211168 219775 211170
rect 219525 211112 219530 211168
rect 219586 211112 219714 211168
rect 219770 211112 219775 211168
rect 219525 211110 219775 211112
rect 219525 211107 219591 211110
rect 219709 211107 219775 211110
rect 223757 211170 223823 211173
rect 223941 211170 224007 211173
rect 223757 211168 224007 211170
rect 223757 211112 223762 211168
rect 223818 211112 223946 211168
rect 224002 211112 224007 211168
rect 223757 211110 224007 211112
rect 223757 211107 223823 211110
rect 223941 211107 224007 211110
rect 238477 211170 238543 211173
rect 238661 211170 238727 211173
rect 238477 211168 238727 211170
rect 238477 211112 238482 211168
rect 238538 211112 238666 211168
rect 238722 211112 238727 211168
rect 238477 211110 238727 211112
rect 238477 211107 238543 211110
rect 238661 211107 238727 211110
rect 374269 211170 374335 211173
rect 374453 211170 374519 211173
rect 374269 211168 374519 211170
rect 374269 211112 374274 211168
rect 374330 211112 374458 211168
rect 374514 211112 374519 211168
rect 374269 211110 374519 211112
rect 374269 211107 374335 211110
rect 374453 211107 374519 211110
rect 152733 208314 152799 208317
rect 614 208312 152799 208314
rect -960 208178 480 208268
rect 614 208256 152738 208312
rect 152794 208256 152799 208312
rect 614 208254 152799 208256
rect 614 208178 674 208254
rect 152733 208251 152799 208254
rect -960 208118 674 208178
rect -960 208028 480 208118
rect 151302 206212 151308 206276
rect 151372 206274 151378 206276
rect 151629 206274 151695 206277
rect 151372 206272 151695 206274
rect 151372 206216 151634 206272
rect 151690 206216 151695 206272
rect 151372 206214 151695 206216
rect 151372 206212 151378 206214
rect 151629 206211 151695 206214
rect 580809 205322 580875 205325
rect 583520 205322 584960 205412
rect 580809 205320 584960 205322
rect 580809 205264 580814 205320
rect 580870 205264 584960 205320
rect 580809 205262 584960 205264
rect 580809 205259 580875 205262
rect 583520 205172 584960 205262
rect 192017 203010 192083 203013
rect 191974 203008 192083 203010
rect 191974 202952 192022 203008
rect 192078 202952 192083 203008
rect 191974 202947 192083 202952
rect 168557 202874 168623 202877
rect 168833 202874 168899 202877
rect 168557 202872 168899 202874
rect 168557 202816 168562 202872
rect 168618 202816 168838 202872
rect 168894 202816 168899 202872
rect 168557 202814 168899 202816
rect 168557 202811 168623 202814
rect 168833 202811 168899 202814
rect 169753 202874 169819 202877
rect 169937 202874 170003 202877
rect 169753 202872 170003 202874
rect 169753 202816 169758 202872
rect 169814 202816 169942 202872
rect 169998 202816 170003 202872
rect 169753 202814 170003 202816
rect 169753 202811 169819 202814
rect 169937 202811 170003 202814
rect 178217 202874 178283 202877
rect 178401 202874 178467 202877
rect 178217 202872 178467 202874
rect 178217 202816 178222 202872
rect 178278 202816 178406 202872
rect 178462 202816 178467 202872
rect 178217 202814 178467 202816
rect 178217 202811 178283 202814
rect 178401 202811 178467 202814
rect 190453 202874 190519 202877
rect 190637 202874 190703 202877
rect 190453 202872 190703 202874
rect 190453 202816 190458 202872
rect 190514 202816 190642 202872
rect 190698 202816 190703 202872
rect 190453 202814 190703 202816
rect 190453 202811 190519 202814
rect 190637 202811 190703 202814
rect 191833 202874 191899 202877
rect 191974 202874 192034 202947
rect 191833 202872 192034 202874
rect 191833 202816 191838 202872
rect 191894 202816 192034 202872
rect 191833 202814 192034 202816
rect 245837 202874 245903 202877
rect 246113 202874 246179 202877
rect 245837 202872 246179 202874
rect 245837 202816 245842 202872
rect 245898 202816 246118 202872
rect 246174 202816 246179 202872
rect 245837 202814 246179 202816
rect 191833 202811 191899 202814
rect 245837 202811 245903 202814
rect 246113 202811 246179 202814
rect 247033 202874 247099 202877
rect 247217 202874 247283 202877
rect 247033 202872 247283 202874
rect 247033 202816 247038 202872
rect 247094 202816 247222 202872
rect 247278 202816 247283 202872
rect 247033 202814 247283 202816
rect 247033 202811 247099 202814
rect 247217 202811 247283 202814
rect 258073 202874 258139 202877
rect 258257 202874 258323 202877
rect 258073 202872 258323 202874
rect 258073 202816 258078 202872
rect 258134 202816 258262 202872
rect 258318 202816 258323 202872
rect 258073 202814 258323 202816
rect 258073 202811 258139 202814
rect 258257 202811 258323 202814
rect 263593 202874 263659 202877
rect 263777 202874 263843 202877
rect 263593 202872 263843 202874
rect 263593 202816 263598 202872
rect 263654 202816 263782 202872
rect 263838 202816 263843 202872
rect 263593 202814 263843 202816
rect 263593 202811 263659 202814
rect 263777 202811 263843 202814
rect 271873 202874 271939 202877
rect 272057 202874 272123 202877
rect 271873 202872 272123 202874
rect 271873 202816 271878 202872
rect 271934 202816 272062 202872
rect 272118 202816 272123 202872
rect 271873 202814 272123 202816
rect 271873 202811 271939 202814
rect 272057 202811 272123 202814
rect 403709 202874 403775 202877
rect 403985 202874 404051 202877
rect 403709 202872 404051 202874
rect 403709 202816 403714 202872
rect 403770 202816 403990 202872
rect 404046 202816 404051 202872
rect 403709 202814 404051 202816
rect 403709 202811 403775 202814
rect 403985 202811 404051 202814
rect 424501 202874 424567 202877
rect 424685 202874 424751 202877
rect 424501 202872 424751 202874
rect 424501 202816 424506 202872
rect 424562 202816 424690 202872
rect 424746 202816 424751 202872
rect 424501 202814 424751 202816
rect 424501 202811 424567 202814
rect 424685 202811 424751 202814
rect 205909 201514 205975 201517
rect 206093 201514 206159 201517
rect 205909 201512 206159 201514
rect 205909 201456 205914 201512
rect 205970 201456 206098 201512
rect 206154 201456 206159 201512
rect 205909 201454 206159 201456
rect 205909 201451 205975 201454
rect 206093 201451 206159 201454
rect 238477 201514 238543 201517
rect 238661 201514 238727 201517
rect 238477 201512 238727 201514
rect 238477 201456 238482 201512
rect 238538 201456 238666 201512
rect 238722 201456 238727 201512
rect 238477 201454 238727 201456
rect 238477 201451 238543 201454
rect 238661 201451 238727 201454
rect 379053 201514 379119 201517
rect 379237 201514 379303 201517
rect 379053 201512 379303 201514
rect 379053 201456 379058 201512
rect 379114 201456 379242 201512
rect 379298 201456 379303 201512
rect 379053 201454 379303 201456
rect 379053 201451 379119 201454
rect 379237 201451 379303 201454
rect 151854 201316 151860 201380
rect 151924 201378 151930 201380
rect 151997 201378 152063 201381
rect 151924 201376 152063 201378
rect 151924 201320 152002 201376
rect 152058 201320 152063 201376
rect 151924 201318 152063 201320
rect 151924 201316 151930 201318
rect 151997 201315 152063 201318
rect 194501 198794 194567 198797
rect 195973 198794 196039 198797
rect 194501 198792 194610 198794
rect 194501 198736 194506 198792
rect 194562 198736 194610 198792
rect 194501 198731 194610 198736
rect 195973 198792 196082 198794
rect 195973 198736 195978 198792
rect 196034 198736 196082 198792
rect 195973 198731 196082 198736
rect 194550 198522 194610 198731
rect 194777 198522 194843 198525
rect 194550 198520 194843 198522
rect 194550 198464 194782 198520
rect 194838 198464 194843 198520
rect 194550 198462 194843 198464
rect 196022 198522 196082 198731
rect 196341 198522 196407 198525
rect 196022 198520 196407 198522
rect 196022 198464 196346 198520
rect 196402 198464 196407 198520
rect 196022 198462 196407 198464
rect 194777 198459 194843 198462
rect 196341 198459 196407 198462
rect 151854 196556 151860 196620
rect 151924 196618 151930 196620
rect 151997 196618 152063 196621
rect 151924 196616 152063 196618
rect 151924 196560 152002 196616
rect 152058 196560 152063 196616
rect 151924 196558 152063 196560
rect 151924 196556 151930 196558
rect 151997 196555 152063 196558
rect -960 193898 480 193988
rect 2773 193898 2839 193901
rect -960 193896 2839 193898
rect -960 193840 2778 193896
rect 2834 193840 2839 193896
rect -960 193838 2839 193840
rect -960 193748 480 193838
rect 2773 193835 2839 193838
rect 583520 193476 584960 193716
rect 151629 193220 151695 193221
rect 151629 193218 151676 193220
rect 151584 193216 151676 193218
rect 151584 193160 151634 193216
rect 151584 193158 151676 193160
rect 151629 193156 151676 193158
rect 151740 193156 151746 193220
rect 151813 193218 151879 193221
rect 151997 193218 152063 193221
rect 151813 193216 152063 193218
rect 151813 193160 151818 193216
rect 151874 193160 152002 193216
rect 152058 193160 152063 193216
rect 151813 193158 152063 193160
rect 151629 193155 151695 193156
rect 151813 193155 151879 193158
rect 151997 193155 152063 193158
rect 190729 193218 190795 193221
rect 190913 193218 190979 193221
rect 190729 193216 190979 193218
rect 190729 193160 190734 193216
rect 190790 193160 190918 193216
rect 190974 193160 190979 193216
rect 190729 193158 190979 193160
rect 190729 193155 190795 193158
rect 190913 193155 190979 193158
rect 192017 193218 192083 193221
rect 192201 193218 192267 193221
rect 192017 193216 192267 193218
rect 192017 193160 192022 193216
rect 192078 193160 192206 193216
rect 192262 193160 192267 193216
rect 192017 193158 192267 193160
rect 192017 193155 192083 193158
rect 192201 193155 192267 193158
rect 234797 193218 234863 193221
rect 234981 193218 235047 193221
rect 234797 193216 235047 193218
rect 234797 193160 234802 193216
rect 234858 193160 234986 193216
rect 235042 193160 235047 193216
rect 234797 193158 235047 193160
rect 234797 193155 234863 193158
rect 234981 193155 235047 193158
rect 239029 193218 239095 193221
rect 239213 193218 239279 193221
rect 239029 193216 239279 193218
rect 239029 193160 239034 193216
rect 239090 193160 239218 193216
rect 239274 193160 239279 193216
rect 239029 193158 239279 193160
rect 239029 193155 239095 193158
rect 239213 193155 239279 193158
rect 424593 193218 424659 193221
rect 424777 193218 424843 193221
rect 424593 193216 424843 193218
rect 424593 193160 424598 193216
rect 424654 193160 424782 193216
rect 424838 193160 424843 193216
rect 424593 193158 424843 193160
rect 424593 193155 424659 193158
rect 424777 193155 424843 193158
rect 208393 191858 208459 191861
rect 208577 191858 208643 191861
rect 208393 191856 208643 191858
rect 208393 191800 208398 191856
rect 208454 191800 208582 191856
rect 208638 191800 208643 191856
rect 208393 191798 208643 191800
rect 208393 191795 208459 191798
rect 208577 191795 208643 191798
rect 374269 191858 374335 191861
rect 374453 191858 374519 191861
rect 374269 191856 374519 191858
rect 374269 191800 374274 191856
rect 374330 191800 374458 191856
rect 374514 191800 374519 191856
rect 374269 191798 374519 191800
rect 374269 191795 374335 191798
rect 374453 191795 374519 191798
rect 226701 190634 226767 190637
rect 226382 190632 226767 190634
rect 226382 190576 226706 190632
rect 226762 190576 226767 190632
rect 226382 190574 226767 190576
rect 226382 190501 226442 190574
rect 226701 190571 226767 190574
rect 226382 190496 226491 190501
rect 226382 190440 226430 190496
rect 226486 190440 226491 190496
rect 226382 190438 226491 190440
rect 226425 190435 226491 190438
rect 154757 183562 154823 183565
rect 154941 183562 155007 183565
rect 154757 183560 155007 183562
rect 154757 183504 154762 183560
rect 154818 183504 154946 183560
rect 155002 183504 155007 183560
rect 154757 183502 155007 183504
rect 154757 183499 154823 183502
rect 154941 183499 155007 183502
rect 168557 183562 168623 183565
rect 168833 183562 168899 183565
rect 168557 183560 168899 183562
rect 168557 183504 168562 183560
rect 168618 183504 168838 183560
rect 168894 183504 168899 183560
rect 168557 183502 168899 183504
rect 168557 183499 168623 183502
rect 168833 183499 168899 183502
rect 169753 183562 169819 183565
rect 169937 183562 170003 183565
rect 169753 183560 170003 183562
rect 169753 183504 169758 183560
rect 169814 183504 169942 183560
rect 169998 183504 170003 183560
rect 169753 183502 170003 183504
rect 169753 183499 169819 183502
rect 169937 183499 170003 183502
rect 173985 183562 174051 183565
rect 174261 183562 174327 183565
rect 173985 183560 174327 183562
rect 173985 183504 173990 183560
rect 174046 183504 174266 183560
rect 174322 183504 174327 183560
rect 173985 183502 174327 183504
rect 173985 183499 174051 183502
rect 174261 183499 174327 183502
rect 178217 183562 178283 183565
rect 178401 183562 178467 183565
rect 178217 183560 178467 183562
rect 178217 183504 178222 183560
rect 178278 183504 178406 183560
rect 178462 183504 178467 183560
rect 178217 183502 178467 183504
rect 178217 183499 178283 183502
rect 178401 183499 178467 183502
rect 216581 183562 216647 183565
rect 216765 183562 216831 183565
rect 216581 183560 216831 183562
rect 216581 183504 216586 183560
rect 216642 183504 216770 183560
rect 216826 183504 216831 183560
rect 216581 183502 216831 183504
rect 216581 183499 216647 183502
rect 216765 183499 216831 183502
rect 245837 183562 245903 183565
rect 246113 183562 246179 183565
rect 245837 183560 246179 183562
rect 245837 183504 245842 183560
rect 245898 183504 246118 183560
rect 246174 183504 246179 183560
rect 245837 183502 246179 183504
rect 245837 183499 245903 183502
rect 246113 183499 246179 183502
rect 247033 183562 247099 183565
rect 247217 183562 247283 183565
rect 247033 183560 247283 183562
rect 247033 183504 247038 183560
rect 247094 183504 247222 183560
rect 247278 183504 247283 183560
rect 247033 183502 247283 183504
rect 247033 183499 247099 183502
rect 247217 183499 247283 183502
rect 252553 183562 252619 183565
rect 252737 183562 252803 183565
rect 252553 183560 252803 183562
rect 252553 183504 252558 183560
rect 252614 183504 252742 183560
rect 252798 183504 252803 183560
rect 252553 183502 252803 183504
rect 252553 183499 252619 183502
rect 252737 183499 252803 183502
rect 258073 183562 258139 183565
rect 258257 183562 258323 183565
rect 258073 183560 258323 183562
rect 258073 183504 258078 183560
rect 258134 183504 258262 183560
rect 258318 183504 258323 183560
rect 258073 183502 258323 183504
rect 258073 183499 258139 183502
rect 258257 183499 258323 183502
rect 263593 183562 263659 183565
rect 263777 183562 263843 183565
rect 263593 183560 263843 183562
rect 263593 183504 263598 183560
rect 263654 183504 263782 183560
rect 263838 183504 263843 183560
rect 263593 183502 263843 183504
rect 263593 183499 263659 183502
rect 263777 183499 263843 183502
rect 271873 183562 271939 183565
rect 272057 183562 272123 183565
rect 271873 183560 272123 183562
rect 271873 183504 271878 183560
rect 271934 183504 272062 183560
rect 272118 183504 272123 183560
rect 271873 183502 272123 183504
rect 271873 183499 271939 183502
rect 272057 183499 272123 183502
rect 284385 183562 284451 183565
rect 284661 183562 284727 183565
rect 284385 183560 284727 183562
rect 284385 183504 284390 183560
rect 284446 183504 284666 183560
rect 284722 183504 284727 183560
rect 284385 183502 284727 183504
rect 284385 183499 284451 183502
rect 284661 183499 284727 183502
rect 307937 183562 308003 183565
rect 308213 183562 308279 183565
rect 307937 183560 308279 183562
rect 307937 183504 307942 183560
rect 307998 183504 308218 183560
rect 308274 183504 308279 183560
rect 307937 183502 308279 183504
rect 307937 183499 308003 183502
rect 308213 183499 308279 183502
rect 346025 183562 346091 183565
rect 346209 183562 346275 183565
rect 346025 183560 346275 183562
rect 346025 183504 346030 183560
rect 346086 183504 346214 183560
rect 346270 183504 346275 183560
rect 346025 183502 346275 183504
rect 346025 183499 346091 183502
rect 346209 183499 346275 183502
rect 357065 183562 357131 183565
rect 357249 183562 357315 183565
rect 357065 183560 357315 183562
rect 357065 183504 357070 183560
rect 357126 183504 357254 183560
rect 357310 183504 357315 183560
rect 357065 183502 357315 183504
rect 357065 183499 357131 183502
rect 357249 183499 357315 183502
rect 403709 183562 403775 183565
rect 403985 183562 404051 183565
rect 403709 183560 404051 183562
rect 403709 183504 403714 183560
rect 403770 183504 403990 183560
rect 404046 183504 404051 183560
rect 403709 183502 404051 183504
rect 403709 183499 403775 183502
rect 403985 183499 404051 183502
rect 424501 183562 424567 183565
rect 424685 183562 424751 183565
rect 424501 183560 424751 183562
rect 424501 183504 424506 183560
rect 424562 183504 424690 183560
rect 424746 183504 424751 183560
rect 424501 183502 424751 183504
rect 424501 183499 424567 183502
rect 424685 183499 424751 183502
rect 223849 182202 223915 182205
rect 224033 182202 224099 182205
rect 223849 182200 224099 182202
rect 223849 182144 223854 182200
rect 223910 182144 224038 182200
rect 224094 182144 224099 182200
rect 223849 182142 224099 182144
rect 223849 182139 223915 182142
rect 224033 182139 224099 182142
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect 226609 180842 226675 180845
rect 226793 180842 226859 180845
rect 226609 180840 226859 180842
rect 226609 180784 226614 180840
rect 226670 180784 226798 180840
rect 226854 180784 226859 180840
rect 226609 180782 226859 180784
rect 226609 180779 226675 180782
rect 226793 180779 226859 180782
rect -960 179482 480 179572
rect 2773 179482 2839 179485
rect -960 179480 2839 179482
rect -960 179424 2778 179480
rect 2834 179424 2839 179480
rect -960 179422 2839 179424
rect -960 179332 480 179422
rect 2773 179419 2839 179422
rect 151302 177244 151308 177308
rect 151372 177306 151378 177308
rect 151445 177306 151511 177309
rect 151372 177304 151511 177306
rect 151372 177248 151450 177304
rect 151506 177248 151511 177304
rect 151372 177246 151511 177248
rect 151372 177244 151378 177246
rect 151445 177243 151511 177246
rect 154849 173906 154915 173909
rect 155033 173906 155099 173909
rect 154849 173904 155099 173906
rect 154849 173848 154854 173904
rect 154910 173848 155038 173904
rect 155094 173848 155099 173904
rect 154849 173846 155099 173848
rect 154849 173843 154915 173846
rect 155033 173843 155099 173846
rect 248137 172546 248203 172549
rect 248321 172546 248387 172549
rect 248137 172544 248387 172546
rect 248137 172488 248142 172544
rect 248198 172488 248326 172544
rect 248382 172488 248387 172544
rect 248137 172486 248387 172488
rect 248137 172483 248203 172486
rect 248321 172483 248387 172486
rect 374269 172546 374335 172549
rect 374453 172546 374519 172549
rect 374269 172544 374519 172546
rect 374269 172488 374274 172544
rect 374330 172488 374458 172544
rect 374514 172488 374519 172544
rect 374269 172486 374519 172488
rect 374269 172483 374335 172486
rect 374453 172483 374519 172486
rect 580441 170098 580507 170101
rect 583520 170098 584960 170188
rect 580441 170096 584960 170098
rect 580441 170040 580446 170096
rect 580502 170040 584960 170096
rect 580441 170038 584960 170040
rect 580441 170035 580507 170038
rect 583520 169948 584960 170038
rect 151854 165610 151860 165612
rect 614 165550 151860 165610
rect -960 165066 480 165156
rect 614 165066 674 165550
rect 151854 165548 151860 165550
rect 151924 165548 151930 165612
rect 151118 165412 151124 165476
rect 151188 165474 151194 165476
rect 151445 165474 151511 165477
rect 151188 165472 151511 165474
rect 151188 165416 151450 165472
rect 151506 165416 151511 165472
rect 151188 165414 151511 165416
rect 151188 165412 151194 165414
rect 151445 165411 151511 165414
rect -960 165006 674 165066
rect -960 164916 480 165006
rect 150709 164386 150775 164389
rect 150709 164384 150818 164386
rect 150709 164328 150714 164384
rect 150770 164328 150818 164384
rect 150709 164323 150818 164328
rect 150758 164253 150818 164323
rect 150758 164248 150867 164253
rect 150758 164192 150806 164248
rect 150862 164192 150867 164248
rect 150758 164190 150867 164192
rect 150801 164187 150867 164190
rect 154849 164250 154915 164253
rect 155033 164250 155099 164253
rect 154849 164248 155099 164250
rect 154849 164192 154854 164248
rect 154910 164192 155038 164248
rect 155094 164192 155099 164248
rect 154849 164190 155099 164192
rect 154849 164187 154915 164190
rect 155033 164187 155099 164190
rect 216857 163026 216923 163029
rect 218329 163026 218395 163029
rect 216814 163024 216923 163026
rect 216814 162968 216862 163024
rect 216918 162968 216923 163024
rect 216814 162963 216923 162968
rect 218286 163024 218395 163026
rect 218286 162968 218334 163024
rect 218390 162968 218395 163024
rect 218286 162963 218395 162968
rect 216814 162893 216874 162963
rect 218286 162893 218346 162963
rect 192017 162890 192083 162893
rect 191974 162888 192083 162890
rect 191974 162832 192022 162888
rect 192078 162832 192083 162888
rect 191974 162827 192083 162832
rect 216765 162888 216874 162893
rect 216765 162832 216770 162888
rect 216826 162832 216874 162888
rect 216765 162830 216874 162832
rect 218237 162888 218346 162893
rect 218237 162832 218242 162888
rect 218298 162832 218346 162888
rect 218237 162830 218346 162832
rect 234797 162890 234863 162893
rect 234981 162890 235047 162893
rect 234797 162888 235047 162890
rect 234797 162832 234802 162888
rect 234858 162832 234986 162888
rect 235042 162832 235047 162888
rect 234797 162830 235047 162832
rect 216765 162827 216831 162830
rect 218237 162827 218303 162830
rect 234797 162827 234863 162830
rect 234981 162827 235047 162830
rect 424777 162890 424843 162893
rect 424961 162890 425027 162893
rect 424777 162888 425027 162890
rect 424777 162832 424782 162888
rect 424838 162832 424966 162888
rect 425022 162832 425027 162888
rect 424777 162830 425027 162832
rect 424777 162827 424843 162830
rect 424961 162827 425027 162830
rect 191974 162754 192034 162827
rect 192109 162754 192175 162757
rect 191974 162752 192175 162754
rect 191974 162696 192114 162752
rect 192170 162696 192175 162752
rect 191974 162694 192175 162696
rect 192109 162691 192175 162694
rect 580073 158402 580139 158405
rect 583520 158402 584960 158492
rect 580073 158400 584960 158402
rect 580073 158344 580078 158400
rect 580134 158344 584960 158400
rect 580073 158342 584960 158344
rect 580073 158339 580139 158342
rect 583520 158252 584960 158342
rect 151118 156572 151124 156636
rect 151188 156634 151194 156636
rect 151486 156634 151492 156636
rect 151188 156574 151492 156634
rect 151188 156572 151194 156574
rect 151486 156572 151492 156574
rect 151556 156572 151562 156636
rect 226517 154730 226583 154733
rect 226517 154728 226626 154730
rect 226517 154672 226522 154728
rect 226578 154672 226626 154728
rect 226517 154667 226626 154672
rect 226566 154597 226626 154667
rect 178217 154594 178283 154597
rect 178401 154594 178467 154597
rect 178217 154592 178467 154594
rect 178217 154536 178222 154592
rect 178278 154536 178406 154592
rect 178462 154536 178467 154592
rect 178217 154534 178467 154536
rect 178217 154531 178283 154534
rect 178401 154531 178467 154534
rect 226517 154592 226626 154597
rect 226517 154536 226522 154592
rect 226578 154536 226626 154592
rect 226517 154534 226626 154536
rect 247033 154594 247099 154597
rect 247309 154594 247375 154597
rect 247033 154592 247375 154594
rect 247033 154536 247038 154592
rect 247094 154536 247314 154592
rect 247370 154536 247375 154592
rect 247033 154534 247375 154536
rect 226517 154531 226583 154534
rect 247033 154531 247099 154534
rect 247309 154531 247375 154534
rect 258073 154594 258139 154597
rect 258349 154594 258415 154597
rect 258073 154592 258415 154594
rect 258073 154536 258078 154592
rect 258134 154536 258354 154592
rect 258410 154536 258415 154592
rect 258073 154534 258415 154536
rect 258073 154531 258139 154534
rect 258349 154531 258415 154534
rect 403525 154594 403591 154597
rect 403801 154594 403867 154597
rect 403525 154592 403867 154594
rect 403525 154536 403530 154592
rect 403586 154536 403806 154592
rect 403862 154536 403867 154592
rect 403525 154534 403867 154536
rect 403525 154531 403591 154534
rect 403801 154531 403867 154534
rect 190453 153234 190519 153237
rect 190729 153234 190795 153237
rect 190453 153232 190795 153234
rect 190453 153176 190458 153232
rect 190514 153176 190734 153232
rect 190790 153176 190795 153232
rect 190453 153174 190795 153176
rect 190453 153171 190519 153174
rect 190729 153171 190795 153174
rect 238385 153234 238451 153237
rect 238569 153234 238635 153237
rect 238385 153232 238635 153234
rect 238385 153176 238390 153232
rect 238446 153176 238574 153232
rect 238630 153176 238635 153232
rect 238385 153174 238635 153176
rect 238385 153171 238451 153174
rect 238569 153171 238635 153174
rect 217961 151874 218027 151877
rect 217961 151872 218162 151874
rect 217961 151816 217966 151872
rect 218022 151816 218162 151872
rect 217961 151814 218162 151816
rect 217961 151811 218027 151814
rect 217961 151738 218027 151741
rect 218102 151738 218162 151814
rect 217961 151736 218162 151738
rect 217961 151680 217966 151736
rect 218022 151680 218162 151736
rect 217961 151678 218162 151680
rect 217961 151675 218027 151678
rect -960 150786 480 150876
rect 3325 150786 3391 150789
rect -960 150784 3391 150786
rect -960 150728 3330 150784
rect 3386 150728 3391 150784
rect -960 150726 3391 150728
rect -960 150636 480 150726
rect 3325 150723 3391 150726
rect 151486 147794 151492 147796
rect 151310 147734 151492 147794
rect 151310 147524 151370 147734
rect 151486 147732 151492 147734
rect 151556 147732 151562 147796
rect 151302 147460 151308 147524
rect 151372 147460 151378 147524
rect 583520 146556 584960 146796
rect 189257 145074 189323 145077
rect 189257 145072 189458 145074
rect 189257 145016 189262 145072
rect 189318 145016 189458 145072
rect 189257 145014 189458 145016
rect 189257 145011 189323 145014
rect 189257 144938 189323 144941
rect 189398 144938 189458 145014
rect 189257 144936 189458 144938
rect 189257 144880 189262 144936
rect 189318 144880 189458 144936
rect 189257 144878 189458 144880
rect 191925 144938 191991 144941
rect 192109 144938 192175 144941
rect 191925 144936 192175 144938
rect 191925 144880 191930 144936
rect 191986 144880 192114 144936
rect 192170 144880 192175 144936
rect 191925 144878 192175 144880
rect 189257 144875 189323 144878
rect 191925 144875 191991 144878
rect 192109 144875 192175 144878
rect 265065 144938 265131 144941
rect 265249 144938 265315 144941
rect 265065 144936 265315 144938
rect 265065 144880 265070 144936
rect 265126 144880 265254 144936
rect 265310 144880 265315 144936
rect 265065 144878 265315 144880
rect 265065 144875 265131 144878
rect 265249 144875 265315 144878
rect 270493 144938 270559 144941
rect 270769 144938 270835 144941
rect 270493 144936 270835 144938
rect 270493 144880 270498 144936
rect 270554 144880 270774 144936
rect 270830 144880 270835 144936
rect 270493 144878 270835 144880
rect 270493 144875 270559 144878
rect 270769 144875 270835 144878
rect 271873 144938 271939 144941
rect 272057 144938 272123 144941
rect 271873 144936 272123 144938
rect 271873 144880 271878 144936
rect 271934 144880 272062 144936
rect 272118 144880 272123 144936
rect 271873 144878 272123 144880
rect 271873 144875 271939 144878
rect 272057 144875 272123 144878
rect 263777 143714 263843 143717
rect 263734 143712 263843 143714
rect 263734 143656 263782 143712
rect 263838 143656 263843 143712
rect 263734 143651 263843 143656
rect 263734 143581 263794 143651
rect 168465 143578 168531 143581
rect 168833 143578 168899 143581
rect 168465 143576 168899 143578
rect 168465 143520 168470 143576
rect 168526 143520 168838 143576
rect 168894 143520 168899 143576
rect 168465 143518 168899 143520
rect 263734 143576 263843 143581
rect 263734 143520 263782 143576
rect 263838 143520 263843 143576
rect 263734 143518 263843 143520
rect 168465 143515 168531 143518
rect 168833 143515 168899 143518
rect 263777 143515 263843 143518
rect 196157 140722 196223 140725
rect 196022 140720 196223 140722
rect 196022 140664 196162 140720
rect 196218 140664 196223 140720
rect 196022 140662 196223 140664
rect 196022 140586 196082 140662
rect 196157 140659 196223 140662
rect 196249 140586 196315 140589
rect 196022 140584 196315 140586
rect 196022 140528 196254 140584
rect 196310 140528 196315 140584
rect 196022 140526 196315 140528
rect 196249 140523 196315 140526
rect -960 136370 480 136460
rect 3877 136370 3943 136373
rect -960 136368 3943 136370
rect -960 136312 3882 136368
rect 3938 136312 3943 136368
rect -960 136310 3943 136312
rect -960 136220 480 136310
rect 3877 136307 3943 136310
rect 169753 135282 169819 135285
rect 170029 135282 170095 135285
rect 169753 135280 170095 135282
rect 169753 135224 169758 135280
rect 169814 135224 170034 135280
rect 170090 135224 170095 135280
rect 169753 135222 170095 135224
rect 169753 135219 169819 135222
rect 170029 135219 170095 135222
rect 178217 135282 178283 135285
rect 178401 135282 178467 135285
rect 178217 135280 178467 135282
rect 178217 135224 178222 135280
rect 178278 135224 178406 135280
rect 178462 135224 178467 135280
rect 178217 135222 178467 135224
rect 178217 135219 178283 135222
rect 178401 135219 178467 135222
rect 191833 135282 191899 135285
rect 192017 135282 192083 135285
rect 191833 135280 192083 135282
rect 191833 135224 191838 135280
rect 191894 135224 192022 135280
rect 192078 135224 192083 135280
rect 191833 135222 192083 135224
rect 191833 135219 191899 135222
rect 192017 135219 192083 135222
rect 207013 135282 207079 135285
rect 207197 135282 207263 135285
rect 207013 135280 207263 135282
rect 207013 135224 207018 135280
rect 207074 135224 207202 135280
rect 207258 135224 207263 135280
rect 207013 135222 207263 135224
rect 207013 135219 207079 135222
rect 207197 135219 207263 135222
rect 222469 135282 222535 135285
rect 222653 135282 222719 135285
rect 222469 135280 222719 135282
rect 222469 135224 222474 135280
rect 222530 135224 222658 135280
rect 222714 135224 222719 135280
rect 222469 135222 222719 135224
rect 222469 135219 222535 135222
rect 222653 135219 222719 135222
rect 223757 135282 223823 135285
rect 223941 135282 224007 135285
rect 223757 135280 224007 135282
rect 223757 135224 223762 135280
rect 223818 135224 223946 135280
rect 224002 135224 224007 135280
rect 223757 135222 224007 135224
rect 223757 135219 223823 135222
rect 223941 135219 224007 135222
rect 226517 135282 226583 135285
rect 226701 135282 226767 135285
rect 226517 135280 226767 135282
rect 226517 135224 226522 135280
rect 226578 135224 226706 135280
rect 226762 135224 226767 135280
rect 226517 135222 226767 135224
rect 226517 135219 226583 135222
rect 226701 135219 226767 135222
rect 229277 135282 229343 135285
rect 229461 135282 229527 135285
rect 229277 135280 229527 135282
rect 229277 135224 229282 135280
rect 229338 135224 229466 135280
rect 229522 135224 229527 135280
rect 229277 135222 229527 135224
rect 229277 135219 229343 135222
rect 229461 135219 229527 135222
rect 234797 135282 234863 135285
rect 234981 135282 235047 135285
rect 234797 135280 235047 135282
rect 234797 135224 234802 135280
rect 234858 135224 234986 135280
rect 235042 135224 235047 135280
rect 234797 135222 235047 135224
rect 234797 135219 234863 135222
rect 234981 135219 235047 135222
rect 258073 135282 258139 135285
rect 258349 135282 258415 135285
rect 258073 135280 258415 135282
rect 258073 135224 258078 135280
rect 258134 135224 258354 135280
rect 258410 135224 258415 135280
rect 258073 135222 258415 135224
rect 258073 135219 258139 135222
rect 258349 135219 258415 135222
rect 265065 135282 265131 135285
rect 265249 135282 265315 135285
rect 265065 135280 265315 135282
rect 265065 135224 265070 135280
rect 265126 135224 265254 135280
rect 265310 135224 265315 135280
rect 265065 135222 265315 135224
rect 265065 135219 265131 135222
rect 265249 135219 265315 135222
rect 384665 135282 384731 135285
rect 384849 135282 384915 135285
rect 384665 135280 384915 135282
rect 384665 135224 384670 135280
rect 384726 135224 384854 135280
rect 384910 135224 384915 135280
rect 384665 135222 384915 135224
rect 384665 135219 384731 135222
rect 384849 135219 384915 135222
rect 580625 134874 580691 134877
rect 583520 134874 584960 134964
rect 580625 134872 584960 134874
rect 580625 134816 580630 134872
rect 580686 134816 584960 134872
rect 580625 134814 584960 134816
rect 580625 134811 580691 134814
rect 583520 134724 584960 134814
rect 153377 133922 153443 133925
rect 153561 133922 153627 133925
rect 153377 133920 153627 133922
rect 153377 133864 153382 133920
rect 153438 133864 153566 133920
rect 153622 133864 153627 133920
rect 153377 133862 153627 133864
rect 153377 133859 153443 133862
rect 153561 133859 153627 133862
rect 156137 133922 156203 133925
rect 156321 133922 156387 133925
rect 156137 133920 156387 133922
rect 156137 133864 156142 133920
rect 156198 133864 156326 133920
rect 156382 133864 156387 133920
rect 156137 133862 156387 133864
rect 156137 133859 156203 133862
rect 156321 133859 156387 133862
rect 190361 133922 190427 133925
rect 190637 133922 190703 133925
rect 190361 133920 190703 133922
rect 190361 133864 190366 133920
rect 190422 133864 190642 133920
rect 190698 133864 190703 133920
rect 190361 133862 190703 133864
rect 190361 133859 190427 133862
rect 190637 133859 190703 133862
rect 189257 125762 189323 125765
rect 189257 125760 189458 125762
rect 189257 125704 189262 125760
rect 189318 125704 189458 125760
rect 189257 125702 189458 125704
rect 189257 125699 189323 125702
rect 189257 125626 189323 125629
rect 189398 125626 189458 125702
rect 189257 125624 189458 125626
rect 189257 125568 189262 125624
rect 189318 125568 189458 125624
rect 189257 125566 189458 125568
rect 271873 125626 271939 125629
rect 272057 125626 272123 125629
rect 271873 125624 272123 125626
rect 271873 125568 271878 125624
rect 271934 125568 272062 125624
rect 272118 125568 272123 125624
rect 271873 125566 272123 125568
rect 189257 125563 189323 125566
rect 271873 125563 271939 125566
rect 272057 125563 272123 125566
rect 403249 125626 403315 125629
rect 403433 125626 403499 125629
rect 403249 125624 403499 125626
rect 403249 125568 403254 125624
rect 403310 125568 403438 125624
rect 403494 125568 403499 125624
rect 403249 125566 403499 125568
rect 403249 125563 403315 125566
rect 403433 125563 403499 125566
rect 190453 124266 190519 124269
rect 190637 124266 190703 124269
rect 190453 124264 190703 124266
rect 190453 124208 190458 124264
rect 190514 124208 190642 124264
rect 190698 124208 190703 124264
rect 190453 124206 190703 124208
rect 190453 124203 190519 124206
rect 190637 124203 190703 124206
rect 423305 124266 423371 124269
rect 423489 124266 423555 124269
rect 423305 124264 423555 124266
rect 423305 124208 423310 124264
rect 423366 124208 423494 124264
rect 423550 124208 423555 124264
rect 423305 124206 423555 124208
rect 423305 124203 423371 124206
rect 423489 124203 423555 124206
rect 580349 123178 580415 123181
rect 583520 123178 584960 123268
rect 580349 123176 584960 123178
rect 580349 123120 580354 123176
rect 580410 123120 584960 123176
rect 580349 123118 584960 123120
rect 580349 123115 580415 123118
rect 583520 123028 584960 123118
rect 2957 122770 3023 122773
rect 152958 122770 152964 122772
rect 2957 122768 152964 122770
rect 2957 122712 2962 122768
rect 3018 122712 152964 122768
rect 2957 122710 152964 122712
rect 2957 122707 3023 122710
rect 152958 122708 152964 122710
rect 153028 122708 153034 122772
rect -960 122090 480 122180
rect 2957 122090 3023 122093
rect -960 122088 3023 122090
rect -960 122032 2962 122088
rect 3018 122032 3023 122088
rect -960 122030 3023 122032
rect -960 121940 480 122030
rect 2957 122027 3023 122030
rect 207105 116106 207171 116109
rect 236361 116106 236427 116109
rect 237649 116106 237715 116109
rect 207062 116104 207171 116106
rect 207062 116048 207110 116104
rect 207166 116048 207171 116104
rect 207062 116043 207171 116048
rect 236318 116104 236427 116106
rect 236318 116048 236366 116104
rect 236422 116048 236427 116104
rect 236318 116043 236427 116048
rect 237606 116104 237715 116106
rect 237606 116048 237654 116104
rect 237710 116048 237715 116104
rect 237606 116043 237715 116048
rect 207062 115973 207122 116043
rect 236318 115973 236378 116043
rect 237606 115973 237666 116043
rect 169753 115970 169819 115973
rect 170029 115970 170095 115973
rect 169753 115968 170095 115970
rect 169753 115912 169758 115968
rect 169814 115912 170034 115968
rect 170090 115912 170095 115968
rect 169753 115910 170095 115912
rect 169753 115907 169819 115910
rect 170029 115907 170095 115910
rect 207013 115968 207122 115973
rect 207013 115912 207018 115968
rect 207074 115912 207122 115968
rect 207013 115910 207122 115912
rect 236269 115968 236378 115973
rect 236269 115912 236274 115968
rect 236330 115912 236378 115968
rect 236269 115910 236378 115912
rect 237557 115968 237666 115973
rect 237557 115912 237562 115968
rect 237618 115912 237666 115968
rect 237557 115910 237666 115912
rect 258073 115970 258139 115973
rect 258349 115970 258415 115973
rect 258073 115968 258415 115970
rect 258073 115912 258078 115968
rect 258134 115912 258354 115968
rect 258410 115912 258415 115968
rect 258073 115910 258415 115912
rect 207013 115907 207079 115910
rect 236269 115907 236335 115910
rect 237557 115907 237623 115910
rect 258073 115907 258139 115910
rect 258349 115907 258415 115910
rect 151302 114684 151308 114748
rect 151372 114746 151378 114748
rect 245745 114746 245811 114749
rect 151372 114686 151554 114746
rect 151372 114684 151378 114686
rect 151494 114612 151554 114686
rect 245745 114744 246130 114746
rect 245745 114688 245750 114744
rect 245806 114688 246130 114744
rect 245745 114686 246130 114688
rect 245745 114683 245811 114686
rect 151486 114548 151492 114612
rect 151556 114548 151562 114612
rect 245929 114610 245995 114613
rect 246070 114610 246130 114686
rect 245929 114608 246130 114610
rect 245929 114552 245934 114608
rect 245990 114552 246130 114608
rect 245929 114550 246130 114552
rect 245929 114547 245995 114550
rect 151486 113052 151492 113116
rect 151556 113052 151562 113116
rect 151494 112981 151554 113052
rect 151494 112976 151603 112981
rect 151494 112920 151542 112976
rect 151598 112920 151603 112976
rect 151494 112918 151603 112920
rect 151537 112915 151603 112918
rect 191741 111754 191807 111757
rect 191925 111754 191991 111757
rect 191741 111752 191991 111754
rect 191741 111696 191746 111752
rect 191802 111696 191930 111752
rect 191986 111696 191991 111752
rect 191741 111694 191991 111696
rect 191741 111691 191807 111694
rect 191925 111691 191991 111694
rect 580625 111482 580691 111485
rect 583520 111482 584960 111572
rect 580625 111480 584960 111482
rect 580625 111424 580630 111480
rect 580686 111424 584960 111480
rect 580625 111422 584960 111424
rect 580625 111419 580691 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3785 107674 3851 107677
rect -960 107672 3851 107674
rect -960 107616 3790 107672
rect 3846 107616 3851 107672
rect -960 107614 3851 107616
rect -960 107524 480 107614
rect 3785 107611 3851 107614
rect 190637 106314 190703 106317
rect 190821 106314 190887 106317
rect 190637 106312 190887 106314
rect 190637 106256 190642 106312
rect 190698 106256 190826 106312
rect 190882 106256 190887 106312
rect 190637 106254 190887 106256
rect 190637 106251 190703 106254
rect 190821 106251 190887 106254
rect 403249 106314 403315 106317
rect 403433 106314 403499 106317
rect 403249 106312 403499 106314
rect 403249 106256 403254 106312
rect 403310 106256 403438 106312
rect 403494 106256 403499 106312
rect 403249 106254 403499 106256
rect 403249 106251 403315 106254
rect 403433 106251 403499 106254
rect 189022 104756 189028 104820
rect 189092 104818 189098 104820
rect 189165 104818 189231 104821
rect 189092 104816 189231 104818
rect 189092 104760 189170 104816
rect 189226 104760 189231 104816
rect 189092 104758 189231 104760
rect 189092 104756 189098 104758
rect 189165 104755 189231 104758
rect 151302 104212 151308 104276
rect 151372 104274 151378 104276
rect 151537 104274 151603 104277
rect 151372 104272 151603 104274
rect 151372 104216 151542 104272
rect 151598 104216 151603 104272
rect 151372 104214 151603 104216
rect 151372 104212 151378 104214
rect 151537 104211 151603 104214
rect 583520 99636 584960 99876
rect 169753 96658 169819 96661
rect 170029 96658 170095 96661
rect 169753 96656 170095 96658
rect 169753 96600 169758 96656
rect 169814 96600 170034 96656
rect 170090 96600 170095 96656
rect 169753 96598 170095 96600
rect 169753 96595 169819 96598
rect 170029 96595 170095 96598
rect 258073 96658 258139 96661
rect 258349 96658 258415 96661
rect 258073 96656 258415 96658
rect 258073 96600 258078 96656
rect 258134 96600 258354 96656
rect 258410 96600 258415 96656
rect 258073 96598 258415 96600
rect 258073 96595 258139 96598
rect 258349 96595 258415 96598
rect 303613 96658 303679 96661
rect 303981 96658 304047 96661
rect 303613 96656 304047 96658
rect 303613 96600 303618 96656
rect 303674 96600 303986 96656
rect 304042 96600 304047 96656
rect 303613 96598 304047 96600
rect 303613 96595 303679 96598
rect 303981 96595 304047 96598
rect 384665 96658 384731 96661
rect 384849 96658 384915 96661
rect 384665 96656 384915 96658
rect 384665 96600 384670 96656
rect 384726 96600 384854 96656
rect 384910 96600 384915 96656
rect 384665 96598 384915 96600
rect 384665 96595 384731 96598
rect 384849 96595 384915 96598
rect 245745 95434 245811 95437
rect 245745 95432 246130 95434
rect 245745 95376 245750 95432
rect 245806 95376 246130 95432
rect 245745 95374 246130 95376
rect 245745 95371 245811 95374
rect 188981 95300 189047 95301
rect 188981 95296 189028 95300
rect 189092 95298 189098 95300
rect 245929 95298 245995 95301
rect 246070 95298 246130 95374
rect 188981 95240 188986 95296
rect 188981 95236 189028 95240
rect 189092 95238 189138 95298
rect 245929 95296 246130 95298
rect 245929 95240 245934 95296
rect 245990 95240 246130 95296
rect 245929 95238 246130 95240
rect 189092 95236 189098 95238
rect 188981 95235 189047 95236
rect 245929 95235 245995 95238
rect -960 93258 480 93348
rect 3693 93258 3759 93261
rect -960 93256 3759 93258
rect -960 93200 3698 93256
rect 3754 93200 3759 93256
rect -960 93198 3759 93200
rect -960 93108 480 93198
rect 3693 93195 3759 93198
rect 151077 92850 151143 92853
rect 151302 92850 151308 92852
rect 151077 92848 151308 92850
rect 151077 92792 151082 92848
rect 151138 92792 151308 92848
rect 151077 92790 151308 92792
rect 151077 92787 151143 92790
rect 151302 92788 151308 92790
rect 151372 92788 151378 92852
rect 150985 92714 151051 92717
rect 150574 92712 151051 92714
rect 150574 92656 150990 92712
rect 151046 92656 151051 92712
rect 150574 92654 151051 92656
rect 150574 92578 150634 92654
rect 150985 92651 151051 92654
rect 150709 92578 150775 92581
rect 150574 92576 150775 92578
rect 150574 92520 150714 92576
rect 150770 92520 150775 92576
rect 150574 92518 150775 92520
rect 150709 92515 150775 92518
rect 151077 91354 151143 91357
rect 150942 91352 151143 91354
rect 150942 91296 151082 91352
rect 151138 91296 151143 91352
rect 150942 91294 151143 91296
rect 150942 91220 151002 91294
rect 151077 91291 151143 91294
rect 150934 91156 150940 91220
rect 151004 91156 151010 91220
rect 580257 87954 580323 87957
rect 583520 87954 584960 88044
rect 580257 87952 584960 87954
rect 580257 87896 580262 87952
rect 580318 87896 584960 87952
rect 580257 87894 584960 87896
rect 580257 87891 580323 87894
rect 583520 87804 584960 87894
rect 162853 87138 162919 87141
rect 224033 87138 224099 87141
rect 234797 87138 234863 87141
rect 237557 87138 237623 87141
rect 162853 87136 162962 87138
rect 162853 87080 162858 87136
rect 162914 87080 162962 87136
rect 162853 87075 162962 87080
rect 162902 87005 162962 87075
rect 223806 87136 224099 87138
rect 223806 87080 224038 87136
rect 224094 87080 224099 87136
rect 223806 87078 224099 87080
rect 223806 87005 223866 87078
rect 224033 87075 224099 87078
rect 234662 87136 234863 87138
rect 234662 87080 234802 87136
rect 234858 87080 234863 87136
rect 234662 87078 234863 87080
rect 234662 87005 234722 87078
rect 234797 87075 234863 87078
rect 237422 87136 237623 87138
rect 237422 87080 237562 87136
rect 237618 87080 237623 87136
rect 237422 87078 237623 87080
rect 237422 87005 237482 87078
rect 237557 87075 237623 87078
rect 154757 87002 154823 87005
rect 154941 87002 155007 87005
rect 154757 87000 155007 87002
rect 154757 86944 154762 87000
rect 154818 86944 154946 87000
rect 155002 86944 155007 87000
rect 154757 86942 155007 86944
rect 162902 87000 163011 87005
rect 162902 86944 162950 87000
rect 163006 86944 163011 87000
rect 162902 86942 163011 86944
rect 154757 86939 154823 86942
rect 154941 86939 155007 86942
rect 162945 86939 163011 86942
rect 190637 87002 190703 87005
rect 190821 87002 190887 87005
rect 190637 87000 190887 87002
rect 190637 86944 190642 87000
rect 190698 86944 190826 87000
rect 190882 86944 190887 87000
rect 190637 86942 190887 86944
rect 223806 87000 223915 87005
rect 223806 86944 223854 87000
rect 223910 86944 223915 87000
rect 223806 86942 223915 86944
rect 234662 87000 234771 87005
rect 234662 86944 234710 87000
rect 234766 86944 234771 87000
rect 234662 86942 234771 86944
rect 237422 87000 237531 87005
rect 237422 86944 237470 87000
rect 237526 86944 237531 87000
rect 237422 86942 237531 86944
rect 190637 86939 190703 86942
rect 190821 86939 190887 86942
rect 223849 86939 223915 86942
rect 234705 86939 234771 86942
rect 237465 86939 237531 86942
rect 384665 87002 384731 87005
rect 384849 87002 384915 87005
rect 384665 87000 384915 87002
rect 384665 86944 384670 87000
rect 384726 86944 384854 87000
rect 384910 86944 384915 87000
rect 384665 86942 384915 86944
rect 384665 86939 384731 86942
rect 384849 86939 384915 86942
rect 403249 87002 403315 87005
rect 403433 87002 403499 87005
rect 403249 87000 403499 87002
rect 403249 86944 403254 87000
rect 403310 86944 403438 87000
rect 403494 86944 403499 87000
rect 403249 86942 403499 86944
rect 403249 86939 403315 86942
rect 403433 86939 403499 86942
rect 208577 85642 208643 85645
rect 208761 85642 208827 85645
rect 208577 85640 208827 85642
rect 208577 85584 208582 85640
rect 208638 85584 208766 85640
rect 208822 85584 208827 85640
rect 208577 85582 208827 85584
rect 208577 85579 208643 85582
rect 208761 85579 208827 85582
rect 189165 85506 189231 85509
rect 189030 85504 189231 85506
rect 189030 85448 189170 85504
rect 189226 85448 189231 85504
rect 189030 85446 189231 85448
rect 189030 85370 189090 85446
rect 189165 85443 189231 85446
rect 189257 85370 189323 85373
rect 189030 85368 189323 85370
rect 189030 85312 189262 85368
rect 189318 85312 189323 85368
rect 189030 85310 189323 85312
rect 189257 85307 189323 85310
rect 150934 82996 150940 83060
rect 151004 83058 151010 83060
rect 151004 82998 151370 83058
rect 151004 82996 151010 82998
rect 151310 82924 151370 82998
rect 151302 82860 151308 82924
rect 151372 82860 151378 82924
rect 151353 81428 151419 81429
rect 151302 81426 151308 81428
rect 151262 81366 151308 81426
rect 151372 81424 151419 81428
rect 151414 81368 151419 81424
rect 151302 81364 151308 81366
rect 151372 81364 151419 81368
rect 151353 81363 151419 81364
rect 3325 80066 3391 80069
rect 152774 80066 152780 80068
rect 3325 80064 152780 80066
rect 3325 80008 3330 80064
rect 3386 80008 152780 80064
rect 3325 80006 152780 80008
rect 3325 80003 3391 80006
rect 152774 80004 152780 80006
rect 152844 80004 152850 80068
rect -960 78978 480 79068
rect 3325 78978 3391 78981
rect -960 78976 3391 78978
rect -960 78920 3330 78976
rect 3386 78920 3391 78976
rect -960 78918 3391 78920
rect -960 78828 480 78918
rect 3325 78915 3391 78918
rect 346117 77210 346183 77213
rect 346301 77210 346367 77213
rect 346117 77208 346367 77210
rect 346117 77152 346122 77208
rect 346178 77152 346306 77208
rect 346362 77152 346367 77208
rect 346117 77150 346367 77152
rect 346117 77147 346183 77150
rect 346301 77147 346367 77150
rect 579613 76258 579679 76261
rect 583520 76258 584960 76348
rect 579613 76256 584960 76258
rect 579613 76200 579618 76256
rect 579674 76200 584960 76256
rect 579613 76198 584960 76200
rect 579613 76195 579679 76198
rect 583520 76108 584960 76198
rect 151353 71906 151419 71909
rect 151486 71906 151492 71908
rect 151353 71904 151492 71906
rect 151353 71848 151358 71904
rect 151414 71848 151492 71904
rect 151353 71846 151492 71848
rect 151353 71843 151419 71846
rect 151486 71844 151492 71846
rect 151556 71844 151562 71908
rect 168649 67826 168715 67829
rect 168422 67824 168715 67826
rect 168422 67768 168654 67824
rect 168710 67768 168715 67824
rect 168422 67766 168715 67768
rect 168422 67656 168482 67766
rect 168649 67763 168715 67766
rect 263777 67826 263843 67829
rect 424777 67826 424843 67829
rect 263777 67824 263978 67826
rect 263777 67768 263782 67824
rect 263838 67768 263978 67824
rect 263777 67766 263978 67768
rect 263777 67763 263843 67766
rect 263777 67690 263843 67693
rect 263918 67690 263978 67766
rect 263777 67688 263978 67690
rect 168557 67656 168623 67659
rect 168422 67654 168623 67656
rect 168422 67598 168562 67654
rect 168618 67598 168623 67654
rect 263777 67632 263782 67688
rect 263838 67632 263978 67688
rect 263777 67630 263978 67632
rect 424550 67824 424843 67826
rect 424550 67768 424782 67824
rect 424838 67768 424843 67824
rect 424550 67766 424843 67768
rect 424550 67690 424610 67766
rect 424777 67763 424843 67766
rect 424685 67690 424751 67693
rect 424550 67688 424751 67690
rect 424550 67632 424690 67688
rect 424746 67632 424751 67688
rect 424550 67630 424751 67632
rect 263777 67627 263843 67630
rect 424685 67627 424751 67630
rect 168422 67596 168623 67598
rect 168557 67593 168623 67596
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 580349 64562 580415 64565
rect 583520 64562 584960 64652
rect 580349 64560 584960 64562
rect 580349 64504 580354 64560
rect 580410 64504 584960 64560
rect 580349 64502 584960 64504
rect 580349 64499 580415 64502
rect 583520 64412 584960 64502
rect 177941 58034 178007 58037
rect 178125 58034 178191 58037
rect 177941 58032 178191 58034
rect 177941 57976 177946 58032
rect 178002 57976 178130 58032
rect 178186 57976 178191 58032
rect 177941 57974 178191 57976
rect 177941 57971 178007 57974
rect 178125 57971 178191 57974
rect 307661 58034 307727 58037
rect 307845 58034 307911 58037
rect 307661 58032 307911 58034
rect 307661 57976 307666 58032
rect 307722 57976 307850 58032
rect 307906 57976 307911 58032
rect 307661 57974 307911 57976
rect 307661 57971 307727 57974
rect 307845 57971 307911 57974
rect 151302 55796 151308 55860
rect 151372 55858 151378 55860
rect 151670 55858 151676 55860
rect 151372 55798 151676 55858
rect 151372 55796 151378 55798
rect 151670 55796 151676 55798
rect 151740 55796 151746 55860
rect 583520 52716 584960 52956
rect 150525 51098 150591 51101
rect 150709 51098 150775 51101
rect 150525 51096 150775 51098
rect 150525 51040 150530 51096
rect 150586 51040 150714 51096
rect 150770 51040 150775 51096
rect 150525 51038 150775 51040
rect 150525 51035 150591 51038
rect 150709 51035 150775 51038
rect -960 50146 480 50236
rect 3601 50146 3667 50149
rect -960 50144 3667 50146
rect -960 50088 3606 50144
rect 3662 50088 3667 50144
rect -960 50086 3667 50088
rect -960 49996 480 50086
rect 3601 50083 3667 50086
rect 263685 48242 263751 48245
rect 307937 48244 308003 48245
rect 263550 48240 263751 48242
rect 263550 48184 263690 48240
rect 263746 48184 263751 48240
rect 263550 48182 263751 48184
rect 263550 48106 263610 48182
rect 263685 48179 263751 48182
rect 307886 48180 307892 48244
rect 307956 48242 308003 48244
rect 307956 48240 308048 48242
rect 307998 48184 308048 48240
rect 307956 48182 308048 48184
rect 307956 48180 308003 48182
rect 307937 48179 308003 48180
rect 263777 48106 263843 48109
rect 263550 48104 263843 48106
rect 263550 48048 263782 48104
rect 263838 48048 263843 48104
rect 263550 48046 263843 48048
rect 263777 48043 263843 48046
rect 191925 44162 191991 44165
rect 192109 44162 192175 44165
rect 191925 44160 192175 44162
rect 191925 44104 191930 44160
rect 191986 44104 192114 44160
rect 192170 44104 192175 44160
rect 191925 44102 192175 44104
rect 191925 44099 191991 44102
rect 192109 44099 192175 44102
rect 194501 44162 194567 44165
rect 194777 44162 194843 44165
rect 194501 44160 194843 44162
rect 194501 44104 194506 44160
rect 194562 44104 194782 44160
rect 194838 44104 194843 44160
rect 194501 44102 194843 44104
rect 194501 44099 194567 44102
rect 194777 44099 194843 44102
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 238661 40626 238727 40629
rect 240041 40626 240107 40629
rect 238661 40624 240107 40626
rect 238661 40568 238666 40624
rect 238722 40568 240046 40624
rect 240102 40568 240107 40624
rect 238661 40566 240107 40568
rect 238661 40563 238727 40566
rect 240041 40563 240107 40566
rect 462262 40428 462268 40492
rect 462332 40490 462338 40492
rect 471881 40490 471947 40493
rect 462332 40488 471947 40490
rect 462332 40432 471886 40488
rect 471942 40432 471947 40488
rect 462332 40430 471947 40432
rect 462332 40428 462338 40430
rect 471881 40427 471947 40430
rect 176377 40354 176443 40357
rect 167686 40352 176443 40354
rect 167686 40296 176382 40352
rect 176438 40296 176443 40352
rect 167686 40294 176443 40296
rect 154062 40020 154068 40084
rect 154132 40082 154138 40084
rect 167686 40082 167746 40294
rect 176377 40291 176443 40294
rect 176561 40354 176627 40357
rect 229001 40354 229067 40357
rect 240041 40354 240107 40357
rect 249742 40354 249748 40356
rect 176561 40352 177314 40354
rect 176561 40296 176566 40352
rect 176622 40296 177314 40352
rect 176561 40294 177314 40296
rect 176561 40291 176627 40294
rect 177254 40218 177314 40294
rect 229001 40352 229202 40354
rect 229001 40296 229006 40352
rect 229062 40296 229202 40352
rect 229001 40294 229202 40296
rect 229001 40291 229067 40294
rect 183502 40218 183508 40220
rect 177254 40158 183508 40218
rect 183502 40156 183508 40158
rect 183572 40156 183578 40220
rect 201493 40218 201559 40221
rect 195286 40216 201559 40218
rect 195286 40160 201498 40216
rect 201554 40160 201559 40216
rect 195286 40158 201559 40160
rect 195286 40082 195346 40158
rect 201493 40155 201559 40158
rect 154132 40022 167746 40082
rect 183694 40022 195346 40082
rect 219341 40084 219407 40085
rect 219341 40080 219388 40084
rect 219452 40082 219458 40084
rect 229142 40082 229202 40294
rect 240041 40352 249748 40354
rect 240041 40296 240046 40352
rect 240102 40296 249748 40352
rect 240041 40294 249748 40296
rect 240041 40291 240107 40294
rect 249742 40292 249748 40294
rect 249812 40292 249818 40356
rect 447225 40354 447291 40357
rect 482921 40354 482987 40357
rect 273118 40294 282930 40354
rect 238661 40082 238727 40085
rect 273118 40082 273178 40294
rect 219341 40024 219346 40080
rect 154132 40020 154138 40022
rect 183502 39884 183508 39948
rect 183572 39946 183578 39948
rect 183694 39946 183754 40022
rect 219341 40020 219388 40024
rect 219452 40022 219534 40082
rect 229142 40080 238727 40082
rect 229142 40024 238666 40080
rect 238722 40024 238727 40080
rect 229142 40022 238727 40024
rect 219452 40020 219458 40022
rect 219341 40019 219407 40020
rect 238661 40019 238727 40022
rect 260790 40022 273178 40082
rect 282870 40082 282930 40294
rect 447225 40352 458834 40354
rect 447225 40296 447230 40352
rect 447286 40296 458834 40352
rect 447225 40294 458834 40296
rect 447225 40291 447291 40294
rect 302141 40218 302207 40221
rect 292622 40216 302207 40218
rect 292622 40160 302146 40216
rect 302202 40160 302207 40216
rect 292622 40158 302207 40160
rect 292622 40082 292682 40158
rect 302141 40155 302207 40158
rect 302325 40218 302391 40221
rect 321277 40218 321343 40221
rect 302325 40216 311818 40218
rect 302325 40160 302330 40216
rect 302386 40160 311818 40216
rect 302325 40158 311818 40160
rect 302325 40155 302391 40158
rect 282870 40022 292682 40082
rect 311758 40082 311818 40158
rect 311942 40216 321343 40218
rect 311942 40160 321282 40216
rect 321338 40160 321343 40216
rect 311942 40158 321343 40160
rect 311942 40082 312002 40158
rect 321277 40155 321343 40158
rect 321553 40218 321619 40221
rect 340689 40218 340755 40221
rect 321553 40216 328378 40218
rect 321553 40160 321558 40216
rect 321614 40160 328378 40216
rect 321553 40158 328378 40160
rect 321553 40155 321619 40158
rect 311758 40022 312002 40082
rect 328318 40082 328378 40158
rect 331262 40216 340755 40218
rect 331262 40160 340694 40216
rect 340750 40160 340755 40216
rect 331262 40158 340755 40160
rect 331262 40082 331322 40158
rect 340689 40155 340755 40158
rect 340965 40218 341031 40221
rect 359917 40218 359983 40221
rect 340965 40216 350458 40218
rect 340965 40160 340970 40216
rect 341026 40160 350458 40216
rect 340965 40158 350458 40160
rect 340965 40155 341031 40158
rect 328318 40022 331322 40082
rect 350398 40082 350458 40158
rect 350582 40216 359983 40218
rect 350582 40160 359922 40216
rect 359978 40160 359983 40216
rect 350582 40158 359983 40160
rect 350582 40082 350642 40158
rect 359917 40155 359983 40158
rect 360193 40218 360259 40221
rect 437197 40218 437263 40221
rect 360193 40216 367018 40218
rect 360193 40160 360198 40216
rect 360254 40160 367018 40216
rect 360193 40158 367018 40160
rect 360193 40155 360259 40158
rect 350398 40022 350642 40082
rect 366958 40082 367018 40158
rect 369902 40158 389098 40218
rect 369902 40082 369962 40158
rect 366958 40022 369962 40082
rect 389038 40082 389098 40158
rect 389222 40158 405658 40218
rect 389222 40082 389282 40158
rect 389038 40022 389282 40082
rect 405598 40082 405658 40158
rect 408542 40158 427738 40218
rect 408542 40082 408602 40158
rect 405598 40022 408602 40082
rect 427678 40082 427738 40158
rect 427862 40216 437263 40218
rect 427862 40160 437202 40216
rect 437258 40160 437263 40216
rect 427862 40158 437263 40160
rect 458774 40218 458834 40294
rect 482921 40352 489930 40354
rect 482921 40296 482926 40352
rect 482982 40296 489930 40352
rect 482921 40294 489930 40296
rect 482921 40291 482987 40294
rect 462262 40218 462268 40220
rect 458774 40158 462268 40218
rect 427862 40082 427922 40158
rect 437197 40155 437263 40158
rect 462262 40156 462268 40158
rect 462332 40156 462338 40220
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 444373 40082 444439 40085
rect 427678 40022 427922 40082
rect 444238 40080 444439 40082
rect 444238 40024 444378 40080
rect 444434 40024 444439 40080
rect 444238 40022 444439 40024
rect 183572 39886 183754 39946
rect 183572 39884 183578 39886
rect 249742 39884 249748 39948
rect 249812 39946 249818 39948
rect 260790 39946 260850 40022
rect 249812 39886 260850 39946
rect 249812 39884 249818 39886
rect 219382 39748 219388 39812
rect 219452 39810 219458 39812
rect 229001 39810 229067 39813
rect 219452 39808 229067 39810
rect 219452 39752 229006 39808
rect 229062 39752 229067 39808
rect 219452 39750 229067 39752
rect 219452 39748 219458 39750
rect 229001 39747 229067 39750
rect 437197 39810 437263 39813
rect 444238 39810 444298 40022
rect 444373 40019 444439 40022
rect 471881 40082 471947 40085
rect 476021 40082 476087 40085
rect 471881 40080 476087 40082
rect 471881 40024 471886 40080
rect 471942 40024 476026 40080
rect 476082 40024 476087 40080
rect 471881 40022 476087 40024
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect 471881 40019 471947 40022
rect 476021 40019 476087 40022
rect 437197 39808 444298 39810
rect 437197 39752 437202 39808
rect 437258 39752 444298 39808
rect 437197 39750 444298 39752
rect 437197 39747 437263 39750
rect 403893 38858 403959 38861
rect 403893 38856 404002 38858
rect 403893 38800 403898 38856
rect 403954 38800 404002 38856
rect 403893 38795 404002 38800
rect 307886 38660 307892 38724
rect 307956 38722 307962 38724
rect 308029 38722 308095 38725
rect 307956 38720 308095 38722
rect 307956 38664 308034 38720
rect 308090 38664 308095 38720
rect 307956 38662 308095 38664
rect 307956 38660 307962 38662
rect 308029 38659 308095 38662
rect 403801 38722 403867 38725
rect 403942 38722 404002 38795
rect 403801 38720 404002 38722
rect 403801 38664 403806 38720
rect 403862 38664 404002 38720
rect 403801 38662 404002 38664
rect 403801 38659 403867 38662
rect 379145 37226 379211 37229
rect 379329 37226 379395 37229
rect 379145 37224 379395 37226
rect 379145 37168 379150 37224
rect 379206 37168 379334 37224
rect 379390 37168 379395 37224
rect 379145 37166 379395 37168
rect 379145 37163 379211 37166
rect 379329 37163 379395 37166
rect -960 35866 480 35956
rect 3509 35866 3575 35869
rect -960 35864 3575 35866
rect -960 35808 3514 35864
rect 3570 35808 3575 35864
rect -960 35806 3575 35808
rect -960 35716 480 35806
rect 3509 35803 3575 35806
rect 150525 33146 150591 33149
rect 150709 33146 150775 33149
rect 150525 33144 150775 33146
rect 150525 33088 150530 33144
rect 150586 33088 150714 33144
rect 150770 33088 150775 33144
rect 150525 33086 150775 33088
rect 150525 33083 150591 33086
rect 150709 33083 150775 33086
rect 579613 29338 579679 29341
rect 583520 29338 584960 29428
rect 579613 29336 584960 29338
rect 579613 29280 579618 29336
rect 579674 29280 584960 29336
rect 579613 29278 584960 29280
rect 579613 29275 579679 29278
rect 583520 29188 584960 29278
rect 189257 27842 189323 27845
rect 189030 27840 189323 27842
rect 189030 27784 189262 27840
rect 189318 27784 189323 27840
rect 189030 27782 189323 27784
rect 189030 27706 189090 27782
rect 189257 27779 189323 27782
rect 189165 27706 189231 27709
rect 189030 27704 189231 27706
rect 189030 27648 189170 27704
rect 189226 27648 189231 27704
rect 189030 27646 189231 27648
rect 189165 27643 189231 27646
rect 191741 26210 191807 26213
rect 191925 26210 191991 26213
rect 191741 26208 191991 26210
rect 191741 26152 191746 26208
rect 191802 26152 191930 26208
rect 191986 26152 191991 26208
rect 191741 26150 191991 26152
rect 191741 26147 191807 26150
rect 191925 26147 191991 26150
rect -960 21450 480 21540
rect 3417 21450 3483 21453
rect -960 21448 3483 21450
rect -960 21392 3422 21448
rect 3478 21392 3483 21448
rect -960 21390 3483 21392
rect -960 21300 480 21390
rect 3417 21387 3483 21390
rect 583520 17642 584960 17732
rect 583342 17582 584960 17642
rect 462262 17036 462268 17100
rect 462332 17098 462338 17100
rect 471881 17098 471947 17101
rect 462332 17096 471947 17098
rect 462332 17040 471886 17096
rect 471942 17040 471947 17096
rect 462332 17038 471947 17040
rect 462332 17036 462338 17038
rect 471881 17035 471947 17038
rect 447225 16962 447291 16965
rect 482921 16962 482987 16965
rect 273118 16902 282930 16962
rect 151670 16628 151676 16692
rect 151740 16690 151746 16692
rect 173893 16690 173959 16693
rect 151740 16688 173959 16690
rect 151740 16632 173898 16688
rect 173954 16632 173959 16688
rect 151740 16630 173959 16632
rect 151740 16628 151746 16630
rect 173893 16627 173959 16630
rect 183461 16690 183527 16693
rect 273118 16690 273178 16902
rect 183461 16688 273178 16690
rect 183461 16632 183466 16688
rect 183522 16632 273178 16688
rect 183461 16630 273178 16632
rect 282870 16690 282930 16902
rect 447225 16960 458834 16962
rect 447225 16904 447230 16960
rect 447286 16904 458834 16960
rect 447225 16902 458834 16904
rect 447225 16899 447291 16902
rect 302141 16826 302207 16829
rect 292622 16824 302207 16826
rect 292622 16768 302146 16824
rect 302202 16768 302207 16824
rect 292622 16766 302207 16768
rect 292622 16690 292682 16766
rect 302141 16763 302207 16766
rect 302325 16826 302391 16829
rect 318793 16826 318859 16829
rect 302325 16824 311818 16826
rect 302325 16768 302330 16824
rect 302386 16768 311818 16824
rect 302325 16766 311818 16768
rect 302325 16763 302391 16766
rect 282870 16630 292682 16690
rect 311758 16690 311818 16766
rect 311942 16824 318859 16826
rect 311942 16768 318798 16824
rect 318854 16768 318859 16824
rect 311942 16766 318859 16768
rect 311942 16690 312002 16766
rect 318793 16763 318859 16766
rect 321553 16826 321619 16829
rect 338205 16826 338271 16829
rect 321553 16824 328378 16826
rect 321553 16768 321558 16824
rect 321614 16768 328378 16824
rect 321553 16766 328378 16768
rect 321553 16763 321619 16766
rect 311758 16630 312002 16690
rect 328318 16690 328378 16766
rect 331262 16824 338271 16826
rect 331262 16768 338210 16824
rect 338266 16768 338271 16824
rect 331262 16766 338271 16768
rect 331262 16690 331322 16766
rect 338205 16763 338271 16766
rect 342621 16826 342687 16829
rect 359917 16826 359983 16829
rect 342621 16824 350458 16826
rect 342621 16768 342626 16824
rect 342682 16768 350458 16824
rect 342621 16766 350458 16768
rect 342621 16763 342687 16766
rect 328318 16630 331322 16690
rect 350398 16690 350458 16766
rect 350582 16824 359983 16826
rect 350582 16768 359922 16824
rect 359978 16768 359983 16824
rect 350582 16766 359983 16768
rect 350582 16690 350642 16766
rect 359917 16763 359983 16766
rect 362217 16826 362283 16829
rect 379237 16826 379303 16829
rect 362217 16824 367018 16826
rect 362217 16768 362222 16824
rect 362278 16768 367018 16824
rect 362217 16766 367018 16768
rect 362217 16763 362283 16766
rect 350398 16630 350642 16690
rect 366958 16690 367018 16766
rect 369902 16824 379303 16826
rect 369902 16768 379242 16824
rect 379298 16768 379303 16824
rect 369902 16766 379303 16768
rect 369902 16690 369962 16766
rect 379237 16763 379303 16766
rect 379605 16826 379671 16829
rect 398649 16826 398715 16829
rect 379605 16824 389098 16826
rect 379605 16768 379610 16824
rect 379666 16768 389098 16824
rect 379605 16766 389098 16768
rect 379605 16763 379671 16766
rect 366958 16630 369962 16690
rect 389038 16690 389098 16766
rect 389222 16824 398715 16826
rect 389222 16768 398654 16824
rect 398710 16768 398715 16824
rect 389222 16766 398715 16768
rect 389222 16690 389282 16766
rect 398649 16763 398715 16766
rect 400857 16826 400923 16829
rect 417969 16826 418035 16829
rect 400857 16824 405658 16826
rect 400857 16768 400862 16824
rect 400918 16768 405658 16824
rect 400857 16766 405658 16768
rect 400857 16763 400923 16766
rect 389038 16630 389282 16690
rect 405598 16690 405658 16766
rect 408542 16824 418035 16826
rect 408542 16768 417974 16824
rect 418030 16768 418035 16824
rect 408542 16766 418035 16768
rect 408542 16690 408602 16766
rect 417969 16763 418035 16766
rect 418245 16826 418311 16829
rect 437197 16826 437263 16829
rect 418245 16824 424978 16826
rect 418245 16768 418250 16824
rect 418306 16768 424978 16824
rect 418245 16766 424978 16768
rect 418245 16763 418311 16766
rect 405598 16630 408602 16690
rect 424918 16690 424978 16766
rect 427862 16824 437263 16826
rect 427862 16768 437202 16824
rect 437258 16768 437263 16824
rect 427862 16766 437263 16768
rect 458774 16826 458834 16902
rect 482921 16960 489930 16962
rect 482921 16904 482926 16960
rect 482982 16904 489930 16960
rect 482921 16902 489930 16904
rect 482921 16899 482987 16902
rect 462262 16826 462268 16828
rect 458774 16766 462268 16826
rect 427862 16690 427922 16766
rect 437197 16763 437263 16766
rect 462262 16764 462268 16766
rect 462332 16764 462338 16828
rect 489870 16826 489930 16902
rect 499622 16902 509250 16962
rect 489870 16766 499498 16826
rect 444373 16690 444439 16693
rect 424918 16630 427922 16690
rect 444238 16688 444439 16690
rect 444238 16632 444378 16688
rect 444434 16632 444439 16688
rect 444238 16630 444439 16632
rect 183461 16627 183527 16630
rect 437197 16418 437263 16421
rect 444238 16418 444298 16630
rect 444373 16627 444439 16630
rect 471881 16690 471947 16693
rect 476021 16690 476087 16693
rect 471881 16688 476087 16690
rect 471881 16632 471886 16688
rect 471942 16632 476026 16688
rect 476082 16632 476087 16688
rect 471881 16630 476087 16632
rect 499438 16690 499498 16766
rect 499622 16690 499682 16902
rect 509190 16826 509250 16902
rect 518942 16902 528570 16962
rect 509190 16766 518818 16826
rect 499438 16630 499682 16690
rect 518758 16690 518818 16766
rect 518942 16690 519002 16902
rect 528510 16826 528570 16902
rect 538262 16902 547890 16962
rect 528510 16766 538138 16826
rect 518758 16630 519002 16690
rect 538078 16690 538138 16766
rect 538262 16690 538322 16902
rect 547830 16826 547890 16902
rect 557582 16902 567210 16962
rect 547830 16766 557458 16826
rect 538078 16630 538322 16690
rect 557398 16690 557458 16766
rect 557582 16690 557642 16902
rect 567150 16826 567210 16902
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 567150 16766 576778 16826
rect 557398 16630 557642 16690
rect 576718 16690 576778 16766
rect 576902 16766 583402 16826
rect 576902 16690 576962 16766
rect 576718 16630 576962 16690
rect 471881 16627 471947 16630
rect 476021 16627 476087 16630
rect 437197 16416 444298 16418
rect 437197 16360 437202 16416
rect 437258 16360 444298 16416
rect 437197 16358 444298 16360
rect 437197 16355 437263 16358
rect 152089 15194 152155 15197
rect 152273 15194 152339 15197
rect 152089 15192 152339 15194
rect 152089 15136 152094 15192
rect 152150 15136 152278 15192
rect 152334 15136 152339 15192
rect 152089 15134 152339 15136
rect 152089 15131 152155 15134
rect 152273 15131 152339 15134
rect 27889 8938 27955 8941
rect 164417 8938 164483 8941
rect 27889 8936 164483 8938
rect 27889 8880 27894 8936
rect 27950 8880 164422 8936
rect 164478 8880 164483 8936
rect 27889 8878 164483 8880
rect 27889 8875 27955 8878
rect 164417 8875 164483 8878
rect 70669 7578 70735 7581
rect 185025 7578 185091 7581
rect 70669 7576 185091 7578
rect 70669 7520 70674 7576
rect 70730 7520 185030 7576
rect 185086 7520 185091 7576
rect 70669 7518 185091 7520
rect 70669 7515 70735 7518
rect 185025 7515 185091 7518
rect 442717 7578 442783 7581
rect 570229 7578 570295 7581
rect 442717 7576 570295 7578
rect 442717 7520 442722 7576
rect 442778 7520 570234 7576
rect 570290 7520 570295 7576
rect 442717 7518 570295 7520
rect 442717 7515 442783 7518
rect 570229 7515 570295 7518
rect -960 7170 480 7260
rect 2773 7170 2839 7173
rect -960 7168 2839 7170
rect -960 7112 2778 7168
rect 2834 7112 2839 7168
rect -960 7110 2839 7112
rect -960 7020 480 7110
rect 2773 7107 2839 7110
rect 44541 6354 44607 6357
rect 172605 6354 172671 6357
rect 44541 6352 172671 6354
rect 44541 6296 44546 6352
rect 44602 6296 172610 6352
rect 172666 6296 172671 6352
rect 44541 6294 172671 6296
rect 44541 6291 44607 6294
rect 172605 6291 172671 6294
rect 37365 6218 37431 6221
rect 168465 6218 168531 6221
rect 37365 6216 168531 6218
rect 37365 6160 37370 6216
rect 37426 6160 168470 6216
rect 168526 6160 168531 6216
rect 37365 6158 168531 6160
rect 37365 6155 37431 6158
rect 168465 6155 168531 6158
rect 440141 6218 440207 6221
rect 563145 6218 563211 6221
rect 440141 6216 563211 6218
rect 440141 6160 440146 6216
rect 440202 6160 563150 6216
rect 563206 6160 563211 6216
rect 440141 6158 563211 6160
rect 440141 6155 440207 6158
rect 563145 6155 563211 6158
rect 583520 5796 584960 6036
rect 151997 5674 152063 5677
rect 152273 5674 152339 5677
rect 151997 5672 152339 5674
rect 151997 5616 152002 5672
rect 152058 5616 152278 5672
rect 152334 5616 152339 5672
rect 151997 5614 152339 5616
rect 151997 5611 152063 5614
rect 152273 5611 152339 5614
rect 93853 5402 93919 5405
rect 103421 5402 103487 5405
rect 93853 5400 103487 5402
rect 93853 5344 93858 5400
rect 93914 5344 103426 5400
rect 103482 5344 103487 5400
rect 93853 5342 103487 5344
rect 93853 5339 93919 5342
rect 103421 5339 103487 5342
rect 113173 5402 113239 5405
rect 122649 5402 122715 5405
rect 113173 5400 122715 5402
rect 113173 5344 113178 5400
rect 113234 5344 122654 5400
rect 122710 5344 122715 5400
rect 113173 5342 122715 5344
rect 113173 5339 113239 5342
rect 122649 5339 122715 5342
rect 132493 5402 132559 5405
rect 141969 5402 142035 5405
rect 132493 5400 142035 5402
rect 132493 5344 132498 5400
rect 132554 5344 141974 5400
rect 142030 5344 142035 5400
rect 132493 5342 142035 5344
rect 132493 5339 132559 5342
rect 141969 5339 142035 5342
rect 178677 5402 178743 5405
rect 183461 5402 183527 5405
rect 178677 5400 183527 5402
rect 178677 5344 178682 5400
rect 178738 5344 183466 5400
rect 183522 5344 183527 5400
rect 178677 5342 183527 5344
rect 178677 5339 178743 5342
rect 183461 5339 183527 5342
rect 420085 5266 420151 5269
rect 424133 5266 424199 5269
rect 420085 5264 424199 5266
rect 420085 5208 420090 5264
rect 420146 5208 424138 5264
rect 424194 5208 424199 5264
rect 420085 5206 424199 5208
rect 420085 5203 420151 5206
rect 424133 5203 424199 5206
rect 142153 4994 142219 4997
rect 150893 4994 150959 4997
rect 142153 4992 150959 4994
rect 142153 4936 142158 4992
rect 142214 4936 150898 4992
rect 150954 4936 150959 4992
rect 142153 4934 150959 4936
rect 142153 4931 142219 4934
rect 150893 4931 150959 4934
rect 379329 4994 379395 4997
rect 379513 4994 379579 4997
rect 379329 4992 379579 4994
rect 379329 4936 379334 4992
rect 379390 4936 379518 4992
rect 379574 4936 379579 4992
rect 379329 4934 379579 4936
rect 379329 4931 379395 4934
rect 379513 4931 379579 4934
rect 398741 4994 398807 4997
rect 403617 4994 403683 4997
rect 398741 4992 403683 4994
rect 398741 4936 398746 4992
rect 398802 4936 403622 4992
rect 403678 4936 403683 4992
rect 398741 4934 403683 4936
rect 398741 4931 398807 4934
rect 403617 4931 403683 4934
rect 12433 4858 12499 4861
rect 155953 4858 156019 4861
rect 12433 4856 156019 4858
rect 12433 4800 12438 4856
rect 12494 4800 155958 4856
rect 156014 4800 156019 4856
rect 12433 4798 156019 4800
rect 12433 4795 12499 4798
rect 155953 4795 156019 4798
rect 380801 4858 380867 4861
rect 447777 4858 447843 4861
rect 380801 4856 447843 4858
rect 380801 4800 380806 4856
rect 380862 4800 447782 4856
rect 447838 4800 447843 4856
rect 380801 4798 447843 4800
rect 380801 4795 380867 4798
rect 447777 4795 447843 4798
rect 448421 4858 448487 4861
rect 579797 4858 579863 4861
rect 448421 4856 579863 4858
rect 448421 4800 448426 4856
rect 448482 4800 579802 4856
rect 579858 4800 579863 4856
rect 448421 4798 579863 4800
rect 448421 4795 448487 4798
rect 579797 4795 579863 4798
rect 398925 4722 398991 4725
rect 404997 4722 405063 4725
rect 398925 4720 405063 4722
rect 398925 4664 398930 4720
rect 398986 4664 405002 4720
rect 405058 4664 405063 4720
rect 398925 4662 405063 4664
rect 398925 4659 398991 4662
rect 404997 4659 405063 4662
rect 391289 4586 391355 4589
rect 394693 4586 394759 4589
rect 391289 4584 394759 4586
rect 391289 4528 391294 4584
rect 391350 4528 394698 4584
rect 394754 4528 394759 4584
rect 391289 4526 394759 4528
rect 391289 4523 391355 4526
rect 394693 4523 394759 4526
rect 398833 4586 398899 4589
rect 401409 4586 401475 4589
rect 398833 4584 401475 4586
rect 398833 4528 398838 4584
rect 398894 4528 401414 4584
rect 401470 4528 401475 4584
rect 398833 4526 401475 4528
rect 398833 4523 398899 4526
rect 401409 4523 401475 4526
rect 427629 4450 427695 4453
rect 427905 4450 427971 4453
rect 427629 4448 427971 4450
rect 427629 4392 427634 4448
rect 427690 4392 427910 4448
rect 427966 4392 427971 4448
rect 427629 4390 427971 4392
rect 427629 4387 427695 4390
rect 427905 4387 427971 4390
rect 231209 3634 231275 3637
rect 232497 3634 232563 3637
rect 231209 3632 232563 3634
rect 231209 3576 231214 3632
rect 231270 3576 232502 3632
rect 232558 3576 232563 3632
rect 231209 3574 232563 3576
rect 231209 3571 231275 3574
rect 232497 3571 232563 3574
rect 5257 3362 5323 3365
rect 151997 3362 152063 3365
rect 5257 3360 152063 3362
rect 5257 3304 5262 3360
rect 5318 3304 152002 3360
rect 152058 3304 152063 3360
rect 5257 3302 152063 3304
rect 5257 3299 5323 3302
rect 151997 3299 152063 3302
rect 449801 3362 449867 3365
rect 582189 3362 582255 3365
rect 449801 3360 582255 3362
rect 449801 3304 449806 3360
rect 449862 3304 582194 3360
rect 582250 3304 582255 3360
rect 449801 3302 582255 3304
rect 449801 3299 449867 3302
rect 582189 3299 582255 3302
<< via3 >>
rect 447732 549068 447796 549132
rect 446628 548932 446692 548996
rect 152780 548796 152844 548860
rect 446444 548660 446508 548724
rect 151860 548524 151924 548588
rect 152228 545260 152292 545324
rect 152964 545124 153028 545188
rect 151676 544580 151740 544644
rect 154068 544640 154132 544644
rect 154068 544584 154082 544640
rect 154082 544584 154132 544640
rect 154068 544580 154132 544584
rect 203196 544640 203260 544644
rect 203196 544584 203210 544640
rect 203210 544584 203260 544640
rect 203196 544580 203260 544584
rect 205404 544640 205468 544644
rect 205404 544584 205454 544640
rect 205454 544584 205468 544640
rect 205404 544580 205468 544584
rect 208164 544580 208228 544644
rect 213500 544640 213564 544644
rect 213500 544584 213514 544640
rect 213514 544584 213564 544640
rect 213500 544580 213564 544584
rect 221412 544580 221476 544644
rect 231532 544640 231596 544644
rect 231532 544584 231582 544640
rect 231582 544584 231596 544640
rect 231532 544580 231596 544584
rect 386460 544640 386524 544644
rect 386460 544584 386510 544640
rect 386510 544584 386524 544640
rect 386460 544580 386524 544584
rect 226932 543900 226996 543964
rect 231716 543900 231780 543964
rect 221412 543628 221476 543692
rect 213500 543492 213564 543556
rect 208164 543356 208228 543420
rect 205404 543220 205468 543284
rect 226932 543220 226996 543284
rect 231532 543220 231596 543284
rect 231716 543220 231780 543284
rect 203196 543084 203260 543148
rect 231164 543084 231228 543148
rect 231348 542948 231412 543012
rect 231900 543084 231964 543148
rect 231716 542948 231780 543012
rect 386460 542948 386524 543012
rect 152228 536148 152292 536212
rect 152964 536148 153028 536212
rect 152780 521596 152844 521660
rect 152596 520236 152660 520300
rect 152044 520100 152108 520164
rect 152596 520100 152660 520164
rect 150756 511940 150820 512004
rect 151492 511940 151556 512004
rect 152044 510580 152108 510644
rect 152780 510580 152844 510644
rect 152964 510444 153028 510508
rect 152964 510036 153028 510100
rect 150756 502556 150820 502620
rect 151124 502420 151188 502484
rect 152596 491404 152660 491468
rect 152780 491268 152844 491332
rect 152780 491132 152844 491196
rect 152044 490860 152108 490924
rect 152044 481612 152108 481676
rect 152780 481612 152844 481676
rect 152228 481476 152292 481540
rect 152780 481476 152844 481540
rect 152228 471956 152292 472020
rect 152780 471956 152844 472020
rect 152780 463524 152844 463588
rect 153148 463524 153212 463588
rect 151492 456860 151556 456924
rect 151308 456588 151372 456652
rect 152780 454140 152844 454204
rect 153148 454140 153212 454204
rect 152228 452508 152292 452572
rect 152780 452508 152844 452572
rect 151308 447204 151372 447268
rect 151492 446932 151556 446996
rect 152228 443124 152292 443188
rect 152596 442988 152660 443052
rect 151492 441492 151556 441556
rect 150940 441356 151004 441420
rect 150940 431972 151004 432036
rect 151676 431972 151740 432036
rect 151676 427892 151740 427956
rect 151676 427756 151740 427820
rect 151676 423676 151740 423740
rect 151676 423540 151740 423604
rect 152228 423540 152292 423604
rect 152780 423540 152844 423604
rect 152228 414156 152292 414220
rect 152780 414020 152844 414084
rect 151308 412524 151372 412588
rect 151492 412388 151556 412452
rect 152228 404228 152292 404292
rect 152780 404228 152844 404292
rect 151492 402868 151556 402932
rect 151124 402732 151188 402796
rect 152228 394844 152292 394908
rect 152780 394708 152844 394772
rect 151124 393348 151188 393412
rect 151676 393348 151740 393412
rect 151676 389268 151740 389332
rect 151492 388996 151556 389060
rect 152228 365604 152292 365668
rect 152780 365604 152844 365668
rect 151492 364380 151556 364444
rect 151676 364380 151740 364444
rect 447732 357716 447796 357780
rect 151676 356220 151740 356284
rect 152228 356220 152292 356284
rect 151492 356084 151556 356148
rect 152780 356084 152844 356148
rect 151492 348468 151556 348532
rect 152228 348468 152292 348532
rect 151860 346564 151924 346628
rect 151860 346156 151924 346220
rect 152044 335412 152108 335476
rect 152228 335412 152292 335476
rect 151860 335276 151924 335340
rect 152044 335140 152108 335204
rect 152228 335140 152292 335204
rect 151860 334052 151924 334116
rect 152780 327524 152844 327588
rect 152964 327524 153028 327588
rect 151860 327388 151924 327452
rect 151492 327116 151556 327180
rect 152780 327116 152844 327180
rect 152964 327116 153028 327180
rect 152228 326980 152292 327044
rect 152780 326980 152844 327044
rect 150756 325620 150820 325684
rect 151492 325620 151556 325684
rect 152228 317596 152292 317660
rect 152780 317460 152844 317524
rect 150756 316236 150820 316300
rect 151308 316236 151372 316300
rect 151308 315964 151372 316028
rect 151492 315964 151556 316028
rect 151308 314604 151372 314668
rect 151492 314604 151556 314668
rect 152228 307668 152292 307732
rect 152780 307668 152844 307732
rect 151124 304948 151188 305012
rect 151308 304948 151372 305012
rect 446628 298420 446692 298484
rect 152228 298284 152292 298348
rect 152780 298148 152844 298212
rect 151124 296788 151188 296852
rect 151676 296788 151740 296852
rect 151676 292708 151740 292772
rect 151492 292436 151556 292500
rect 152228 288356 152292 288420
rect 152780 288356 152844 288420
rect 151124 280740 151188 280804
rect 151492 280740 151556 280804
rect 152228 278972 152292 279036
rect 152780 278836 152844 278900
rect 151124 275980 151188 276044
rect 151492 275980 151556 276044
rect 151124 266188 151188 266252
rect 151492 266188 151556 266252
rect 152780 259388 152844 259452
rect 152596 259252 152660 259316
rect 151124 256668 151188 256732
rect 151492 256668 151556 256732
rect 446812 251500 446876 251564
rect 152596 248508 152660 248572
rect 152780 248372 152844 248436
rect 152780 248236 152844 248300
rect 153516 248236 153580 248300
rect 151124 246876 151188 246940
rect 151492 246876 151556 246940
rect 152964 244428 153028 244492
rect 152964 244156 153028 244220
rect 153148 238716 153212 238780
rect 153516 238716 153580 238780
rect 151124 237356 151188 237420
rect 151492 237356 151556 237420
rect 151492 237220 151556 237284
rect 153148 222260 153212 222324
rect 153332 221988 153396 222052
rect 151492 220900 151556 220964
rect 152780 215248 152844 215252
rect 152780 215192 152794 215248
rect 152794 215192 152844 215248
rect 152780 215188 152844 215192
rect 152780 215052 152844 215116
rect 153148 215052 153212 215116
rect 151492 212468 151556 212532
rect 151308 212332 151372 212396
rect 151308 206212 151372 206276
rect 151860 201316 151924 201380
rect 151860 196556 151924 196620
rect 151676 193216 151740 193220
rect 151676 193160 151690 193216
rect 151690 193160 151740 193216
rect 151676 193156 151740 193160
rect 151308 177244 151372 177308
rect 151860 165548 151924 165612
rect 151124 165412 151188 165476
rect 151124 156572 151188 156636
rect 151492 156572 151556 156636
rect 151492 147732 151556 147796
rect 151308 147460 151372 147524
rect 152964 122708 153028 122772
rect 151308 114684 151372 114748
rect 151492 114548 151556 114612
rect 151492 113052 151556 113116
rect 189028 104756 189092 104820
rect 151308 104212 151372 104276
rect 189028 95296 189092 95300
rect 189028 95240 189042 95296
rect 189042 95240 189092 95296
rect 189028 95236 189092 95240
rect 151308 92788 151372 92852
rect 150940 91156 151004 91220
rect 150940 82996 151004 83060
rect 151308 82860 151372 82924
rect 151308 81424 151372 81428
rect 151308 81368 151358 81424
rect 151358 81368 151372 81424
rect 151308 81364 151372 81368
rect 152780 80004 152844 80068
rect 151492 71844 151556 71908
rect 151308 55796 151372 55860
rect 151676 55796 151740 55860
rect 307892 48240 307956 48244
rect 307892 48184 307942 48240
rect 307942 48184 307956 48240
rect 307892 48180 307956 48184
rect 462268 40428 462332 40492
rect 154068 40020 154132 40084
rect 183508 40156 183572 40220
rect 219388 40080 219452 40084
rect 249748 40292 249812 40356
rect 219388 40024 219402 40080
rect 219402 40024 219452 40080
rect 183508 39884 183572 39948
rect 219388 40020 219452 40024
rect 462268 40156 462332 40220
rect 249748 39884 249812 39948
rect 219388 39748 219452 39812
rect 307892 38660 307956 38724
rect 462268 17036 462332 17100
rect 151676 16628 151740 16692
rect 462268 16764 462332 16828
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 547136 149004 581498
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 151859 548588 151925 548589
rect 151859 548524 151860 548588
rect 151924 548524 151925 548588
rect 151859 548523 151925 548524
rect 151675 544644 151741 544645
rect 151675 544580 151676 544644
rect 151740 544580 151741 544644
rect 151675 544579 151741 544580
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 151678 534170 151738 544579
rect 151494 534110 151738 534170
rect 151494 512005 151554 534110
rect 150755 512004 150821 512005
rect 150755 511940 150756 512004
rect 150820 511940 150821 512004
rect 150755 511939 150821 511940
rect 151491 512004 151557 512005
rect 151491 511940 151492 512004
rect 151556 511940 151557 512004
rect 151491 511939 151557 511940
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 150758 502621 150818 511939
rect 150755 502620 150821 502621
rect 150755 502556 150756 502620
rect 150820 502556 150821 502620
rect 150755 502555 150821 502556
rect 151123 502484 151189 502485
rect 151123 502420 151124 502484
rect 151188 502420 151189 502484
rect 151123 502419 151189 502420
rect 151126 495410 151186 502419
rect 151126 495350 151370 495410
rect 151310 485210 151370 495350
rect 151310 485150 151554 485210
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 151494 456925 151554 485150
rect 151491 456924 151557 456925
rect 151491 456860 151492 456924
rect 151556 456860 151557 456924
rect 151491 456859 151557 456860
rect 151307 456652 151373 456653
rect 151307 456588 151308 456652
rect 151372 456588 151373 456652
rect 151307 456587 151373 456588
rect 151310 447269 151370 456587
rect 151307 447268 151373 447269
rect 151307 447204 151308 447268
rect 151372 447204 151373 447268
rect 151307 447203 151373 447204
rect 151491 446996 151557 446997
rect 151491 446932 151492 446996
rect 151556 446932 151557 446996
rect 151491 446931 151557 446932
rect 151494 441557 151554 446931
rect 151491 441556 151557 441557
rect 151491 441492 151492 441556
rect 151556 441492 151557 441556
rect 151491 441491 151557 441492
rect 150939 441420 151005 441421
rect 150939 441356 150940 441420
rect 151004 441356 151005 441420
rect 150939 441355 151005 441356
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 150942 432037 151002 441355
rect 150939 432036 151005 432037
rect 150939 431972 150940 432036
rect 151004 431972 151005 432036
rect 150939 431971 151005 431972
rect 151675 432036 151741 432037
rect 151675 431972 151676 432036
rect 151740 431972 151741 432036
rect 151675 431971 151741 431972
rect 151678 427957 151738 431971
rect 151675 427956 151741 427957
rect 151675 427892 151676 427956
rect 151740 427892 151741 427956
rect 151675 427891 151741 427892
rect 151675 427820 151741 427821
rect 151675 427756 151676 427820
rect 151740 427756 151741 427820
rect 151675 427755 151741 427756
rect 151678 423741 151738 427755
rect 151675 423740 151741 423741
rect 151675 423676 151676 423740
rect 151740 423676 151741 423740
rect 151675 423675 151741 423676
rect 151675 423604 151741 423605
rect 151675 423540 151676 423604
rect 151740 423540 151741 423604
rect 151675 423539 151741 423540
rect 151678 417890 151738 423539
rect 151310 417830 151738 417890
rect 151310 412589 151370 417830
rect 151307 412588 151373 412589
rect 151307 412524 151308 412588
rect 151372 412524 151373 412588
rect 151307 412523 151373 412524
rect 151491 412452 151557 412453
rect 151491 412388 151492 412452
rect 151556 412388 151557 412452
rect 151491 412387 151557 412388
rect 151494 402933 151554 412387
rect 151491 402932 151557 402933
rect 151491 402868 151492 402932
rect 151556 402868 151557 402932
rect 151491 402867 151557 402868
rect 151123 402796 151189 402797
rect 151123 402732 151124 402796
rect 151188 402732 151189 402796
rect 151123 402731 151189 402732
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 151126 393413 151186 402731
rect 151123 393412 151189 393413
rect 151123 393348 151124 393412
rect 151188 393348 151189 393412
rect 151123 393347 151189 393348
rect 151675 393412 151741 393413
rect 151675 393348 151676 393412
rect 151740 393348 151741 393412
rect 151675 393347 151741 393348
rect 151678 389333 151738 393347
rect 151675 389332 151741 389333
rect 151675 389268 151676 389332
rect 151740 389268 151741 389332
rect 151675 389267 151741 389268
rect 151491 389060 151557 389061
rect 151491 388996 151492 389060
rect 151556 388996 151557 389060
rect 151491 388995 151557 388996
rect 151494 364445 151554 388995
rect 151491 364444 151557 364445
rect 151491 364380 151492 364444
rect 151556 364380 151557 364444
rect 151491 364379 151557 364380
rect 151675 364444 151741 364445
rect 151675 364380 151676 364444
rect 151740 364380 151741 364444
rect 151675 364379 151741 364380
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 151678 356285 151738 364379
rect 151675 356284 151741 356285
rect 151675 356220 151676 356284
rect 151740 356220 151741 356284
rect 151675 356219 151741 356220
rect 151491 356148 151557 356149
rect 151491 356084 151492 356148
rect 151556 356084 151557 356148
rect 151491 356083 151557 356084
rect 151494 348533 151554 356083
rect 151491 348532 151557 348533
rect 151491 348468 151492 348532
rect 151556 348468 151557 348532
rect 151491 348467 151557 348468
rect 151862 346629 151922 548523
rect 152004 547136 152604 549098
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 152779 548860 152845 548861
rect 152779 548796 152780 548860
rect 152844 548796 152845 548860
rect 152779 548795 152845 548796
rect 152227 545324 152293 545325
rect 152227 545260 152228 545324
rect 152292 545260 152293 545324
rect 152227 545259 152293 545260
rect 152230 536213 152290 545259
rect 152782 539610 152842 548795
rect 155604 547136 156204 552698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 547136 163404 559898
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 547136 167004 563498
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 547136 170604 567098
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 547136 174204 570698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 547136 181404 577898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 547136 185004 581498
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 547136 188604 549098
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 547136 192204 552698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 547136 199404 559898
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 547136 203004 563498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 547136 206604 567098
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 547136 210204 570698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 547136 217404 577898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 547136 221004 581498
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 547136 224604 549098
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 547136 228204 552698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 547136 235404 559898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 547136 239004 563498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 547136 242604 567098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 547136 246204 570698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 547136 253404 577898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 547136 257004 581498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 547136 260604 549098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 547136 264204 552698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 547136 271404 559898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 547136 275004 563498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 547136 278604 567098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 547136 282204 570698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 547136 289404 577898
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 547136 293004 581498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 547136 296604 549098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 547136 300204 552698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 547136 307404 559898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 547136 311004 563498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 547136 314604 567098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 547136 318204 570698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 547136 325404 577898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 547136 329004 581498
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 547136 332604 549098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 547136 336204 552698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 547136 343404 559898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 547136 347004 563498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 547136 350604 567098
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 547136 354204 570698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 547136 361404 577898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 547136 365004 581498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 547136 368604 549098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 547136 372204 552698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 547136 379404 559898
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 547136 383004 563498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 547136 386604 567098
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 547136 390204 570698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 547136 397404 577898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 547136 401004 581498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 547136 404604 549098
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 547136 408204 552698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 547136 415404 559898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 547136 419004 563498
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 547136 422604 567098
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 547136 426204 570698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 547136 433404 577898
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 547136 437004 581498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 547136 440604 549098
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 547136 444204 552698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 447731 549132 447797 549133
rect 447731 549068 447732 549132
rect 447796 549068 447797 549132
rect 447731 549067 447797 549068
rect 446627 548996 446693 548997
rect 446627 548932 446628 548996
rect 446692 548932 446693 548996
rect 446627 548931 446693 548932
rect 446443 548724 446509 548725
rect 446443 548660 446444 548724
rect 446508 548660 446509 548724
rect 446443 548659 446509 548660
rect 152963 545188 153029 545189
rect 152963 545124 152964 545188
rect 153028 545124 153029 545188
rect 152963 545123 153029 545124
rect 152414 539550 152842 539610
rect 152227 536212 152293 536213
rect 152227 536148 152228 536212
rect 152292 536148 152293 536212
rect 152227 536147 152293 536148
rect 152043 520164 152109 520165
rect 152043 520100 152044 520164
rect 152108 520100 152109 520164
rect 152043 520099 152109 520100
rect 152046 510645 152106 520099
rect 152043 510644 152109 510645
rect 152043 510580 152044 510644
rect 152108 510580 152109 510644
rect 152043 510579 152109 510580
rect 152043 490924 152109 490925
rect 152043 490860 152044 490924
rect 152108 490860 152109 490924
rect 152043 490859 152109 490860
rect 152046 481677 152106 490859
rect 152043 481676 152109 481677
rect 152043 481612 152044 481676
rect 152108 481612 152109 481676
rect 152043 481611 152109 481612
rect 152227 481540 152293 481541
rect 152227 481476 152228 481540
rect 152292 481476 152293 481540
rect 152227 481475 152293 481476
rect 152230 472021 152290 481475
rect 152227 472020 152293 472021
rect 152227 471956 152228 472020
rect 152292 471956 152293 472020
rect 152227 471955 152293 471956
rect 152227 452572 152293 452573
rect 152227 452508 152228 452572
rect 152292 452508 152293 452572
rect 152227 452507 152293 452508
rect 152230 443189 152290 452507
rect 152227 443188 152293 443189
rect 152227 443124 152228 443188
rect 152292 443124 152293 443188
rect 152227 443123 152293 443124
rect 152227 423604 152293 423605
rect 152227 423540 152228 423604
rect 152292 423540 152293 423604
rect 152227 423539 152293 423540
rect 152230 414221 152290 423539
rect 152227 414220 152293 414221
rect 152227 414156 152228 414220
rect 152292 414156 152293 414220
rect 152227 414155 152293 414156
rect 152227 404292 152293 404293
rect 152227 404228 152228 404292
rect 152292 404228 152293 404292
rect 152227 404227 152293 404228
rect 152230 394909 152290 404227
rect 152227 394908 152293 394909
rect 152227 394844 152228 394908
rect 152292 394844 152293 394908
rect 152227 394843 152293 394844
rect 152227 365668 152293 365669
rect 152227 365604 152228 365668
rect 152292 365604 152293 365668
rect 152227 365603 152293 365604
rect 152230 356285 152290 365603
rect 152227 356284 152293 356285
rect 152227 356220 152228 356284
rect 152292 356220 152293 356284
rect 152227 356219 152293 356220
rect 152227 348532 152293 348533
rect 152227 348468 152228 348532
rect 152292 348468 152293 348532
rect 152227 348467 152293 348468
rect 151859 346628 151925 346629
rect 151859 346564 151860 346628
rect 151924 346564 151925 346628
rect 151859 346563 151925 346564
rect 151859 346220 151925 346221
rect 151859 346156 151860 346220
rect 151924 346156 151925 346220
rect 151859 346155 151925 346156
rect 151862 335341 151922 346155
rect 152230 335477 152290 348467
rect 152043 335476 152109 335477
rect 152043 335412 152044 335476
rect 152108 335412 152109 335476
rect 152043 335411 152109 335412
rect 152227 335476 152293 335477
rect 152227 335412 152228 335476
rect 152292 335412 152293 335476
rect 152227 335411 152293 335412
rect 151859 335340 151925 335341
rect 151859 335276 151860 335340
rect 151924 335276 151925 335340
rect 151859 335275 151925 335276
rect 152046 335205 152106 335411
rect 152043 335204 152109 335205
rect 152043 335140 152044 335204
rect 152108 335140 152109 335204
rect 152043 335139 152109 335140
rect 152227 335204 152293 335205
rect 152227 335140 152228 335204
rect 152292 335140 152293 335204
rect 152227 335139 152293 335140
rect 151859 334116 151925 334117
rect 151859 334052 151860 334116
rect 151924 334052 151925 334116
rect 151859 334051 151925 334052
rect 151862 327453 151922 334051
rect 151859 327452 151925 327453
rect 151859 327388 151860 327452
rect 151924 327388 151925 327452
rect 151859 327387 151925 327388
rect 151491 327180 151557 327181
rect 151491 327116 151492 327180
rect 151556 327116 151557 327180
rect 152230 327178 152290 335139
rect 151491 327115 151557 327116
rect 151862 327118 152290 327178
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 151494 325685 151554 327115
rect 150755 325684 150821 325685
rect 150755 325620 150756 325684
rect 150820 325620 150821 325684
rect 150755 325619 150821 325620
rect 151491 325684 151557 325685
rect 151491 325620 151492 325684
rect 151556 325620 151557 325684
rect 151491 325619 151557 325620
rect 150758 316301 150818 325619
rect 150755 316300 150821 316301
rect 150755 316236 150756 316300
rect 150820 316236 150821 316300
rect 150755 316235 150821 316236
rect 151307 316300 151373 316301
rect 151307 316236 151308 316300
rect 151372 316236 151373 316300
rect 151307 316235 151373 316236
rect 151310 316029 151370 316235
rect 151307 316028 151373 316029
rect 151307 315964 151308 316028
rect 151372 315964 151373 316028
rect 151307 315963 151373 315964
rect 151491 316028 151557 316029
rect 151491 315964 151492 316028
rect 151556 315964 151557 316028
rect 151491 315963 151557 315964
rect 151494 314669 151554 315963
rect 151307 314668 151373 314669
rect 151307 314604 151308 314668
rect 151372 314604 151373 314668
rect 151307 314603 151373 314604
rect 151491 314668 151557 314669
rect 151491 314604 151492 314668
rect 151556 314604 151557 314668
rect 151491 314603 151557 314604
rect 151310 305013 151370 314603
rect 151123 305012 151189 305013
rect 151123 304948 151124 305012
rect 151188 304948 151189 305012
rect 151123 304947 151189 304948
rect 151307 305012 151373 305013
rect 151307 304948 151308 305012
rect 151372 304948 151373 305012
rect 151307 304947 151373 304948
rect 151126 296853 151186 304947
rect 151123 296852 151189 296853
rect 151123 296788 151124 296852
rect 151188 296788 151189 296852
rect 151123 296787 151189 296788
rect 151675 296852 151741 296853
rect 151675 296788 151676 296852
rect 151740 296788 151741 296852
rect 151675 296787 151741 296788
rect 151678 292773 151738 296787
rect 151675 292772 151741 292773
rect 151675 292708 151676 292772
rect 151740 292708 151741 292772
rect 151675 292707 151741 292708
rect 151491 292500 151557 292501
rect 151491 292436 151492 292500
rect 151556 292436 151557 292500
rect 151491 292435 151557 292436
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 151494 280805 151554 292435
rect 151123 280804 151189 280805
rect 151123 280740 151124 280804
rect 151188 280740 151189 280804
rect 151123 280739 151189 280740
rect 151491 280804 151557 280805
rect 151491 280740 151492 280804
rect 151556 280740 151557 280804
rect 151491 280739 151557 280740
rect 151126 276045 151186 280739
rect 151123 276044 151189 276045
rect 151123 275980 151124 276044
rect 151188 275980 151189 276044
rect 151123 275979 151189 275980
rect 151491 276044 151557 276045
rect 151491 275980 151492 276044
rect 151556 275980 151557 276044
rect 151491 275979 151557 275980
rect 151494 266253 151554 275979
rect 151123 266252 151189 266253
rect 151123 266188 151124 266252
rect 151188 266188 151189 266252
rect 151123 266187 151189 266188
rect 151491 266252 151557 266253
rect 151491 266188 151492 266252
rect 151556 266188 151557 266252
rect 151491 266187 151557 266188
rect 151126 256733 151186 266187
rect 151123 256732 151189 256733
rect 151123 256668 151124 256732
rect 151188 256668 151189 256732
rect 151123 256667 151189 256668
rect 151491 256732 151557 256733
rect 151491 256668 151492 256732
rect 151556 256668 151557 256732
rect 151491 256667 151557 256668
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 151494 246941 151554 256667
rect 151123 246940 151189 246941
rect 151123 246876 151124 246940
rect 151188 246876 151189 246940
rect 151123 246875 151189 246876
rect 151491 246940 151557 246941
rect 151491 246876 151492 246940
rect 151556 246876 151557 246940
rect 151491 246875 151557 246876
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 222054 149004 243136
rect 151126 237421 151186 246875
rect 151123 237420 151189 237421
rect 151123 237356 151124 237420
rect 151188 237356 151189 237420
rect 151123 237355 151189 237356
rect 151491 237420 151557 237421
rect 151491 237356 151492 237420
rect 151556 237356 151557 237420
rect 151491 237355 151557 237356
rect 151494 237285 151554 237355
rect 151491 237284 151557 237285
rect 151491 237220 151492 237284
rect 151556 237220 151557 237284
rect 151491 237219 151557 237220
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 151491 220964 151557 220965
rect 151491 220900 151492 220964
rect 151556 220900 151557 220964
rect 151491 220899 151557 220900
rect 151494 212533 151554 220899
rect 151491 212532 151557 212533
rect 151491 212468 151492 212532
rect 151556 212468 151557 212532
rect 151491 212467 151557 212468
rect 151307 212396 151373 212397
rect 151307 212332 151308 212396
rect 151372 212332 151373 212396
rect 151307 212331 151373 212332
rect 151310 206277 151370 212331
rect 151307 206276 151373 206277
rect 151307 206212 151308 206276
rect 151372 206212 151373 206276
rect 151307 206211 151373 206212
rect 151862 201381 151922 327118
rect 152227 327044 152293 327045
rect 152227 326980 152228 327044
rect 152292 326980 152293 327044
rect 152227 326979 152293 326980
rect 152230 317661 152290 326979
rect 152227 317660 152293 317661
rect 152227 317596 152228 317660
rect 152292 317596 152293 317660
rect 152227 317595 152293 317596
rect 152227 307732 152293 307733
rect 152227 307668 152228 307732
rect 152292 307668 152293 307732
rect 152227 307667 152293 307668
rect 152230 298349 152290 307667
rect 152227 298348 152293 298349
rect 152227 298284 152228 298348
rect 152292 298284 152293 298348
rect 152227 298283 152293 298284
rect 152227 288420 152293 288421
rect 152227 288356 152228 288420
rect 152292 288356 152293 288420
rect 152227 288355 152293 288356
rect 152230 279037 152290 288355
rect 152227 279036 152293 279037
rect 152227 278972 152228 279036
rect 152292 278972 152293 279036
rect 152227 278971 152293 278972
rect 152414 243810 152474 539550
rect 152966 537570 153026 545123
rect 154067 544644 154133 544645
rect 154067 544580 154068 544644
rect 154132 544580 154133 544644
rect 154067 544579 154133 544580
rect 203195 544644 203261 544645
rect 203195 544580 203196 544644
rect 203260 544580 203261 544644
rect 203195 544579 203261 544580
rect 205403 544644 205469 544645
rect 205403 544580 205404 544644
rect 205468 544580 205469 544644
rect 205403 544579 205469 544580
rect 208163 544644 208229 544645
rect 208163 544580 208164 544644
rect 208228 544580 208229 544644
rect 208163 544579 208229 544580
rect 213499 544644 213565 544645
rect 213499 544580 213500 544644
rect 213564 544580 213565 544644
rect 213499 544579 213565 544580
rect 221411 544644 221477 544645
rect 221411 544580 221412 544644
rect 221476 544580 221477 544644
rect 221411 544579 221477 544580
rect 231531 544644 231597 544645
rect 231531 544580 231532 544644
rect 231596 544580 231597 544644
rect 231531 544579 231597 544580
rect 386459 544644 386525 544645
rect 386459 544580 386460 544644
rect 386524 544580 386525 544644
rect 386459 544579 386525 544580
rect 152598 537510 153026 537570
rect 152598 531450 152658 537510
rect 152963 536212 153029 536213
rect 152963 536148 152964 536212
rect 153028 536148 153029 536212
rect 152963 536147 153029 536148
rect 152598 531390 152842 531450
rect 152782 521661 152842 531390
rect 152779 521660 152845 521661
rect 152779 521596 152780 521660
rect 152844 521596 152845 521660
rect 152779 521595 152845 521596
rect 152595 520300 152661 520301
rect 152595 520236 152596 520300
rect 152660 520236 152661 520300
rect 152595 520235 152661 520236
rect 152598 520165 152658 520235
rect 152595 520164 152661 520165
rect 152595 520100 152596 520164
rect 152660 520100 152661 520164
rect 152595 520099 152661 520100
rect 152779 510644 152845 510645
rect 152779 510580 152780 510644
rect 152844 510580 152845 510644
rect 152779 510579 152845 510580
rect 152782 500850 152842 510579
rect 152966 510509 153026 536147
rect 152963 510508 153029 510509
rect 152963 510444 152964 510508
rect 153028 510444 153029 510508
rect 152963 510443 153029 510444
rect 152963 510100 153029 510101
rect 152963 510036 152964 510100
rect 153028 510036 153029 510100
rect 152963 510035 153029 510036
rect 152598 500790 152842 500850
rect 152598 491469 152658 500790
rect 152595 491468 152661 491469
rect 152595 491404 152596 491468
rect 152660 491404 152661 491468
rect 152595 491403 152661 491404
rect 152779 491332 152845 491333
rect 152779 491268 152780 491332
rect 152844 491268 152845 491332
rect 152779 491267 152845 491268
rect 152782 491197 152842 491267
rect 152779 491196 152845 491197
rect 152779 491132 152780 491196
rect 152844 491132 152845 491196
rect 152779 491131 152845 491132
rect 152779 481676 152845 481677
rect 152779 481612 152780 481676
rect 152844 481612 152845 481676
rect 152779 481611 152845 481612
rect 152782 481541 152842 481611
rect 152779 481540 152845 481541
rect 152779 481476 152780 481540
rect 152844 481476 152845 481540
rect 152779 481475 152845 481476
rect 152779 472020 152845 472021
rect 152779 471956 152780 472020
rect 152844 471956 152845 472020
rect 152779 471955 152845 471956
rect 152782 463589 152842 471955
rect 152779 463588 152845 463589
rect 152779 463524 152780 463588
rect 152844 463524 152845 463588
rect 152779 463523 152845 463524
rect 152779 454204 152845 454205
rect 152779 454140 152780 454204
rect 152844 454140 152845 454204
rect 152779 454139 152845 454140
rect 152782 452573 152842 454139
rect 152779 452572 152845 452573
rect 152779 452508 152780 452572
rect 152844 452508 152845 452572
rect 152779 452507 152845 452508
rect 152595 443052 152661 443053
rect 152595 442988 152596 443052
rect 152660 443050 152661 443052
rect 152660 442990 152842 443050
rect 152660 442988 152661 442990
rect 152595 442987 152661 442988
rect 152782 423605 152842 442990
rect 152779 423604 152845 423605
rect 152779 423540 152780 423604
rect 152844 423540 152845 423604
rect 152779 423539 152845 423540
rect 152779 414084 152845 414085
rect 152779 414020 152780 414084
rect 152844 414020 152845 414084
rect 152779 414019 152845 414020
rect 152782 404293 152842 414019
rect 152779 404292 152845 404293
rect 152779 404228 152780 404292
rect 152844 404228 152845 404292
rect 152779 404227 152845 404228
rect 152779 394772 152845 394773
rect 152779 394708 152780 394772
rect 152844 394708 152845 394772
rect 152779 394707 152845 394708
rect 152782 365669 152842 394707
rect 152779 365668 152845 365669
rect 152779 365604 152780 365668
rect 152844 365604 152845 365668
rect 152779 365603 152845 365604
rect 152779 356148 152845 356149
rect 152779 356084 152780 356148
rect 152844 356084 152845 356148
rect 152779 356083 152845 356084
rect 152782 327589 152842 356083
rect 152966 327589 153026 510035
rect 153147 463588 153213 463589
rect 153147 463524 153148 463588
rect 153212 463524 153213 463588
rect 153147 463523 153213 463524
rect 153150 454205 153210 463523
rect 153147 454204 153213 454205
rect 153147 454140 153148 454204
rect 153212 454140 153213 454204
rect 153147 454139 153213 454140
rect 152779 327588 152845 327589
rect 152779 327524 152780 327588
rect 152844 327524 152845 327588
rect 152779 327523 152845 327524
rect 152963 327588 153029 327589
rect 152963 327524 152964 327588
rect 153028 327524 153029 327588
rect 152963 327523 153029 327524
rect 152779 327180 152845 327181
rect 152779 327116 152780 327180
rect 152844 327116 152845 327180
rect 152779 327115 152845 327116
rect 152963 327180 153029 327181
rect 152963 327116 152964 327180
rect 153028 327116 153029 327180
rect 152963 327115 153029 327116
rect 152782 327045 152842 327115
rect 152779 327044 152845 327045
rect 152779 326980 152780 327044
rect 152844 326980 152845 327044
rect 152779 326979 152845 326980
rect 152779 317524 152845 317525
rect 152779 317460 152780 317524
rect 152844 317460 152845 317524
rect 152779 317459 152845 317460
rect 152782 307733 152842 317459
rect 152779 307732 152845 307733
rect 152779 307668 152780 307732
rect 152844 307668 152845 307732
rect 152779 307667 152845 307668
rect 152779 298212 152845 298213
rect 152779 298148 152780 298212
rect 152844 298148 152845 298212
rect 152779 298147 152845 298148
rect 152782 288421 152842 298147
rect 152779 288420 152845 288421
rect 152779 288356 152780 288420
rect 152844 288356 152845 288420
rect 152779 288355 152845 288356
rect 152779 278900 152845 278901
rect 152779 278836 152780 278900
rect 152844 278836 152845 278900
rect 152779 278835 152845 278836
rect 152782 259453 152842 278835
rect 152779 259452 152845 259453
rect 152779 259388 152780 259452
rect 152844 259388 152845 259452
rect 152779 259387 152845 259388
rect 152595 259316 152661 259317
rect 152595 259252 152596 259316
rect 152660 259252 152661 259316
rect 152595 259251 152661 259252
rect 152598 248573 152658 259251
rect 152595 248572 152661 248573
rect 152595 248508 152596 248572
rect 152660 248508 152661 248572
rect 152595 248507 152661 248508
rect 152779 248436 152845 248437
rect 152779 248372 152780 248436
rect 152844 248372 152845 248436
rect 152779 248371 152845 248372
rect 152782 248301 152842 248371
rect 152779 248300 152845 248301
rect 152779 248236 152780 248300
rect 152844 248236 152845 248300
rect 152779 248235 152845 248236
rect 152966 244493 153026 327115
rect 153515 248300 153581 248301
rect 153515 248236 153516 248300
rect 153580 248236 153581 248300
rect 153515 248235 153581 248236
rect 152963 244492 153029 244493
rect 152963 244428 152964 244492
rect 153028 244428 153029 244492
rect 152963 244427 153029 244428
rect 152963 244220 153029 244221
rect 152963 244156 152964 244220
rect 153028 244156 153029 244220
rect 152963 244155 153029 244156
rect 152414 243750 152842 243810
rect 152004 225654 152604 243136
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 151859 201380 151925 201381
rect 151859 201316 151860 201380
rect 151924 201316 151925 201380
rect 151859 201315 151925 201316
rect 151859 196620 151925 196621
rect 151859 196556 151860 196620
rect 151924 196556 151925 196620
rect 151859 196555 151925 196556
rect 151675 193220 151741 193221
rect 151675 193156 151676 193220
rect 151740 193156 151741 193220
rect 151675 193155 151741 193156
rect 151678 188050 151738 193155
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 151310 187990 151738 188050
rect 151310 177309 151370 187990
rect 151307 177308 151373 177309
rect 151307 177244 151308 177308
rect 151372 177244 151373 177308
rect 151307 177243 151373 177244
rect 151862 165613 151922 196555
rect 152004 189654 152604 225098
rect 152782 215253 152842 243750
rect 152779 215252 152845 215253
rect 152779 215188 152780 215252
rect 152844 215188 152845 215252
rect 152779 215187 152845 215188
rect 152779 215116 152845 215117
rect 152779 215052 152780 215116
rect 152844 215052 152845 215116
rect 152779 215051 152845 215052
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 151859 165612 151925 165613
rect 151859 165548 151860 165612
rect 151924 165548 151925 165612
rect 151859 165547 151925 165548
rect 151123 165476 151189 165477
rect 151123 165412 151124 165476
rect 151188 165412 151189 165476
rect 151123 165411 151189 165412
rect 151126 156637 151186 165411
rect 151123 156636 151189 156637
rect 151123 156572 151124 156636
rect 151188 156572 151189 156636
rect 151123 156571 151189 156572
rect 151491 156636 151557 156637
rect 151491 156572 151492 156636
rect 151556 156572 151557 156636
rect 151491 156571 151557 156572
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 151494 147797 151554 156571
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 151491 147796 151557 147797
rect 151491 147732 151492 147796
rect 151556 147732 151557 147796
rect 151491 147731 151557 147732
rect 151307 147524 151373 147525
rect 151307 147460 151308 147524
rect 151372 147460 151373 147524
rect 151307 147459 151373 147460
rect 151310 114749 151370 147459
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 151307 114748 151373 114749
rect 151307 114684 151308 114748
rect 151372 114684 151373 114748
rect 151307 114683 151373 114684
rect 151491 114612 151557 114613
rect 151491 114548 151492 114612
rect 151556 114548 151557 114612
rect 151491 114547 151557 114548
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 151494 113117 151554 114547
rect 151491 113116 151557 113117
rect 151491 113052 151492 113116
rect 151556 113052 151557 113116
rect 151491 113051 151557 113052
rect 151307 104276 151373 104277
rect 151307 104212 151308 104276
rect 151372 104212 151373 104276
rect 151307 104211 151373 104212
rect 151310 92853 151370 104211
rect 151307 92852 151373 92853
rect 151307 92788 151308 92852
rect 151372 92788 151373 92852
rect 151307 92787 151373 92788
rect 150939 91220 151005 91221
rect 150939 91156 150940 91220
rect 151004 91156 151005 91220
rect 150939 91155 151005 91156
rect 150942 83061 151002 91155
rect 150939 83060 151005 83061
rect 150939 82996 150940 83060
rect 151004 82996 151005 83060
rect 150939 82995 151005 82996
rect 151307 82924 151373 82925
rect 151307 82860 151308 82924
rect 151372 82860 151373 82924
rect 151307 82859 151373 82860
rect 151310 81429 151370 82859
rect 152004 81654 152604 117098
rect 151307 81428 151373 81429
rect 151307 81364 151308 81428
rect 151372 81364 151373 81428
rect 151307 81363 151373 81364
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 151491 71908 151557 71909
rect 151491 71844 151492 71908
rect 151556 71844 151557 71908
rect 151491 71843 151557 71844
rect 151494 69730 151554 71843
rect 151310 69670 151554 69730
rect 151310 55861 151370 69670
rect 151307 55860 151373 55861
rect 151307 55796 151308 55860
rect 151372 55796 151373 55860
rect 151307 55795 151373 55796
rect 151675 55860 151741 55861
rect 151675 55796 151676 55860
rect 151740 55796 151741 55860
rect 151675 55795 151741 55796
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 151678 33010 151738 55795
rect 152004 45654 152604 81098
rect 152782 80069 152842 215051
rect 152966 122773 153026 244155
rect 153518 238781 153578 248235
rect 153147 238780 153213 238781
rect 153147 238716 153148 238780
rect 153212 238716 153213 238780
rect 153147 238715 153213 238716
rect 153515 238780 153581 238781
rect 153515 238716 153516 238780
rect 153580 238716 153581 238780
rect 153515 238715 153581 238716
rect 153150 222325 153210 238715
rect 153147 222324 153213 222325
rect 153147 222260 153148 222324
rect 153212 222260 153213 222324
rect 153147 222259 153213 222260
rect 153331 222052 153397 222053
rect 153331 221988 153332 222052
rect 153396 221988 153397 222052
rect 153331 221987 153397 221988
rect 153334 220690 153394 221987
rect 153150 220630 153394 220690
rect 153150 215117 153210 220630
rect 153147 215116 153213 215117
rect 153147 215052 153148 215116
rect 153212 215052 153213 215116
rect 153147 215051 153213 215052
rect 152963 122772 153029 122773
rect 152963 122708 152964 122772
rect 153028 122708 153029 122772
rect 152963 122707 153029 122708
rect 152779 80068 152845 80069
rect 152779 80004 152780 80068
rect 152844 80004 152845 80068
rect 152779 80003 152845 80004
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 151678 32950 151922 33010
rect 151862 23490 151922 32950
rect 151678 23430 151922 23490
rect 151678 16693 151738 23430
rect 151675 16692 151741 16693
rect 151675 16628 151676 16692
rect 151740 16628 151741 16692
rect 151675 16627 151741 16628
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 9654 152604 45098
rect 154070 40085 154130 544579
rect 203198 543149 203258 544579
rect 205406 543285 205466 544579
rect 208166 543421 208226 544579
rect 213502 543557 213562 544579
rect 221414 543693 221474 544579
rect 226931 543964 226997 543965
rect 226931 543900 226932 543964
rect 226996 543900 226997 543964
rect 226931 543899 226997 543900
rect 221411 543692 221477 543693
rect 221411 543628 221412 543692
rect 221476 543628 221477 543692
rect 221411 543627 221477 543628
rect 213499 543556 213565 543557
rect 213499 543492 213500 543556
rect 213564 543492 213565 543556
rect 213499 543491 213565 543492
rect 208163 543420 208229 543421
rect 208163 543356 208164 543420
rect 208228 543356 208229 543420
rect 208163 543355 208229 543356
rect 226934 543285 226994 543899
rect 231534 543285 231594 544579
rect 231715 543964 231781 543965
rect 231715 543900 231716 543964
rect 231780 543900 231781 543964
rect 231715 543899 231781 543900
rect 231718 543285 231778 543899
rect 205403 543284 205469 543285
rect 205403 543220 205404 543284
rect 205468 543220 205469 543284
rect 205403 543219 205469 543220
rect 226931 543284 226997 543285
rect 226931 543220 226932 543284
rect 226996 543220 226997 543284
rect 226931 543219 226997 543220
rect 231531 543284 231597 543285
rect 231531 543220 231532 543284
rect 231596 543220 231597 543284
rect 231531 543219 231597 543220
rect 231715 543284 231781 543285
rect 231715 543220 231716 543284
rect 231780 543220 231781 543284
rect 231715 543219 231781 543220
rect 203195 543148 203261 543149
rect 203195 543084 203196 543148
rect 203260 543084 203261 543148
rect 203195 543083 203261 543084
rect 231163 543148 231229 543149
rect 231163 543084 231164 543148
rect 231228 543084 231229 543148
rect 231163 543083 231229 543084
rect 231899 543148 231965 543149
rect 231899 543084 231900 543148
rect 231964 543084 231965 543148
rect 231899 543083 231965 543084
rect 231166 542874 231226 543083
rect 231347 543012 231413 543013
rect 231347 542948 231348 543012
rect 231412 543010 231413 543012
rect 231715 543012 231781 543013
rect 231715 543010 231716 543012
rect 231412 542950 231716 543010
rect 231412 542948 231413 542950
rect 231347 542947 231413 542948
rect 231715 542948 231716 542950
rect 231780 542948 231781 543012
rect 231715 542947 231781 542948
rect 231902 542874 231962 543083
rect 386462 543013 386522 544579
rect 386459 543012 386525 543013
rect 386459 542948 386460 543012
rect 386524 542948 386525 543012
rect 386459 542947 386525 542948
rect 231166 542814 231962 542874
rect 446446 254690 446506 548659
rect 446630 298485 446690 548931
rect 447734 357781 447794 549067
rect 450804 547136 451404 559898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 447731 357780 447797 357781
rect 447731 357716 447732 357780
rect 447796 357716 447797 357780
rect 447731 357715 447797 357716
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 446627 298484 446693 298485
rect 446627 298420 446628 298484
rect 446692 298420 446693 298484
rect 446627 298419 446693 298420
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 446446 254630 446874 254690
rect 446814 251565 446874 254630
rect 446811 251564 446877 251565
rect 446811 251500 446812 251564
rect 446876 251500 446877 251564
rect 446811 251499 446877 251500
rect 155604 229254 156204 243136
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 154067 40084 154133 40085
rect 154067 40020 154068 40084
rect 154132 40020 154133 40084
rect 154067 40019 154133 40020
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 236454 163404 243136
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 240054 167004 243136
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 207654 170604 243136
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 211254 174204 243136
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 218454 181404 243136
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 184404 222054 185004 243136
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 183507 40220 183573 40221
rect 183507 40156 183508 40220
rect 183572 40156 183573 40220
rect 183507 40155 183573 40156
rect 183510 39949 183570 40155
rect 183507 39948 183573 39949
rect 183507 39884 183508 39948
rect 183572 39884 183573 39948
rect 183507 39883 183573 39884
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 225654 188604 243136
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 191604 229254 192204 243136
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 189027 104820 189093 104821
rect 189027 104756 189028 104820
rect 189092 104756 189093 104820
rect 189027 104755 189093 104756
rect 189030 95301 189090 104755
rect 189027 95300 189093 95301
rect 189027 95236 189028 95300
rect 189092 95236 189093 95300
rect 189027 95235 189093 95236
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 236454 199404 243136
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 240054 203004 243136
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 207654 206604 243136
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 211254 210204 243136
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 218454 217404 243136
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 220404 222054 221004 243136
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 219387 40084 219453 40085
rect 219387 40020 219388 40084
rect 219452 40020 219453 40084
rect 219387 40019 219453 40020
rect 219390 39813 219450 40019
rect 219387 39812 219453 39813
rect 219387 39748 219388 39812
rect 219452 39748 219453 39812
rect 219387 39747 219453 39748
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 225654 224604 243136
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 229254 228204 243136
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 236454 235404 243136
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 240054 239004 243136
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 207654 242604 243136
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 211254 246204 243136
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 252804 218454 253404 243136
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 249747 40356 249813 40357
rect 249747 40292 249748 40356
rect 249812 40292 249813 40356
rect 249747 40291 249813 40292
rect 249750 39949 249810 40291
rect 249747 39948 249813 39949
rect 249747 39884 249748 39948
rect 249812 39884 249813 39948
rect 249747 39883 249813 39884
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 222054 257004 243136
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 225654 260604 243136
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 229254 264204 243136
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 236454 271404 243136
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 240054 275004 243136
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 207654 278604 243136
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 211254 282204 243136
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 218454 289404 243136
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 222054 293004 243136
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 225654 296604 243136
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 229254 300204 243136
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 236454 307404 243136
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 310404 240054 311004 243136
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 307891 48244 307957 48245
rect 307891 48180 307892 48244
rect 307956 48180 307957 48244
rect 307891 48179 307957 48180
rect 307894 38725 307954 48179
rect 307891 38724 307957 38725
rect 307891 38660 307892 38724
rect 307956 38660 307957 38724
rect 307891 38659 307957 38660
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 207654 314604 243136
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 211254 318204 243136
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 218454 325404 243136
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 222054 329004 243136
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 225654 332604 243136
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 229254 336204 243136
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 236454 343404 243136
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 240054 347004 243136
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 207654 350604 243136
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 211254 354204 243136
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 218454 361404 243136
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 222054 365004 243136
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 225654 368604 243136
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 229254 372204 243136
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 236454 379404 243136
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 240054 383004 243136
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 207654 386604 243136
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 211254 390204 243136
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 218454 397404 243136
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 222054 401004 243136
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 225654 404604 243136
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 229254 408204 243136
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 236454 415404 243136
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 240054 419004 243136
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 207654 422604 243136
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 211254 426204 243136
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 218454 433404 243136
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 222054 437004 243136
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 225654 440604 243136
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 229254 444204 243136
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 236454 451404 243136
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 462267 40492 462333 40493
rect 462267 40428 462268 40492
rect 462332 40428 462333 40492
rect 462267 40427 462333 40428
rect 462270 40221 462330 40427
rect 462267 40220 462333 40221
rect 462267 40156 462268 40220
rect 462332 40156 462333 40220
rect 462267 40155 462333 40156
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 462267 17100 462333 17101
rect 462267 17036 462268 17100
rect 462332 17036 462333 17100
rect 462267 17035 462333 17036
rect 462270 16829 462330 17035
rect 462267 16828 462333 16829
rect 462267 16764 462268 16828
rect 462332 16764 462333 16828
rect 462267 16763 462333 16764
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 152186 81418 152422 81654
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 152186 81098 152422 81334
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 147992 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 147992 546054
rect -4756 545734 147992 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 147992 545734
rect -4756 545476 147992 545498
rect 451992 546054 588680 546076
rect 451992 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect 451992 545734 588680 545818
rect 451992 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect 451992 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 147992 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 147992 542454
rect -2916 542134 147992 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 147992 542134
rect -2916 541876 147992 541898
rect 451992 542454 586840 542476
rect 451992 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect 451992 542134 586840 542218
rect 451992 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect 451992 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 147992 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 147992 535254
rect -8436 534934 147992 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 147992 534934
rect -8436 534676 147992 534698
rect 451992 535254 592360 535276
rect 451992 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect 451992 534934 592360 535018
rect 451992 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect 451992 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 147992 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 147992 531654
rect -6596 531334 147992 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 147992 531334
rect -6596 531076 147992 531098
rect 451992 531654 590520 531676
rect 451992 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect 451992 531334 590520 531418
rect 451992 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect 451992 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 147992 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 147992 528054
rect -4756 527734 147992 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 147992 527734
rect -4756 527476 147992 527498
rect 451992 528054 588680 528076
rect 451992 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect 451992 527734 588680 527818
rect 451992 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect 451992 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 147992 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 147992 524454
rect -2916 524134 147992 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 147992 524134
rect -2916 523876 147992 523898
rect 451992 524454 586840 524476
rect 451992 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect 451992 524134 586840 524218
rect 451992 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect 451992 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 147992 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 147992 517254
rect -8436 516934 147992 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 147992 516934
rect -8436 516676 147992 516698
rect 451992 517254 592360 517276
rect 451992 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect 451992 516934 592360 517018
rect 451992 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect 451992 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 147992 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 147992 513654
rect -6596 513334 147992 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 147992 513334
rect -6596 513076 147992 513098
rect 451992 513654 590520 513676
rect 451992 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect 451992 513334 590520 513418
rect 451992 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect 451992 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 147992 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 147992 510054
rect -4756 509734 147992 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 147992 509734
rect -4756 509476 147992 509498
rect 451992 510054 588680 510076
rect 451992 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect 451992 509734 588680 509818
rect 451992 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect 451992 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 147992 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 147992 506454
rect -2916 506134 147992 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 147992 506134
rect -2916 505876 147992 505898
rect 451992 506454 586840 506476
rect 451992 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect 451992 506134 586840 506218
rect 451992 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect 451992 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 147992 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 147992 499254
rect -8436 498934 147992 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 147992 498934
rect -8436 498676 147992 498698
rect 451992 499254 592360 499276
rect 451992 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect 451992 498934 592360 499018
rect 451992 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect 451992 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 147992 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 147992 495654
rect -6596 495334 147992 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 147992 495334
rect -6596 495076 147992 495098
rect 451992 495654 590520 495676
rect 451992 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect 451992 495334 590520 495418
rect 451992 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect 451992 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 147992 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 147992 492054
rect -4756 491734 147992 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 147992 491734
rect -4756 491476 147992 491498
rect 451992 492054 588680 492076
rect 451992 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect 451992 491734 588680 491818
rect 451992 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect 451992 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 147992 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 147992 488454
rect -2916 488134 147992 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 147992 488134
rect -2916 487876 147992 487898
rect 451992 488454 586840 488476
rect 451992 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect 451992 488134 586840 488218
rect 451992 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect 451992 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 147992 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 147992 481254
rect -8436 480934 147992 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 147992 480934
rect -8436 480676 147992 480698
rect 451992 481254 592360 481276
rect 451992 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect 451992 480934 592360 481018
rect 451992 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect 451992 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 147992 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 147992 477654
rect -6596 477334 147992 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 147992 477334
rect -6596 477076 147992 477098
rect 451992 477654 590520 477676
rect 451992 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect 451992 477334 590520 477418
rect 451992 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect 451992 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 147992 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 147992 474054
rect -4756 473734 147992 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 147992 473734
rect -4756 473476 147992 473498
rect 451992 474054 588680 474076
rect 451992 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect 451992 473734 588680 473818
rect 451992 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect 451992 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 147992 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 147992 470454
rect -2916 470134 147992 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 147992 470134
rect -2916 469876 147992 469898
rect 451992 470454 586840 470476
rect 451992 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect 451992 470134 586840 470218
rect 451992 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect 451992 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 147992 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 147992 463254
rect -8436 462934 147992 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 147992 462934
rect -8436 462676 147992 462698
rect 451992 463254 592360 463276
rect 451992 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect 451992 462934 592360 463018
rect 451992 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect 451992 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 147992 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 147992 459654
rect -6596 459334 147992 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 147992 459334
rect -6596 459076 147992 459098
rect 451992 459654 590520 459676
rect 451992 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect 451992 459334 590520 459418
rect 451992 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect 451992 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 147992 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 147992 456054
rect -4756 455734 147992 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 147992 455734
rect -4756 455476 147992 455498
rect 451992 456054 588680 456076
rect 451992 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect 451992 455734 588680 455818
rect 451992 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect 451992 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 147992 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 147992 452454
rect -2916 452134 147992 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 147992 452134
rect -2916 451876 147992 451898
rect 451992 452454 586840 452476
rect 451992 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect 451992 452134 586840 452218
rect 451992 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect 451992 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 147992 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 147992 445254
rect -8436 444934 147992 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 147992 444934
rect -8436 444676 147992 444698
rect 451992 445254 592360 445276
rect 451992 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect 451992 444934 592360 445018
rect 451992 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect 451992 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 147992 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 147992 441654
rect -6596 441334 147992 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 147992 441334
rect -6596 441076 147992 441098
rect 451992 441654 590520 441676
rect 451992 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect 451992 441334 590520 441418
rect 451992 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect 451992 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 147992 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 147992 438054
rect -4756 437734 147992 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 147992 437734
rect -4756 437476 147992 437498
rect 451992 438054 588680 438076
rect 451992 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect 451992 437734 588680 437818
rect 451992 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect 451992 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 147992 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 147992 434454
rect -2916 434134 147992 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 147992 434134
rect -2916 433876 147992 433898
rect 451992 434454 586840 434476
rect 451992 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect 451992 434134 586840 434218
rect 451992 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect 451992 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 147992 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 147992 427254
rect -8436 426934 147992 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 147992 426934
rect -8436 426676 147992 426698
rect 451992 427254 592360 427276
rect 451992 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect 451992 426934 592360 427018
rect 451992 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect 451992 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 147992 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 147992 423654
rect -6596 423334 147992 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 147992 423334
rect -6596 423076 147992 423098
rect 451992 423654 590520 423676
rect 451992 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect 451992 423334 590520 423418
rect 451992 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect 451992 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 147992 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 147992 420054
rect -4756 419734 147992 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 147992 419734
rect -4756 419476 147992 419498
rect 451992 420054 588680 420076
rect 451992 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect 451992 419734 588680 419818
rect 451992 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect 451992 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 147992 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 147992 416454
rect -2916 416134 147992 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 147992 416134
rect -2916 415876 147992 415898
rect 451992 416454 586840 416476
rect 451992 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect 451992 416134 586840 416218
rect 451992 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect 451992 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 147992 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 147992 409254
rect -8436 408934 147992 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 147992 408934
rect -8436 408676 147992 408698
rect 451992 409254 592360 409276
rect 451992 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect 451992 408934 592360 409018
rect 451992 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect 451992 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 147992 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 147992 405654
rect -6596 405334 147992 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 147992 405334
rect -6596 405076 147992 405098
rect 451992 405654 590520 405676
rect 451992 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect 451992 405334 590520 405418
rect 451992 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect 451992 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 147992 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 147992 402054
rect -4756 401734 147992 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 147992 401734
rect -4756 401476 147992 401498
rect 451992 402054 588680 402076
rect 451992 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect 451992 401734 588680 401818
rect 451992 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect 451992 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 147992 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 147992 398454
rect -2916 398134 147992 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 147992 398134
rect -2916 397876 147992 397898
rect 451992 398454 586840 398476
rect 451992 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect 451992 398134 586840 398218
rect 451992 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect 451992 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 147992 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 147992 391254
rect -8436 390934 147992 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 147992 390934
rect -8436 390676 147992 390698
rect 451992 391254 592360 391276
rect 451992 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect 451992 390934 592360 391018
rect 451992 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect 451992 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 147992 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 147992 387654
rect -6596 387334 147992 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 147992 387334
rect -6596 387076 147992 387098
rect 451992 387654 590520 387676
rect 451992 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect 451992 387334 590520 387418
rect 451992 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect 451992 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 147992 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 147992 384054
rect -4756 383734 147992 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 147992 383734
rect -4756 383476 147992 383498
rect 451992 384054 588680 384076
rect 451992 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect 451992 383734 588680 383818
rect 451992 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect 451992 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 147992 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 147992 380454
rect -2916 380134 147992 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 147992 380134
rect -2916 379876 147992 379898
rect 451992 380454 586840 380476
rect 451992 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect 451992 380134 586840 380218
rect 451992 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect 451992 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 147992 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 147992 373254
rect -8436 372934 147992 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 147992 372934
rect -8436 372676 147992 372698
rect 451992 373254 592360 373276
rect 451992 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect 451992 372934 592360 373018
rect 451992 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect 451992 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 147992 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 147992 369654
rect -6596 369334 147992 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 147992 369334
rect -6596 369076 147992 369098
rect 451992 369654 590520 369676
rect 451992 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect 451992 369334 590520 369418
rect 451992 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect 451992 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 147992 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 147992 366054
rect -4756 365734 147992 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 147992 365734
rect -4756 365476 147992 365498
rect 451992 366054 588680 366076
rect 451992 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect 451992 365734 588680 365818
rect 451992 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect 451992 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 147992 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 147992 362454
rect -2916 362134 147992 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 147992 362134
rect -2916 361876 147992 361898
rect 451992 362454 586840 362476
rect 451992 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect 451992 362134 586840 362218
rect 451992 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect 451992 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 147992 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 147992 355254
rect -8436 354934 147992 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 147992 354934
rect -8436 354676 147992 354698
rect 451992 355254 592360 355276
rect 451992 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect 451992 354934 592360 355018
rect 451992 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect 451992 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 147992 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 147992 351654
rect -6596 351334 147992 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 147992 351334
rect -6596 351076 147992 351098
rect 451992 351654 590520 351676
rect 451992 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect 451992 351334 590520 351418
rect 451992 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect 451992 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 147992 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 147992 348054
rect -4756 347734 147992 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 147992 347734
rect -4756 347476 147992 347498
rect 451992 348054 588680 348076
rect 451992 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect 451992 347734 588680 347818
rect 451992 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect 451992 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 147992 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 147992 344454
rect -2916 344134 147992 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 147992 344134
rect -2916 343876 147992 343898
rect 451992 344454 586840 344476
rect 451992 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect 451992 344134 586840 344218
rect 451992 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect 451992 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 147992 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 147992 337254
rect -8436 336934 147992 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 147992 336934
rect -8436 336676 147992 336698
rect 451992 337254 592360 337276
rect 451992 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect 451992 336934 592360 337018
rect 451992 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect 451992 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 147992 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 147992 333654
rect -6596 333334 147992 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 147992 333334
rect -6596 333076 147992 333098
rect 451992 333654 590520 333676
rect 451992 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect 451992 333334 590520 333418
rect 451992 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect 451992 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 147992 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 147992 330054
rect -4756 329734 147992 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 147992 329734
rect -4756 329476 147992 329498
rect 451992 330054 588680 330076
rect 451992 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect 451992 329734 588680 329818
rect 451992 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect 451992 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 147992 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 147992 326454
rect -2916 326134 147992 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 147992 326134
rect -2916 325876 147992 325898
rect 451992 326454 586840 326476
rect 451992 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect 451992 326134 586840 326218
rect 451992 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect 451992 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 147992 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 147992 319254
rect -8436 318934 147992 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 147992 318934
rect -8436 318676 147992 318698
rect 451992 319254 592360 319276
rect 451992 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect 451992 318934 592360 319018
rect 451992 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect 451992 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 147992 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 147992 315654
rect -6596 315334 147992 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 147992 315334
rect -6596 315076 147992 315098
rect 451992 315654 590520 315676
rect 451992 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect 451992 315334 590520 315418
rect 451992 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect 451992 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 147992 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 147992 312054
rect -4756 311734 147992 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 147992 311734
rect -4756 311476 147992 311498
rect 451992 312054 588680 312076
rect 451992 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect 451992 311734 588680 311818
rect 451992 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect 451992 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 147992 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 147992 308454
rect -2916 308134 147992 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 147992 308134
rect -2916 307876 147992 307898
rect 451992 308454 586840 308476
rect 451992 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect 451992 308134 586840 308218
rect 451992 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect 451992 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 147992 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 147992 301254
rect -8436 300934 147992 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 147992 300934
rect -8436 300676 147992 300698
rect 451992 301254 592360 301276
rect 451992 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect 451992 300934 592360 301018
rect 451992 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect 451992 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 147992 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 147992 297654
rect -6596 297334 147992 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 147992 297334
rect -6596 297076 147992 297098
rect 451992 297654 590520 297676
rect 451992 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect 451992 297334 590520 297418
rect 451992 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect 451992 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 147992 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 147992 294054
rect -4756 293734 147992 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 147992 293734
rect -4756 293476 147992 293498
rect 451992 294054 588680 294076
rect 451992 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect 451992 293734 588680 293818
rect 451992 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect 451992 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 147992 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 147992 290454
rect -2916 290134 147992 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 147992 290134
rect -2916 289876 147992 289898
rect 451992 290454 586840 290476
rect 451992 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect 451992 290134 586840 290218
rect 451992 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect 451992 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 147992 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 147992 283254
rect -8436 282934 147992 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 147992 282934
rect -8436 282676 147992 282698
rect 451992 283254 592360 283276
rect 451992 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect 451992 282934 592360 283018
rect 451992 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect 451992 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 147992 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 147992 279654
rect -6596 279334 147992 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 147992 279334
rect -6596 279076 147992 279098
rect 451992 279654 590520 279676
rect 451992 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect 451992 279334 590520 279418
rect 451992 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect 451992 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 147992 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 147992 276054
rect -4756 275734 147992 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 147992 275734
rect -4756 275476 147992 275498
rect 451992 276054 588680 276076
rect 451992 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect 451992 275734 588680 275818
rect 451992 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect 451992 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 147992 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 147992 272454
rect -2916 272134 147992 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 147992 272134
rect -2916 271876 147992 271898
rect 451992 272454 586840 272476
rect 451992 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect 451992 272134 586840 272218
rect 451992 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect 451992 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 147992 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 147992 265254
rect -8436 264934 147992 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 147992 264934
rect -8436 264676 147992 264698
rect 451992 265254 592360 265276
rect 451992 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect 451992 264934 592360 265018
rect 451992 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect 451992 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 147992 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 147992 261654
rect -6596 261334 147992 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 147992 261334
rect -6596 261076 147992 261098
rect 451992 261654 590520 261676
rect 451992 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect 451992 261334 590520 261418
rect 451992 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect 451992 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 147992 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 147992 258054
rect -4756 257734 147992 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 147992 257734
rect -4756 257476 147992 257498
rect 451992 258054 588680 258076
rect 451992 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect 451992 257734 588680 257818
rect 451992 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect 451992 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 147992 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 147992 254454
rect -2916 254134 147992 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 147992 254134
rect -2916 253876 147992 253898
rect 451992 254454 586840 254476
rect 451992 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect 451992 254134 586840 254218
rect 451992 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect 451992 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 147992 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 147992 247254
rect -8436 246934 147992 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 147992 246934
rect -8436 246676 147992 246698
rect 451992 247254 592360 247276
rect 451992 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect 451992 246934 592360 247018
rect 451992 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect 451992 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 147992 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 147992 243654
rect -6596 243334 147992 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 147992 243334
rect -6596 243076 147992 243098
rect 451992 243654 590520 243676
rect 451992 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect 451992 243334 590520 243418
rect 451992 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect 451992 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1608069679
transform 1 0 149992 0 1 245136
box -1200 -1200 301200 301200
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
