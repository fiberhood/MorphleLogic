VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dummy_slave
  CLASS BLOCK ;
  FOREIGN dummy_slave ;
  ORIGIN 0.000 0.000 ;
  SIZE 107.040 BY 106.320 ;
  PIN wb_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END wb_ack_o
  PIN wb_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.000 0.000 6.280 4.000 ;
    END
  END wb_adr_i[0]
  PIN wb_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.500 0.000 40.780 4.000 ;
    END
  END wb_adr_i[10]
  PIN wb_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.720 0.000 44.000 4.000 ;
    END
  END wb_adr_i[11]
  PIN wb_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.480 0.000 46.760 4.000 ;
    END
  END wb_adr_i[12]
  PIN wb_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.700 0.000 49.980 4.000 ;
    END
  END wb_adr_i[13]
  PIN wb_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.920 0.000 53.200 4.000 ;
    END
  END wb_adr_i[14]
  PIN wb_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.680 0.000 55.960 4.000 ;
    END
  END wb_adr_i[15]
  PIN wb_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.900 0.000 59.180 4.000 ;
    END
  END wb_adr_i[16]
  PIN wb_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.120 0.000 62.400 4.000 ;
    END
  END wb_adr_i[17]
  PIN wb_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.880 0.000 65.160 4.000 ;
    END
  END wb_adr_i[18]
  PIN wb_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.100 0.000 68.380 4.000 ;
    END
  END wb_adr_i[19]
  PIN wb_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.140 0.000 10.420 4.000 ;
    END
  END wb_adr_i[1]
  PIN wb_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.320 0.000 71.600 4.000 ;
    END
  END wb_adr_i[20]
  PIN wb_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.080 0.000 74.360 4.000 ;
    END
  END wb_adr_i[21]
  PIN wb_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.300 0.000 77.580 4.000 ;
    END
  END wb_adr_i[22]
  PIN wb_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.520 0.000 80.800 4.000 ;
    END
  END wb_adr_i[23]
  PIN wb_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.280 0.000 83.560 4.000 ;
    END
  END wb_adr_i[24]
  PIN wb_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.500 0.000 86.780 4.000 ;
    END
  END wb_adr_i[25]
  PIN wb_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.720 0.000 90.000 4.000 ;
    END
  END wb_adr_i[26]
  PIN wb_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.480 0.000 92.760 4.000 ;
    END
  END wb_adr_i[27]
  PIN wb_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.700 0.000 95.980 4.000 ;
    END
  END wb_adr_i[28]
  PIN wb_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.920 0.000 99.200 4.000 ;
    END
  END wb_adr_i[29]
  PIN wb_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.280 0.000 14.560 4.000 ;
    END
  END wb_adr_i[2]
  PIN wb_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.680 0.000 101.960 4.000 ;
    END
  END wb_adr_i[30]
  PIN wb_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.900 0.000 105.180 4.000 ;
    END
  END wb_adr_i[31]
  PIN wb_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.960 0.000 18.240 4.000 ;
    END
  END wb_adr_i[3]
  PIN wb_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.100 0.000 22.380 4.000 ;
    END
  END wb_adr_i[4]
  PIN wb_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.320 0.000 25.600 4.000 ;
    END
  END wb_adr_i[5]
  PIN wb_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.540 0.000 28.820 4.000 ;
    END
  END wb_adr_i[6]
  PIN wb_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.300 0.000 31.580 4.000 ;
    END
  END wb_adr_i[7]
  PIN wb_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.520 0.000 34.800 4.000 ;
    END
  END wb_adr_i[8]
  PIN wb_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.740 0.000 38.020 4.000 ;
    END
  END wb_adr_i[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.940 0.000 1.220 4.000 ;
    END
  END wb_clk_i
  PIN wb_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.860 0.000 2.140 4.000 ;
    END
  END wb_cyc_i
  PIN wb_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.920 0.000 7.200 4.000 ;
    END
  END wb_dat_i[0]
  PIN wb_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.420 0.000 41.700 4.000 ;
    END
  END wb_dat_i[10]
  PIN wb_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.640 0.000 44.920 4.000 ;
    END
  END wb_dat_i[11]
  PIN wb_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.860 0.000 48.140 4.000 ;
    END
  END wb_dat_i[12]
  PIN wb_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.620 0.000 50.900 4.000 ;
    END
  END wb_dat_i[13]
  PIN wb_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.840 0.000 54.120 4.000 ;
    END
  END wb_dat_i[14]
  PIN wb_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.060 0.000 57.340 4.000 ;
    END
  END wb_dat_i[15]
  PIN wb_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.820 0.000 60.100 4.000 ;
    END
  END wb_dat_i[16]
  PIN wb_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.040 0.000 63.320 4.000 ;
    END
  END wb_dat_i[17]
  PIN wb_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.260 0.000 66.540 4.000 ;
    END
  END wb_dat_i[18]
  PIN wb_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.020 0.000 69.300 4.000 ;
    END
  END wb_dat_i[19]
  PIN wb_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.060 0.000 11.340 4.000 ;
    END
  END wb_dat_i[1]
  PIN wb_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.240 0.000 72.520 4.000 ;
    END
  END wb_dat_i[20]
  PIN wb_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.460 0.000 75.740 4.000 ;
    END
  END wb_dat_i[21]
  PIN wb_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.220 0.000 78.500 4.000 ;
    END
  END wb_dat_i[22]
  PIN wb_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.440 0.000 81.720 4.000 ;
    END
  END wb_dat_i[23]
  PIN wb_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.660 0.000 84.940 4.000 ;
    END
  END wb_dat_i[24]
  PIN wb_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.420 0.000 87.700 4.000 ;
    END
  END wb_dat_i[25]
  PIN wb_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.640 0.000 90.920 4.000 ;
    END
  END wb_dat_i[26]
  PIN wb_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.400 0.000 93.680 4.000 ;
    END
  END wb_dat_i[27]
  PIN wb_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.620 0.000 96.900 4.000 ;
    END
  END wb_dat_i[28]
  PIN wb_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.840 0.000 100.120 4.000 ;
    END
  END wb_dat_i[29]
  PIN wb_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.200 0.000 15.480 4.000 ;
    END
  END wb_dat_i[2]
  PIN wb_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 102.600 0.000 102.880 4.000 ;
    END
  END wb_dat_i[30]
  PIN wb_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.820 0.000 106.100 4.000 ;
    END
  END wb_dat_i[31]
  PIN wb_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.340 0.000 19.620 4.000 ;
    END
  END wb_dat_i[3]
  PIN wb_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.020 0.000 23.300 4.000 ;
    END
  END wb_dat_i[4]
  PIN wb_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.240 0.000 26.520 4.000 ;
    END
  END wb_dat_i[5]
  PIN wb_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.460 0.000 29.740 4.000 ;
    END
  END wb_dat_i[6]
  PIN wb_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.220 0.000 32.500 4.000 ;
    END
  END wb_dat_i[7]
  PIN wb_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.440 0.000 35.720 4.000 ;
    END
  END wb_dat_i[8]
  PIN wb_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.660 0.000 38.940 4.000 ;
    END
  END wb_dat_i[9]
  PIN wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.840 0.000 8.120 4.000 ;
    END
  END wb_dat_o[0]
  PIN wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 42.800 0.000 43.080 4.000 ;
    END
  END wb_dat_o[10]
  PIN wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.560 0.000 45.840 4.000 ;
    END
  END wb_dat_o[11]
  PIN wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.780 0.000 49.060 4.000 ;
    END
  END wb_dat_o[12]
  PIN wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 52.000 0.000 52.280 4.000 ;
    END
  END wb_dat_o[13]
  PIN wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.760 0.000 55.040 4.000 ;
    END
  END wb_dat_o[14]
  PIN wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.980 0.000 58.260 4.000 ;
    END
  END wb_dat_o[15]
  PIN wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.200 0.000 61.480 4.000 ;
    END
  END wb_dat_o[16]
  PIN wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.960 0.000 64.240 4.000 ;
    END
  END wb_dat_o[17]
  PIN wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.180 0.000 67.460 4.000 ;
    END
  END wb_dat_o[18]
  PIN wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.940 0.000 70.220 4.000 ;
    END
  END wb_dat_o[19]
  PIN wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.980 0.000 12.260 4.000 ;
    END
  END wb_dat_o[1]
  PIN wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.160 0.000 73.440 4.000 ;
    END
  END wb_dat_o[20]
  PIN wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.380 0.000 76.660 4.000 ;
    END
  END wb_dat_o[21]
  PIN wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.140 0.000 79.420 4.000 ;
    END
  END wb_dat_o[22]
  PIN wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.360 0.000 82.640 4.000 ;
    END
  END wb_dat_o[23]
  PIN wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.580 0.000 85.860 4.000 ;
    END
  END wb_dat_o[24]
  PIN wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.340 0.000 88.620 4.000 ;
    END
  END wb_dat_o[25]
  PIN wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.560 0.000 91.840 4.000 ;
    END
  END wb_dat_o[26]
  PIN wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.780 0.000 95.060 4.000 ;
    END
  END wb_dat_o[27]
  PIN wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.540 0.000 97.820 4.000 ;
    END
  END wb_dat_o[28]
  PIN wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.760 0.000 101.040 4.000 ;
    END
  END wb_dat_o[29]
  PIN wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.120 0.000 16.400 4.000 ;
    END
  END wb_dat_o[2]
  PIN wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.980 0.000 104.260 4.000 ;
    END
  END wb_dat_o[30]
  PIN wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.740 0.000 107.020 4.000 ;
    END
  END wb_dat_o[31]
  PIN wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.260 0.000 20.540 4.000 ;
    END
  END wb_dat_o[3]
  PIN wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.400 0.000 24.680 4.000 ;
    END
  END wb_dat_o[4]
  PIN wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.160 0.000 27.440 4.000 ;
    END
  END wb_dat_o[5]
  PIN wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.380 0.000 30.660 4.000 ;
    END
  END wb_dat_o[6]
  PIN wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.600 0.000 33.880 4.000 ;
    END
  END wb_dat_o[7]
  PIN wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.360 0.000 36.640 4.000 ;
    END
  END wb_dat_o[8]
  PIN wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.580 0.000 39.860 4.000 ;
    END
  END wb_dat_o[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.780 0.000 3.060 4.000 ;
    END
  END wb_rst_i
  PIN wb_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.760 0.000 9.040 4.000 ;
    END
  END wb_sel_i[0]
  PIN wb_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.900 0.000 13.180 4.000 ;
    END
  END wb_sel_i[1]
  PIN wb_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.040 0.000 17.320 4.000 ;
    END
  END wb_sel_i[2]
  PIN wb_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.180 0.000 21.460 4.000 ;
    END
  END wb_sel_i[3]
  PIN wb_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.700 0.000 3.980 4.000 ;
    END
  END wb_stb_i
  PIN wb_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.080 0.000 5.360 4.000 ;
    END
  END wb_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.290 10.640 21.890 106.320 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 36.390 10.640 37.990 106.320 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.990 10.795 101.590 106.165 ;
      LAYER met1 ;
        RECT 0.000 6.840 107.040 106.320 ;
      LAYER met2 ;
        RECT 0.030 4.280 107.010 106.320 ;
        RECT 0.580 4.000 0.660 4.280 ;
        RECT 1.500 4.000 1.580 4.280 ;
        RECT 2.420 4.000 2.500 4.280 ;
        RECT 3.340 4.000 3.420 4.280 ;
        RECT 4.260 4.000 4.800 4.280 ;
        RECT 5.640 4.000 5.720 4.280 ;
        RECT 6.560 4.000 6.640 4.280 ;
        RECT 7.480 4.000 7.560 4.280 ;
        RECT 8.400 4.000 8.480 4.280 ;
        RECT 9.320 4.000 9.860 4.280 ;
        RECT 10.700 4.000 10.780 4.280 ;
        RECT 11.620 4.000 11.700 4.280 ;
        RECT 12.540 4.000 12.620 4.280 ;
        RECT 13.460 4.000 14.000 4.280 ;
        RECT 14.840 4.000 14.920 4.280 ;
        RECT 15.760 4.000 15.840 4.280 ;
        RECT 16.680 4.000 16.760 4.280 ;
        RECT 17.600 4.000 17.680 4.280 ;
        RECT 18.520 4.000 19.060 4.280 ;
        RECT 19.900 4.000 19.980 4.280 ;
        RECT 20.820 4.000 20.900 4.280 ;
        RECT 21.740 4.000 21.820 4.280 ;
        RECT 22.660 4.000 22.740 4.280 ;
        RECT 23.580 4.000 24.120 4.280 ;
        RECT 24.960 4.000 25.040 4.280 ;
        RECT 25.880 4.000 25.960 4.280 ;
        RECT 26.800 4.000 26.880 4.280 ;
        RECT 27.720 4.000 28.260 4.280 ;
        RECT 29.100 4.000 29.180 4.280 ;
        RECT 30.020 4.000 30.100 4.280 ;
        RECT 30.940 4.000 31.020 4.280 ;
        RECT 31.860 4.000 31.940 4.280 ;
        RECT 32.780 4.000 33.320 4.280 ;
        RECT 34.160 4.000 34.240 4.280 ;
        RECT 35.080 4.000 35.160 4.280 ;
        RECT 36.000 4.000 36.080 4.280 ;
        RECT 36.920 4.000 37.460 4.280 ;
        RECT 38.300 4.000 38.380 4.280 ;
        RECT 39.220 4.000 39.300 4.280 ;
        RECT 40.140 4.000 40.220 4.280 ;
        RECT 41.060 4.000 41.140 4.280 ;
        RECT 41.980 4.000 42.520 4.280 ;
        RECT 43.360 4.000 43.440 4.280 ;
        RECT 44.280 4.000 44.360 4.280 ;
        RECT 45.200 4.000 45.280 4.280 ;
        RECT 46.120 4.000 46.200 4.280 ;
        RECT 47.040 4.000 47.580 4.280 ;
        RECT 48.420 4.000 48.500 4.280 ;
        RECT 49.340 4.000 49.420 4.280 ;
        RECT 50.260 4.000 50.340 4.280 ;
        RECT 51.180 4.000 51.720 4.280 ;
        RECT 52.560 4.000 52.640 4.280 ;
        RECT 53.480 4.000 53.560 4.280 ;
        RECT 54.400 4.000 54.480 4.280 ;
        RECT 55.320 4.000 55.400 4.280 ;
        RECT 56.240 4.000 56.780 4.280 ;
        RECT 57.620 4.000 57.700 4.280 ;
        RECT 58.540 4.000 58.620 4.280 ;
        RECT 59.460 4.000 59.540 4.280 ;
        RECT 60.380 4.000 60.920 4.280 ;
        RECT 61.760 4.000 61.840 4.280 ;
        RECT 62.680 4.000 62.760 4.280 ;
        RECT 63.600 4.000 63.680 4.280 ;
        RECT 64.520 4.000 64.600 4.280 ;
        RECT 65.440 4.000 65.980 4.280 ;
        RECT 66.820 4.000 66.900 4.280 ;
        RECT 67.740 4.000 67.820 4.280 ;
        RECT 68.660 4.000 68.740 4.280 ;
        RECT 69.580 4.000 69.660 4.280 ;
        RECT 70.500 4.000 71.040 4.280 ;
        RECT 71.880 4.000 71.960 4.280 ;
        RECT 72.800 4.000 72.880 4.280 ;
        RECT 73.720 4.000 73.800 4.280 ;
        RECT 74.640 4.000 75.180 4.280 ;
        RECT 76.020 4.000 76.100 4.280 ;
        RECT 76.940 4.000 77.020 4.280 ;
        RECT 77.860 4.000 77.940 4.280 ;
        RECT 78.780 4.000 78.860 4.280 ;
        RECT 79.700 4.000 80.240 4.280 ;
        RECT 81.080 4.000 81.160 4.280 ;
        RECT 82.000 4.000 82.080 4.280 ;
        RECT 82.920 4.000 83.000 4.280 ;
        RECT 83.840 4.000 84.380 4.280 ;
        RECT 85.220 4.000 85.300 4.280 ;
        RECT 86.140 4.000 86.220 4.280 ;
        RECT 87.060 4.000 87.140 4.280 ;
        RECT 87.980 4.000 88.060 4.280 ;
        RECT 88.900 4.000 89.440 4.280 ;
        RECT 90.280 4.000 90.360 4.280 ;
        RECT 91.200 4.000 91.280 4.280 ;
        RECT 92.120 4.000 92.200 4.280 ;
        RECT 93.040 4.000 93.120 4.280 ;
        RECT 93.960 4.000 94.500 4.280 ;
        RECT 95.340 4.000 95.420 4.280 ;
        RECT 96.260 4.000 96.340 4.280 ;
        RECT 97.180 4.000 97.260 4.280 ;
        RECT 98.100 4.000 98.640 4.280 ;
        RECT 99.480 4.000 99.560 4.280 ;
        RECT 100.400 4.000 100.480 4.280 ;
        RECT 101.320 4.000 101.400 4.280 ;
        RECT 102.240 4.000 102.320 4.280 ;
        RECT 103.160 4.000 103.700 4.280 ;
        RECT 104.540 4.000 104.620 4.280 ;
        RECT 105.460 4.000 105.540 4.280 ;
        RECT 106.380 4.000 106.460 4.280 ;
      LAYER met3 ;
        RECT 5.055 10.715 96.925 106.245 ;
      LAYER met4 ;
        RECT 14.485 10.640 19.890 106.320 ;
        RECT 22.290 10.640 35.990 106.320 ;
        RECT 38.390 10.640 95.775 106.320 ;
  END
END dummy_slave
END LIBRARY

