* NGSPICE file created from user_proj_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for ycell abstract view
.subckt ycell cbitin cbitout confclk confclko dempty din[0] din[1] dout[0] dout[1]
+ hempty hempty2 lempty lin[0] lin[1] lout[0] lout[1] rempty reset reseto rin[0] rin[1]
+ rout[0] rout[1] uempty uin[0] uin[1] uout[0] uout[1] vempty vempty2 VPWR VGND
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i VPWR VGND
XFILLER_42_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_223_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_501_ VGND VGND VPWR VPWR _501_/HI _501_/LO sky130_fd_sc_hd__conb_1
XFILLER_499_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_432_ VGND VGND VPWR VPWR _432_/HI _432_/LO sky130_fd_sc_hd__conb_1
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_363_ _363_/A VGND VGND VPWR VPWR _363_/Y sky130_fd_sc_hd__inv_2
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_294_ _807_/Q VGND VGND VPWR VPWR _294_/Y sky130_fd_sc_hd__inv_2
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[2\].yc blk.column\[8\].row\[2\].yc/cbitin blk.column\[8\].row\[3\].yc/cbitin
+ blk.column\[8\].row\[2\].yc/confclk blk.column\[8\].row\[3\].yc/confclk blk.column\[8\].row\[2\].yc/dempty
+ blk.column\[8\].row\[2\].yc/din[0] blk.column\[8\].row\[2\].yc/din[1] blk.column\[8\].row\[3\].yc/uin[0]
+ blk.column\[8\].row\[3\].yc/uin[1] blk.column\[8\].row\[2\].yc/hempty blk.column\[7\].row\[2\].yc/lempty
+ blk.column\[8\].row\[2\].yc/lempty blk.column\[8\].row\[2\].yc/lin[0] blk.column\[8\].row\[2\].yc/lin[1]
+ blk.column\[9\].row\[2\].yc/rin[0] blk.column\[9\].row\[2\].yc/rin[1] blk.column\[7\].row\[2\].yc/hempty
+ blk.column\[8\].row\[2\].yc/reset blk.column\[8\].row\[3\].yc/reset blk.column\[8\].row\[2\].yc/rin[0]
+ blk.column\[8\].row\[2\].yc/rin[1] blk.column\[7\].row\[2\].yc/lin[0] blk.column\[7\].row\[2\].yc/lin[1]
+ blk.column\[8\].row\[2\].yc/uempty blk.column\[8\].row\[2\].yc/uin[0] blk.column\[8\].row\[2\].yc/uin[1]
+ blk.column\[8\].row\[1\].yc/din[0] blk.column\[8\].row\[1\].yc/din[1] blk.column\[8\].row\[1\].yc/dempty
+ blk.column\[8\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_515_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_457_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_482_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_523_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_539_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_338_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_492_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[10\].yc blk.column\[2\].row\[9\].yc/cbitout blk.column\[2\].row\[11\].yc/cbitin
+ blk.column\[2\].row\[9\].yc/confclko blk.column\[2\].row\[11\].yc/confclk blk.column\[2\].row\[10\].yc/dempty
+ blk.column\[2\].row\[10\].yc/din[0] blk.column\[2\].row\[10\].yc/din[1] blk.column\[2\].row\[11\].yc/uin[0]
+ blk.column\[2\].row\[11\].yc/uin[1] blk.column\[2\].row\[10\].yc/hempty blk.column\[1\].row\[10\].yc/lempty
+ blk.column\[2\].row\[10\].yc/lempty blk.column\[2\].row\[10\].yc/lin[0] blk.column\[2\].row\[10\].yc/lin[1]
+ blk.column\[3\].row\[10\].yc/rin[0] blk.column\[3\].row\[10\].yc/rin[1] blk.column\[1\].row\[10\].yc/hempty
+ blk.column\[2\].row\[9\].yc/reseto blk.column\[2\].row\[11\].yc/reset blk.column\[2\].row\[10\].yc/rin[0]
+ blk.column\[2\].row\[10\].yc/rin[1] blk.column\[1\].row\[10\].yc/lin[0] blk.column\[1\].row\[10\].yc/lin[1]
+ blk.column\[2\].row\[9\].yc/vempty2 blk.column\[2\].row\[9\].yc/dout[0] blk.column\[2\].row\[9\].yc/dout[1]
+ blk.column\[2\].row\[9\].yc/din[0] blk.column\[2\].row\[9\].yc/din[1] blk.column\[2\].row\[9\].yc/dempty
+ blk.column\[2\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_511_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_448_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_515_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_528_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_531_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_384_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_492_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_492_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_352_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_486_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_273_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_415_ _412_/X wbs_dat_o[8] _335_/A _410_/X VGND VGND VPWR VPWR _752_/D sky130_fd_sc_hd__o22a_4
XPHY_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_501_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_346_ _344_/Y _340_/X wbs_dat_i[21] _345_/X VGND VGND VPWR VPWR _789_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_538_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_358_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_532_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_229_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_451_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_369_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_384_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[9\].yc blk.column\[13\].row\[9\].yc/cbitin blk.column\[13\].row\[9\].yc/cbitout
+ blk.column\[13\].row\[9\].yc/confclk blk.column\[13\].row\[9\].yc/confclko blk.column\[13\].row\[9\].yc/dempty
+ blk.column\[13\].row\[9\].yc/din[0] blk.column\[13\].row\[9\].yc/din[1] blk.column\[13\].row\[9\].yc/dout[0]
+ blk.column\[13\].row\[9\].yc/dout[1] blk.column\[13\].row\[9\].yc/hempty blk.column\[12\].row\[9\].yc/lempty
+ blk.column\[13\].row\[9\].yc/lempty blk.column\[13\].row\[9\].yc/lin[0] blk.column\[13\].row\[9\].yc/lin[1]
+ blk.column\[14\].row\[9\].yc/rin[0] blk.column\[14\].row\[9\].yc/rin[1] blk.column\[12\].row\[9\].yc/hempty
+ blk.column\[13\].row\[9\].yc/reset blk.column\[13\].row\[9\].yc/reseto blk.column\[13\].row\[9\].yc/rin[0]
+ blk.column\[13\].row\[9\].yc/rin[1] blk.column\[12\].row\[9\].yc/lin[0] blk.column\[12\].row\[9\].yc/lin[1]
+ blk.column\[13\].row\[9\].yc/uempty blk.column\[13\].row\[9\].yc/uin[0] blk.column\[13\].row\[9\].yc/uin[1]
+ blk.column\[13\].row\[8\].yc/din[0] blk.column\[13\].row\[8\].yc/din[1] blk.column\[13\].row\[8\].yc/dempty
+ blk.column\[13\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_499_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_464_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_284_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_348_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_3019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_540_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_329_ _328_/Y _324_/X wbs_dat_i[11] _324_/X VGND VGND VPWR VPWR _795_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_524_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_493_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_390_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_514_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_680_ VGND VGND VPWR VPWR _680_/HI la_data_out[64] sky130_fd_sc_hd__conb_1
XPHY_6857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_324_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_498_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[4\].yc blk.column\[9\].row\[4\].yc/cbitin blk.column\[9\].row\[5\].yc/cbitin
+ blk.column\[9\].row\[4\].yc/confclk blk.column\[9\].row\[5\].yc/confclk blk.column\[9\].row\[4\].yc/dempty
+ blk.column\[9\].row\[4\].yc/din[0] blk.column\[9\].row\[4\].yc/din[1] blk.column\[9\].row\[5\].yc/uin[0]
+ blk.column\[9\].row\[5\].yc/uin[1] blk.column\[9\].row\[4\].yc/hempty blk.column\[8\].row\[4\].yc/lempty
+ blk.column\[9\].row\[4\].yc/lempty blk.column\[9\].row\[4\].yc/lin[0] blk.column\[9\].row\[4\].yc/lin[1]
+ blk.column\[9\].row\[4\].yc/lout[0] blk.column\[9\].row\[4\].yc/lout[1] blk.column\[8\].row\[4\].yc/hempty
+ blk.column\[9\].row\[4\].yc/reset blk.column\[9\].row\[5\].yc/reset blk.column\[9\].row\[4\].yc/rin[0]
+ blk.column\[9\].row\[4\].yc/rin[1] blk.column\[8\].row\[4\].yc/lin[0] blk.column\[8\].row\[4\].yc/lin[1]
+ blk.column\[9\].row\[4\].yc/uempty blk.column\[9\].row\[4\].yc/uin[0] blk.column\[9\].row\[4\].yc/uin[1]
+ blk.column\[9\].row\[3\].yc/din[0] blk.column\[9\].row\[3\].yc/din[1] blk.column\[9\].row\[3\].yc/dempty
+ blk.column\[9\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_203_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_455_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_517_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_537_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_474_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[13\].yc blk.column\[6\].row\[13\].yc/cbitin blk.column\[6\].row\[14\].yc/cbitin
+ blk.column\[6\].row\[13\].yc/confclk blk.column\[6\].row\[14\].yc/confclk blk.column\[6\].row\[13\].yc/dempty
+ blk.column\[6\].row\[13\].yc/din[0] blk.column\[6\].row\[13\].yc/din[1] blk.column\[6\].row\[14\].yc/uin[0]
+ blk.column\[6\].row\[14\].yc/uin[1] blk.column\[6\].row\[13\].yc/hempty blk.column\[5\].row\[13\].yc/lempty
+ blk.column\[6\].row\[13\].yc/lempty blk.column\[6\].row\[13\].yc/lin[0] blk.column\[6\].row\[13\].yc/lin[1]
+ blk.column\[7\].row\[13\].yc/rin[0] blk.column\[7\].row\[13\].yc/rin[1] blk.column\[5\].row\[13\].yc/hempty
+ blk.column\[6\].row\[13\].yc/reset blk.column\[6\].row\[14\].yc/reset blk.column\[6\].row\[13\].yc/rin[0]
+ blk.column\[6\].row\[13\].yc/rin[1] blk.column\[5\].row\[13\].yc/lin[0] blk.column\[5\].row\[13\].yc/lin[1]
+ blk.column\[6\].row\[13\].yc/uempty blk.column\[6\].row\[13\].yc/uin[0] blk.column\[6\].row\[13\].yc/uin[1]
+ blk.column\[6\].row\[12\].yc/din[0] blk.column\[6\].row\[12\].yc/din[1] blk.column\[6\].row\[12\].yc/dempty
+ blk.column\[6\].row\[14\].yc/uempty VPWR VGND ycell
XPHY_9494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_282_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_495_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_468_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_304_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_531_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_540_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_801_ wb_clk_i _313_/X VGND VGND VPWR VPWR _312_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_40_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_732_ VGND VGND VPWR VPWR _732_/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XPHY_7377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_663_ VGND VGND VPWR VPWR _663_/HI io_out[37] sky130_fd_sc_hd__conb_1
XFILLER_483_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_594_ VGND VGND VPWR VPWR _594_/HI io_oeb[6] sky130_fd_sc_hd__conb_1
XPHY_5986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_318_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_430_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_522_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_380_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[13\].row\[15\].yc blk.column\[13\].row\[15\].yc/cbitin la_data_out[45]
+ blk.column\[13\].row\[15\].yc/confclk blk.column\[13\].row\[15\].yc/confclko _448_/HI
+ _521_/LO _522_/LO blk.column\[13\].row\[15\].yc/dout[0] blk.column\[13\].row\[15\].yc/dout[1]
+ blk.column\[13\].row\[15\].yc/hempty blk.column\[12\].row\[15\].yc/lempty blk.column\[13\].row\[15\].yc/lempty
+ blk.column\[13\].row\[15\].yc/lin[0] blk.column\[13\].row\[15\].yc/lin[1] blk.column\[14\].row\[15\].yc/rin[0]
+ blk.column\[14\].row\[15\].yc/rin[1] blk.column\[12\].row\[15\].yc/hempty blk.column\[13\].row\[15\].yc/reset
+ blk.column\[13\].row\[15\].yc/reseto blk.column\[13\].row\[15\].yc/rin[0] blk.column\[13\].row\[15\].yc/rin[1]
+ blk.column\[12\].row\[15\].yc/lin[0] blk.column\[12\].row\[15\].yc/lin[1] blk.column\[13\].row\[15\].yc/uempty
+ blk.column\[13\].row\[15\].yc/uin[0] blk.column\[13\].row\[15\].yc/uin[1] blk.column\[13\].row\[14\].yc/din[0]
+ blk.column\[13\].row\[14\].yc/din[1] blk.column\[13\].row\[14\].yc/dempty blk.column\[13\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_360_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_260_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_213_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_401_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_313_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_715_ VGND VGND VPWR VPWR _715_/HI la_data_out[99] sky130_fd_sc_hd__conb_1
XPHY_6473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_389_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_646_ VGND VGND VPWR VPWR _646_/HI io_out[20] sky130_fd_sc_hd__conb_1
XFILLER_504_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_320_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_577_ VGND VGND VPWR VPWR _577_/HI _577_/LO sky130_fd_sc_hd__conb_1
XFILLER_400_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_272_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_487_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_411_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_356_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_533_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_510_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_500_ VGND VGND VPWR VPWR _500_/HI _500_/LO sky130_fd_sc_hd__conb_1
XPHY_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_431_ VGND VGND VPWR VPWR _431_/HI _431_/LO sky130_fd_sc_hd__conb_1
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_362_ _358_/Y _361_/X wbs_dat_i[31] _361_/X VGND VGND VPWR VPWR _362_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_332_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_439_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_469_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_629_ VGND VGND VPWR VPWR _629_/HI io_out[3] sky130_fd_sc_hd__conb_1
XFILLER_500_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_359_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_338_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_255_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_530_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_303_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[5\].yc blk.column\[0\].row\[5\].yc/cbitin blk.column\[0\].row\[6\].yc/cbitin
+ blk.column\[0\].row\[5\].yc/confclk blk.column\[0\].row\[6\].yc/confclk blk.column\[0\].row\[5\].yc/dempty
+ blk.column\[0\].row\[5\].yc/din[0] blk.column\[0\].row\[5\].yc/din[1] blk.column\[0\].row\[6\].yc/uin[0]
+ blk.column\[0\].row\[6\].yc/uin[1] blk.column\[0\].row\[5\].yc/hempty blk.column\[0\].row\[5\].yc/hempty2
+ blk.column\[0\].row\[5\].yc/lempty blk.column\[0\].row\[5\].yc/lin[0] blk.column\[0\].row\[5\].yc/lin[1]
+ blk.column\[1\].row\[5\].yc/rin[0] blk.column\[1\].row\[5\].yc/rin[1] _440_/HI blk.column\[0\].row\[5\].yc/reset
+ blk.column\[0\].row\[6\].yc/reset _501_/LO _502_/LO blk.column\[0\].row\[5\].yc/rout[0]
+ blk.column\[0\].row\[5\].yc/rout[1] blk.column\[0\].row\[5\].yc/uempty blk.column\[0\].row\[5\].yc/uin[0]
+ blk.column\[0\].row\[5\].yc/uin[1] blk.column\[0\].row\[4\].yc/din[0] blk.column\[0\].row\[4\].yc/din[1]
+ blk.column\[0\].row\[4\].yc/dempty blk.column\[0\].row\[6\].yc/uempty VPWR VGND
+ ycell
XPHY_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_369_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_400_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_250_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_476_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_453_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_529_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_523_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_407_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_414_ _412_/X wbs_dat_o[9] _333_/A _410_/X VGND VGND VPWR VPWR _753_/D sky130_fd_sc_hd__o22a_4
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_345_ _339_/X VGND VGND VPWR VPWR _345_/X sky130_fd_sc_hd__buf_2
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_521_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_278_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_303_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[14\].yc blk.column\[1\].row\[14\].yc/cbitin blk.column\[1\].row\[15\].yc/cbitin
+ blk.column\[1\].row\[14\].yc/confclk blk.column\[1\].row\[15\].yc/confclk blk.column\[1\].row\[14\].yc/dempty
+ blk.column\[1\].row\[14\].yc/din[0] blk.column\[1\].row\[14\].yc/din[1] blk.column\[1\].row\[15\].yc/uin[0]
+ blk.column\[1\].row\[15\].yc/uin[1] blk.column\[1\].row\[14\].yc/hempty blk.column\[0\].row\[14\].yc/lempty
+ blk.column\[1\].row\[14\].yc/lempty blk.column\[1\].row\[14\].yc/lin[0] blk.column\[1\].row\[14\].yc/lin[1]
+ blk.column\[2\].row\[14\].yc/rin[0] blk.column\[2\].row\[14\].yc/rin[1] blk.column\[0\].row\[14\].yc/hempty
+ blk.column\[1\].row\[14\].yc/reset blk.column\[1\].row\[15\].yc/reset blk.column\[1\].row\[14\].yc/rin[0]
+ blk.column\[1\].row\[14\].yc/rin[1] blk.column\[0\].row\[14\].yc/lin[0] blk.column\[0\].row\[14\].yc/lin[1]
+ blk.column\[1\].row\[14\].yc/uempty blk.column\[1\].row\[14\].yc/uin[0] blk.column\[1\].row\[14\].yc/uin[1]
+ blk.column\[1\].row\[13\].yc/din[0] blk.column\[1\].row\[13\].yc/din[1] blk.column\[1\].row\[13\].yc/dempty
+ blk.column\[1\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_390_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_414_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[10\].yc blk.column\[15\].row\[9\].yc/cbitout blk.column\[15\].row\[11\].yc/cbitin
+ blk.column\[15\].row\[9\].yc/confclko blk.column\[15\].row\[11\].yc/confclk blk.column\[15\].row\[10\].yc/dempty
+ blk.column\[15\].row\[10\].yc/din[0] blk.column\[15\].row\[10\].yc/din[1] blk.column\[15\].row\[11\].yc/uin[0]
+ blk.column\[15\].row\[11\].yc/uin[1] blk.column\[15\].row\[10\].yc/hempty blk.column\[14\].row\[10\].yc/lempty
+ _451_/HI _529_/LO _530_/LO blk.column\[15\].row\[10\].yc/lout[0] blk.column\[15\].row\[10\].yc/lout[1]
+ blk.column\[14\].row\[10\].yc/hempty blk.column\[15\].row\[9\].yc/reseto blk.column\[15\].row\[11\].yc/reset
+ blk.column\[15\].row\[10\].yc/rin[0] blk.column\[15\].row\[10\].yc/rin[1] blk.column\[14\].row\[10\].yc/lin[0]
+ blk.column\[14\].row\[10\].yc/lin[1] blk.column\[15\].row\[9\].yc/vempty2 blk.column\[15\].row\[9\].yc/dout[0]
+ blk.column\[15\].row\[9\].yc/dout[1] blk.column\[15\].row\[9\].yc/din[0] blk.column\[15\].row\[9\].yc/din[1]
+ blk.column\[15\].row\[9\].yc/dempty blk.column\[15\].row\[11\].yc/uempty VPWR VGND
+ ycell
XFILLER_441_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_372_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_536_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_517_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_255_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_494_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_372_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_535_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_483_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_501_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_348_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_401_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_328_ _795_/Q VGND VGND VPWR VPWR _328_/Y sky130_fd_sc_hd__inv_2
XFILLER_501_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_252_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_541_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_257_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_268_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_344_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_363_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_404_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_355_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_529_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_423_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_488_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[6\].yc blk.column\[10\].row\[6\].yc/cbitin blk.column\[10\].row\[7\].yc/cbitin
+ blk.column\[10\].row\[6\].yc/confclk blk.column\[10\].row\[7\].yc/confclk blk.column\[10\].row\[6\].yc/dempty
+ blk.column\[10\].row\[6\].yc/din[0] blk.column\[10\].row\[6\].yc/din[1] blk.column\[10\].row\[7\].yc/uin[0]
+ blk.column\[10\].row\[7\].yc/uin[1] blk.column\[10\].row\[6\].yc/hempty blk.column\[9\].row\[6\].yc/lempty
+ blk.column\[10\].row\[6\].yc/lempty blk.column\[10\].row\[6\].yc/lin[0] blk.column\[10\].row\[6\].yc/lin[1]
+ blk.column\[11\].row\[6\].yc/rin[0] blk.column\[11\].row\[6\].yc/rin[1] blk.column\[9\].row\[6\].yc/hempty
+ blk.column\[10\].row\[6\].yc/reset blk.column\[10\].row\[7\].yc/reset blk.column\[9\].row\[6\].yc/lout[0]
+ blk.column\[9\].row\[6\].yc/lout[1] blk.column\[9\].row\[6\].yc/lin[0] blk.column\[9\].row\[6\].yc/lin[1]
+ blk.column\[10\].row\[6\].yc/uempty blk.column\[10\].row\[6\].yc/uin[0] blk.column\[10\].row\[6\].yc/uin[1]
+ blk.column\[10\].row\[5\].yc/din[0] blk.column\[10\].row\[5\].yc/din[1] blk.column\[10\].row\[5\].yc/dempty
+ blk.column\[10\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_363_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_484_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[7\].yc blk.column\[1\].row\[7\].yc/cbitin blk.column\[1\].row\[8\].yc/cbitin
+ blk.column\[1\].row\[7\].yc/confclk blk.column\[1\].row\[8\].yc/confclk blk.column\[1\].row\[7\].yc/dempty
+ blk.column\[1\].row\[7\].yc/din[0] blk.column\[1\].row\[7\].yc/din[1] blk.column\[1\].row\[8\].yc/uin[0]
+ blk.column\[1\].row\[8\].yc/uin[1] blk.column\[1\].row\[7\].yc/hempty blk.column\[0\].row\[7\].yc/lempty
+ blk.column\[1\].row\[7\].yc/lempty blk.column\[1\].row\[7\].yc/lin[0] blk.column\[1\].row\[7\].yc/lin[1]
+ blk.column\[2\].row\[7\].yc/rin[0] blk.column\[2\].row\[7\].yc/rin[1] blk.column\[0\].row\[7\].yc/hempty
+ blk.column\[1\].row\[7\].yc/reset blk.column\[1\].row\[8\].yc/reset blk.column\[1\].row\[7\].yc/rin[0]
+ blk.column\[1\].row\[7\].yc/rin[1] blk.column\[0\].row\[7\].yc/lin[0] blk.column\[0\].row\[7\].yc/lin[1]
+ blk.column\[1\].row\[7\].yc/uempty blk.column\[1\].row\[7\].yc/uin[0] blk.column\[1\].row\[7\].yc/uin[1]
+ blk.column\[1\].row\[6\].yc/din[0] blk.column\[1\].row\[6\].yc/din[1] blk.column\[1\].row\[6\].yc/dempty
+ blk.column\[1\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_484_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_484_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_267_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_274_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_496_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_800_ wb_clk_i _800_/D VGND VGND VPWR VPWR _314_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_44_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_731_ VGND VGND VPWR VPWR _731_/HI la_data_out[115] sky130_fd_sc_hd__conb_1
XFILLER_152_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_662_ VGND VGND VPWR VPWR _662_/HI io_out[36] sky130_fd_sc_hd__conb_1
XPHY_6677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_362_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_507_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_593_ VGND VGND VPWR VPWR _593_/HI io_oeb[5] sky130_fd_sc_hd__conb_1
XFILLER_496_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_420_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_385_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_535_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_535_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[0\].yc la_data_in[111] blk.column\[15\].row\[1\].yc/cbitin
+ la_data_in[112] blk.column\[15\].row\[1\].yc/confclk blk.column\[15\].row\[0\].yc/dempty
+ blk.column\[15\].row\[0\].yc/din[0] blk.column\[15\].row\[0\].yc/din[1] blk.column\[15\].row\[1\].yc/uin[0]
+ blk.column\[15\].row\[1\].yc/uin[1] blk.column\[15\].row\[0\].yc/hempty blk.column\[14\].row\[0\].yc/lempty
+ _450_/HI _526_/LO _527_/LO blk.column\[15\].row\[0\].yc/lout[0] blk.column\[15\].row\[0\].yc/lout[1]
+ blk.column\[14\].row\[0\].yc/hempty la_data_in[113] blk.column\[15\].row\[1\].yc/reset
+ blk.column\[15\].row\[0\].yc/rin[0] blk.column\[15\].row\[0\].yc/rin[1] blk.column\[14\].row\[0\].yc/lin[0]
+ blk.column\[14\].row\[0\].yc/lin[1] _528_/LO la_data_in[94] la_data_in[95] la_data_out[30]
+ la_data_out[31] blk.column\[15\].row\[0\].yc/vempty blk.column\[15\].row\[1\].yc/uempty
+ VPWR VGND ycell
XFILLER_68_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_531_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_364_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[1\].yc blk.column\[6\].row\[1\].yc/cbitin blk.column\[6\].row\[2\].yc/cbitin
+ blk.column\[6\].row\[1\].yc/confclk blk.column\[6\].row\[2\].yc/confclk blk.column\[6\].row\[1\].yc/dempty
+ blk.column\[6\].row\[1\].yc/din[0] blk.column\[6\].row\[1\].yc/din[1] blk.column\[6\].row\[2\].yc/uin[0]
+ blk.column\[6\].row\[2\].yc/uin[1] blk.column\[6\].row\[1\].yc/hempty blk.column\[5\].row\[1\].yc/lempty
+ blk.column\[6\].row\[1\].yc/lempty blk.column\[6\].row\[1\].yc/lin[0] blk.column\[6\].row\[1\].yc/lin[1]
+ blk.column\[7\].row\[1\].yc/rin[0] blk.column\[7\].row\[1\].yc/rin[1] blk.column\[5\].row\[1\].yc/hempty
+ blk.column\[6\].row\[1\].yc/reset blk.column\[6\].row\[2\].yc/reset blk.column\[6\].row\[1\].yc/rin[0]
+ blk.column\[6\].row\[1\].yc/rin[1] blk.column\[5\].row\[1\].yc/lin[0] blk.column\[5\].row\[1\].yc/lin[1]
+ blk.column\[6\].row\[1\].yc/uempty blk.column\[6\].row\[1\].yc/uin[0] blk.column\[6\].row\[1\].yc/uin[1]
+ blk.column\[6\].row\[0\].yc/din[0] blk.column\[6\].row\[0\].yc/din[1] blk.column\[6\].row\[0\].yc/dempty
+ blk.column\[6\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_522_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_520_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_451_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_351_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_380_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_402_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_506_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_401_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_327_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_519_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_714_ VGND VGND VPWR VPWR _714_/HI la_data_out[98] sky130_fd_sc_hd__conb_1
XFILLER_166_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_251_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_645_ VGND VGND VPWR VPWR _645_/HI io_out[19] sky130_fd_sc_hd__conb_1
XPHY_5762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_389_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_576_ VGND VGND VPWR VPWR _576_/HI _576_/LO sky130_fd_sc_hd__conb_1
XFILLER_400_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_515_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[11\].yc blk.column\[10\].row\[11\].yc/cbitin blk.column\[10\].row\[12\].yc/cbitin
+ blk.column\[10\].row\[11\].yc/confclk blk.column\[10\].row\[12\].yc/confclk blk.column\[10\].row\[11\].yc/dempty
+ blk.column\[10\].row\[11\].yc/din[0] blk.column\[10\].row\[11\].yc/din[1] blk.column\[10\].row\[12\].yc/uin[0]
+ blk.column\[10\].row\[12\].yc/uin[1] blk.column\[10\].row\[11\].yc/hempty blk.column\[9\].row\[11\].yc/lempty
+ blk.column\[10\].row\[11\].yc/lempty blk.column\[10\].row\[11\].yc/lin[0] blk.column\[10\].row\[11\].yc/lin[1]
+ blk.column\[11\].row\[11\].yc/rin[0] blk.column\[11\].row\[11\].yc/rin[1] blk.column\[9\].row\[11\].yc/hempty
+ blk.column\[10\].row\[11\].yc/reset blk.column\[10\].row\[12\].yc/reset blk.column\[9\].row\[11\].yc/lout[0]
+ blk.column\[9\].row\[11\].yc/lout[1] blk.column\[9\].row\[11\].yc/lin[0] blk.column\[9\].row\[11\].yc/lin[1]
+ blk.column\[10\].row\[11\].yc/uempty blk.column\[10\].row\[11\].yc/uin[0] blk.column\[10\].row\[11\].yc/uin[1]
+ blk.column\[10\].row\[10\].yc/din[0] blk.column\[10\].row\[10\].yc/din[1] blk.column\[10\].row\[10\].yc/dempty
+ blk.column\[10\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_509_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_299_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_320_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_495_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_492_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_451_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_490_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_430_ VGND VGND VPWR VPWR _430_/HI _430_/LO sky130_fd_sc_hd__conb_1
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_361_ _361_/A VGND VGND VPWR VPWR _361_/X sky130_fd_sc_hd__buf_2
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_521_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_393_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_315_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_485_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_343_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[8\].yc blk.column\[11\].row\[8\].yc/cbitin blk.column\[11\].row\[9\].yc/cbitin
+ blk.column\[11\].row\[8\].yc/confclk blk.column\[11\].row\[9\].yc/confclk blk.column\[11\].row\[8\].yc/dempty
+ blk.column\[11\].row\[8\].yc/din[0] blk.column\[11\].row\[8\].yc/din[1] blk.column\[11\].row\[9\].yc/uin[0]
+ blk.column\[11\].row\[9\].yc/uin[1] blk.column\[11\].row\[8\].yc/hempty blk.column\[10\].row\[8\].yc/lempty
+ blk.column\[11\].row\[8\].yc/lempty blk.column\[11\].row\[8\].yc/lin[0] blk.column\[11\].row\[8\].yc/lin[1]
+ blk.column\[12\].row\[8\].yc/rin[0] blk.column\[12\].row\[8\].yc/rin[1] blk.column\[10\].row\[8\].yc/hempty
+ blk.column\[11\].row\[8\].yc/reset blk.column\[11\].row\[9\].yc/reset blk.column\[11\].row\[8\].yc/rin[0]
+ blk.column\[11\].row\[8\].yc/rin[1] blk.column\[10\].row\[8\].yc/lin[0] blk.column\[10\].row\[8\].yc/lin[1]
+ blk.column\[11\].row\[8\].yc/uempty blk.column\[11\].row\[8\].yc/uin[0] blk.column\[11\].row\[8\].yc/uin[1]
+ blk.column\[11\].row\[7\].yc/din[0] blk.column\[11\].row\[7\].yc/din[1] blk.column\[11\].row\[7\].yc/dempty
+ blk.column\[11\].row\[9\].yc/uempty VPWR VGND ycell
X_628_ VGND VGND VPWR VPWR _628_/HI io_out[2] sky130_fd_sc_hd__conb_1
XFILLER_526_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_559_ VGND VGND VPWR VPWR _559_/HI _559_/LO sky130_fd_sc_hd__conb_1
XFILLER_359_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_534_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[9\].yc blk.column\[2\].row\[9\].yc/cbitin blk.column\[2\].row\[9\].yc/cbitout
+ blk.column\[2\].row\[9\].yc/confclk blk.column\[2\].row\[9\].yc/confclko blk.column\[2\].row\[9\].yc/dempty
+ blk.column\[2\].row\[9\].yc/din[0] blk.column\[2\].row\[9\].yc/din[1] blk.column\[2\].row\[9\].yc/dout[0]
+ blk.column\[2\].row\[9\].yc/dout[1] blk.column\[2\].row\[9\].yc/hempty blk.column\[1\].row\[9\].yc/lempty
+ blk.column\[2\].row\[9\].yc/lempty blk.column\[2\].row\[9\].yc/lin[0] blk.column\[2\].row\[9\].yc/lin[1]
+ blk.column\[3\].row\[9\].yc/rin[0] blk.column\[3\].row\[9\].yc/rin[1] blk.column\[1\].row\[9\].yc/hempty
+ blk.column\[2\].row\[9\].yc/reset blk.column\[2\].row\[9\].yc/reseto blk.column\[2\].row\[9\].yc/rin[0]
+ blk.column\[2\].row\[9\].yc/rin[1] blk.column\[1\].row\[9\].yc/lin[0] blk.column\[1\].row\[9\].yc/lin[1]
+ blk.column\[2\].row\[9\].yc/uempty blk.column\[2\].row\[9\].yc/uin[0] blk.column\[2\].row\[9\].yc/uin[1]
+ blk.column\[2\].row\[8\].yc/din[0] blk.column\[2\].row\[8\].yc/din[1] blk.column\[2\].row\[8\].yc/dempty
+ blk.column\[2\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_172_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[12\].yc blk.column\[7\].row\[12\].yc/cbitin blk.column\[7\].row\[13\].yc/cbitin
+ blk.column\[7\].row\[12\].yc/confclk blk.column\[7\].row\[13\].yc/confclk blk.column\[7\].row\[12\].yc/dempty
+ blk.column\[7\].row\[12\].yc/din[0] blk.column\[7\].row\[12\].yc/din[1] blk.column\[7\].row\[13\].yc/uin[0]
+ blk.column\[7\].row\[13\].yc/uin[1] blk.column\[7\].row\[12\].yc/hempty blk.column\[6\].row\[12\].yc/lempty
+ blk.column\[7\].row\[12\].yc/lempty blk.column\[7\].row\[12\].yc/lin[0] blk.column\[7\].row\[12\].yc/lin[1]
+ blk.column\[8\].row\[12\].yc/rin[0] blk.column\[8\].row\[12\].yc/rin[1] blk.column\[6\].row\[12\].yc/hempty
+ blk.column\[7\].row\[12\].yc/reset blk.column\[7\].row\[13\].yc/reset blk.column\[7\].row\[12\].yc/rin[0]
+ blk.column\[7\].row\[12\].yc/rin[1] blk.column\[6\].row\[12\].yc/lin[0] blk.column\[6\].row\[12\].yc/lin[1]
+ blk.column\[7\].row\[12\].yc/uempty blk.column\[7\].row\[12\].yc/uin[0] blk.column\[7\].row\[12\].yc/uin[1]
+ blk.column\[7\].row\[11\].yc/din[0] blk.column\[7\].row\[11\].yc/din[1] blk.column\[7\].row\[11\].yc/dempty
+ blk.column\[7\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_160_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_541_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_431_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_369_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_503_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_384_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_492_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_259_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_275_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_352_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_533_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_413_ _412_/X wbs_dat_o[10] _330_/A _410_/X VGND VGND VPWR VPWR _754_/D sky130_fd_sc_hd__o22a_4
XFILLER_14_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_540_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_344_ _344_/A VGND VGND VPWR VPWR _344_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_343_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[3\].yc blk.column\[7\].row\[3\].yc/cbitin blk.column\[7\].row\[4\].yc/cbitin
+ blk.column\[7\].row\[3\].yc/confclk blk.column\[7\].row\[4\].yc/confclk blk.column\[7\].row\[3\].yc/dempty
+ blk.column\[7\].row\[3\].yc/din[0] blk.column\[7\].row\[3\].yc/din[1] blk.column\[7\].row\[4\].yc/uin[0]
+ blk.column\[7\].row\[4\].yc/uin[1] blk.column\[7\].row\[3\].yc/hempty blk.column\[6\].row\[3\].yc/lempty
+ blk.column\[7\].row\[3\].yc/lempty blk.column\[7\].row\[3\].yc/lin[0] blk.column\[7\].row\[3\].yc/lin[1]
+ blk.column\[8\].row\[3\].yc/rin[0] blk.column\[8\].row\[3\].yc/rin[1] blk.column\[6\].row\[3\].yc/hempty
+ blk.column\[7\].row\[3\].yc/reset blk.column\[7\].row\[4\].yc/reset blk.column\[7\].row\[3\].yc/rin[0]
+ blk.column\[7\].row\[3\].yc/rin[1] blk.column\[6\].row\[3\].yc/lin[0] blk.column\[6\].row\[3\].yc/lin[1]
+ blk.column\[7\].row\[3\].yc/uempty blk.column\[7\].row\[3\].yc/uin[0] blk.column\[7\].row\[3\].yc/uin[1]
+ blk.column\[7\].row\[2\].yc/din[0] blk.column\[7\].row\[2\].yc/din[1] blk.column\[7\].row\[2\].yc/dempty
+ blk.column\[7\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_482_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_485_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_508_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_517_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_389_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3029 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_511_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_392_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_522_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_369_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_499_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_372_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_513_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_353_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_392_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_3206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_483_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[14\].yc blk.column\[14\].row\[14\].yc/cbitin blk.column\[14\].row\[15\].yc/cbitin
+ blk.column\[14\].row\[14\].yc/confclk blk.column\[14\].row\[15\].yc/confclk blk.column\[14\].row\[14\].yc/dempty
+ blk.column\[14\].row\[14\].yc/din[0] blk.column\[14\].row\[14\].yc/din[1] blk.column\[14\].row\[15\].yc/uin[0]
+ blk.column\[14\].row\[15\].yc/uin[1] blk.column\[14\].row\[14\].yc/hempty blk.column\[13\].row\[14\].yc/lempty
+ blk.column\[14\].row\[14\].yc/lempty blk.column\[14\].row\[14\].yc/lin[0] blk.column\[14\].row\[14\].yc/lin[1]
+ blk.column\[15\].row\[14\].yc/rin[0] blk.column\[15\].row\[14\].yc/rin[1] blk.column\[13\].row\[14\].yc/hempty
+ blk.column\[14\].row\[14\].yc/reset blk.column\[14\].row\[15\].yc/reset blk.column\[14\].row\[14\].yc/rin[0]
+ blk.column\[14\].row\[14\].yc/rin[1] blk.column\[13\].row\[14\].yc/lin[0] blk.column\[13\].row\[14\].yc/lin[1]
+ blk.column\[14\].row\[14\].yc/uempty blk.column\[14\].row\[14\].yc/uin[0] blk.column\[14\].row\[14\].yc/uin[1]
+ blk.column\[14\].row\[13\].yc/din[0] blk.column\[14\].row\[13\].yc/din[1] blk.column\[14\].row\[13\].yc/dempty
+ blk.column\[14\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_21_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_327_ _326_/Y _324_/X wbs_dat_i[12] _324_/X VGND VGND VPWR VPWR _327_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_509_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_486_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_263_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_504_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_366_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_322_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_487_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_344_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_238_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_390_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_490_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_447_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_450_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_411_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_327_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_442_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_399_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_336_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_242_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_386_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_528_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_730_ VGND VGND VPWR VPWR _730_/HI la_data_out[114] sky130_fd_sc_hd__conb_1
XFILLER_131_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_661_ VGND VGND VPWR VPWR _661_/HI io_out[35] sky130_fd_sc_hd__conb_1
XFILLER_526_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_508_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_592_ VGND VGND VPWR VPWR _592_/HI io_oeb[4] sky130_fd_sc_hd__conb_1
XPHY_5966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_355_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_385_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[8\].row\[5\].yc blk.column\[8\].row\[5\].yc/cbitin blk.column\[8\].row\[6\].yc/cbitin
+ blk.column\[8\].row\[5\].yc/confclk blk.column\[8\].row\[6\].yc/confclk blk.column\[8\].row\[5\].yc/dempty
+ blk.column\[8\].row\[5\].yc/din[0] blk.column\[8\].row\[5\].yc/din[1] blk.column\[8\].row\[6\].yc/uin[0]
+ blk.column\[8\].row\[6\].yc/uin[1] blk.column\[8\].row\[5\].yc/hempty blk.column\[7\].row\[5\].yc/lempty
+ blk.column\[8\].row\[5\].yc/lempty blk.column\[8\].row\[5\].yc/lin[0] blk.column\[8\].row\[5\].yc/lin[1]
+ blk.column\[9\].row\[5\].yc/rin[0] blk.column\[9\].row\[5\].yc/rin[1] blk.column\[7\].row\[5\].yc/hempty
+ blk.column\[8\].row\[5\].yc/reset blk.column\[8\].row\[6\].yc/reset blk.column\[8\].row\[5\].yc/rin[0]
+ blk.column\[8\].row\[5\].yc/rin[1] blk.column\[7\].row\[5\].yc/lin[0] blk.column\[7\].row\[5\].yc/lin[1]
+ blk.column\[8\].row\[5\].yc/uempty blk.column\[8\].row\[5\].yc/uin[0] blk.column\[8\].row\[5\].yc/uin[1]
+ blk.column\[8\].row\[4\].yc/din[0] blk.column\[8\].row\[4\].yc/din[1] blk.column\[8\].row\[4\].yc/dempty
+ blk.column\[8\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_535_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_502_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_531_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_364_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_483_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_520_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[2\].row\[13\].yc blk.column\[2\].row\[13\].yc/cbitin blk.column\[2\].row\[14\].yc/cbitin
+ blk.column\[2\].row\[13\].yc/confclk blk.column\[2\].row\[14\].yc/confclk blk.column\[2\].row\[13\].yc/dempty
+ blk.column\[2\].row\[13\].yc/din[0] blk.column\[2\].row\[13\].yc/din[1] blk.column\[2\].row\[14\].yc/uin[0]
+ blk.column\[2\].row\[14\].yc/uin[1] blk.column\[2\].row\[13\].yc/hempty blk.column\[1\].row\[13\].yc/lempty
+ blk.column\[2\].row\[13\].yc/lempty blk.column\[2\].row\[13\].yc/lin[0] blk.column\[2\].row\[13\].yc/lin[1]
+ blk.column\[3\].row\[13\].yc/rin[0] blk.column\[3\].row\[13\].yc/rin[1] blk.column\[1\].row\[13\].yc/hempty
+ blk.column\[2\].row\[13\].yc/reset blk.column\[2\].row\[14\].yc/reset blk.column\[2\].row\[13\].yc/rin[0]
+ blk.column\[2\].row\[13\].yc/rin[1] blk.column\[1\].row\[13\].yc/lin[0] blk.column\[1\].row\[13\].yc/lin[1]
+ blk.column\[2\].row\[13\].yc/uempty blk.column\[2\].row\[13\].yc/uin[0] blk.column\[2\].row\[13\].yc/uin[1]
+ blk.column\[2\].row\[12\].yc/din[0] blk.column\[2\].row\[12\].yc/din[1] blk.column\[2\].row\[12\].yc/dempty
+ blk.column\[2\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_258_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_457_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_334_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_406_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_402_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_440_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_472_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_713_ VGND VGND VPWR VPWR _713_/HI la_data_out[97] sky130_fd_sc_hd__conb_1
XPHY_7187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_644_ VGND VGND VPWR VPWR _644_/HI io_out[18] sky130_fd_sc_hd__conb_1
XPHY_6486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_389_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_575_ VGND VGND VPWR VPWR _575_/HI _575_/LO sky130_fd_sc_hd__conb_1
XPHY_5796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_537_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_430_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_360_ _359_/X VGND VGND VPWR VPWR _361_/A sky130_fd_sc_hd__buf_2
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_495_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_354_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_318_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_428_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_471_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_10953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_343_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_627_ VGND VGND VPWR VPWR _627_/HI io_out[1] sky130_fd_sc_hd__conb_1
XFILLER_402_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_378_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_558_ VGND VGND VPWR VPWR _558_/HI _558_/LO sky130_fd_sc_hd__conb_1
XFILLER_539_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_474_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_489_ VGND VGND VPWR VPWR _489_/HI _489_/LO sky130_fd_sc_hd__conb_1
XFILLER_439_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_349_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_475_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_396_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_503_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_352_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_412_ _419_/A VGND VGND VPWR VPWR _412_/X sky130_fd_sc_hd__buf_2
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[9\].row\[7\].yc blk.column\[9\].row\[7\].yc/cbitin blk.column\[9\].row\[8\].yc/cbitin
+ blk.column\[9\].row\[7\].yc/confclk blk.column\[9\].row\[8\].yc/confclk blk.column\[9\].row\[7\].yc/dempty
+ blk.column\[9\].row\[7\].yc/din[0] blk.column\[9\].row\[7\].yc/din[1] blk.column\[9\].row\[8\].yc/uin[0]
+ blk.column\[9\].row\[8\].yc/uin[1] blk.column\[9\].row\[7\].yc/hempty blk.column\[8\].row\[7\].yc/lempty
+ blk.column\[9\].row\[7\].yc/lempty blk.column\[9\].row\[7\].yc/lin[0] blk.column\[9\].row\[7\].yc/lin[1]
+ blk.column\[9\].row\[7\].yc/lout[0] blk.column\[9\].row\[7\].yc/lout[1] blk.column\[8\].row\[7\].yc/hempty
+ blk.column\[9\].row\[7\].yc/reset blk.column\[9\].row\[8\].yc/reset blk.column\[9\].row\[7\].yc/rin[0]
+ blk.column\[9\].row\[7\].yc/rin[1] blk.column\[8\].row\[7\].yc/lin[0] blk.column\[8\].row\[7\].yc/lin[1]
+ blk.column\[9\].row\[7\].yc/uempty blk.column\[9\].row\[7\].yc/uin[0] blk.column\[9\].row\[7\].yc/uin[1]
+ blk.column\[9\].row\[6\].yc/din[0] blk.column\[9\].row\[6\].yc/din[1] blk.column\[9\].row\[6\].yc/dempty
+ blk.column\[9\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_501_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_343_ _342_/Y _340_/X wbs_dat_i[22] _340_/X VGND VGND VPWR VPWR _790_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_528_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_511_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_383_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_481_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_270_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_418_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_527_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_333_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_516_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_483_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_429_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_395_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_326_ _326_/A VGND VGND VPWR VPWR _326_/Y sky130_fd_sc_hd__inv_2
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_517_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_531_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_517_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[0\].yc la_data_in[100] blk.column\[4\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[4\].row\[1\].yc/confclk blk.column\[4\].row\[0\].yc/dempty blk.column\[4\].row\[0\].yc/din[0]
+ blk.column\[4\].row\[0\].yc/din[1] blk.column\[4\].row\[1\].yc/uin[0] blk.column\[4\].row\[1\].yc/uin[1]
+ blk.column\[4\].row\[0\].yc/hempty blk.column\[3\].row\[0\].yc/lempty blk.column\[4\].row\[0\].yc/lempty
+ blk.column\[4\].row\[0\].yc/lin[0] blk.column\[4\].row\[0\].yc/lin[1] blk.column\[5\].row\[0\].yc/rin[0]
+ blk.column\[5\].row\[0\].yc/rin[1] blk.column\[3\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[4\].row\[1\].yc/reset blk.column\[4\].row\[0\].yc/rin[0] blk.column\[4\].row\[0\].yc/rin[1]
+ blk.column\[3\].row\[0\].yc/lin[0] blk.column\[3\].row\[0\].yc/lin[1] _570_/LO la_data_in[72]
+ la_data_in[73] la_data_out[8] la_data_out[9] blk.column\[4\].row\[0\].yc/vempty
+ blk.column\[4\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[11\].row\[10\].yc blk.column\[11\].row\[9\].yc/cbitout blk.column\[11\].row\[11\].yc/cbitin
+ blk.column\[11\].row\[9\].yc/confclko blk.column\[11\].row\[11\].yc/confclk blk.column\[11\].row\[10\].yc/dempty
+ blk.column\[11\].row\[10\].yc/din[0] blk.column\[11\].row\[10\].yc/din[1] blk.column\[11\].row\[11\].yc/uin[0]
+ blk.column\[11\].row\[11\].yc/uin[1] blk.column\[11\].row\[10\].yc/hempty blk.column\[10\].row\[10\].yc/lempty
+ blk.column\[11\].row\[10\].yc/lempty blk.column\[11\].row\[10\].yc/lin[0] blk.column\[11\].row\[10\].yc/lin[1]
+ blk.column\[12\].row\[10\].yc/rin[0] blk.column\[12\].row\[10\].yc/rin[1] blk.column\[10\].row\[10\].yc/hempty
+ blk.column\[11\].row\[9\].yc/reseto blk.column\[11\].row\[11\].yc/reset blk.column\[11\].row\[10\].yc/rin[0]
+ blk.column\[11\].row\[10\].yc/rin[1] blk.column\[10\].row\[10\].yc/lin[0] blk.column\[10\].row\[10\].yc/lin[1]
+ blk.column\[11\].row\[9\].yc/vempty2 blk.column\[11\].row\[9\].yc/dout[0] blk.column\[11\].row\[9\].yc/dout[1]
+ blk.column\[11\].row\[9\].yc/din[0] blk.column\[11\].row\[9\].yc/din[1] blk.column\[11\].row\[9\].yc/dempty
+ blk.column\[11\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_512_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_476_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_409_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_383_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_363_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_345_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_390_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_300_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_332_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_442_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_499_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_309_ _802_/Q VGND VGND VPWR VPWR _309_/Y sky130_fd_sc_hd__inv_2
XFILLER_536_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_256_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_505_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_421_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_225_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_507_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_339_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_517_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[11\].yc blk.column\[8\].row\[11\].yc/cbitin blk.column\[8\].row\[12\].yc/cbitin
+ blk.column\[8\].row\[11\].yc/confclk blk.column\[8\].row\[12\].yc/confclk blk.column\[8\].row\[11\].yc/dempty
+ blk.column\[8\].row\[11\].yc/din[0] blk.column\[8\].row\[11\].yc/din[1] blk.column\[8\].row\[12\].yc/uin[0]
+ blk.column\[8\].row\[12\].yc/uin[1] blk.column\[8\].row\[11\].yc/hempty blk.column\[7\].row\[11\].yc/lempty
+ blk.column\[8\].row\[11\].yc/lempty blk.column\[8\].row\[11\].yc/lin[0] blk.column\[8\].row\[11\].yc/lin[1]
+ blk.column\[9\].row\[11\].yc/rin[0] blk.column\[9\].row\[11\].yc/rin[1] blk.column\[7\].row\[11\].yc/hempty
+ blk.column\[8\].row\[11\].yc/reset blk.column\[8\].row\[12\].yc/reset blk.column\[8\].row\[11\].yc/rin[0]
+ blk.column\[8\].row\[11\].yc/rin[1] blk.column\[7\].row\[11\].yc/lin[0] blk.column\[7\].row\[11\].yc/lin[1]
+ blk.column\[8\].row\[11\].yc/uempty blk.column\[8\].row\[11\].yc/uin[0] blk.column\[8\].row\[11\].yc/uin[1]
+ blk.column\[8\].row\[10\].yc/din[0] blk.column\[8\].row\[10\].yc/din[1] blk.column\[8\].row\[10\].yc/dempty
+ blk.column\[8\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_161_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_660_ VGND VGND VPWR VPWR _660_/HI io_out[34] sky130_fd_sc_hd__conb_1
XPHY_6646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_591_ VGND VGND VPWR VPWR _591_/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_502_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_524_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_515_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_433_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_253_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_470_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_327_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_789_ wb_clk_i _789_/D VGND VGND VPWR VPWR _344_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_143_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_525_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_531_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[8\].yc blk.column\[0\].row\[8\].yc/cbitin blk.column\[0\].row\[9\].yc/cbitin
+ blk.column\[0\].row\[8\].yc/confclk blk.column\[0\].row\[9\].yc/confclk blk.column\[0\].row\[8\].yc/dempty
+ blk.column\[0\].row\[8\].yc/din[0] blk.column\[0\].row\[8\].yc/din[1] blk.column\[0\].row\[9\].yc/uin[0]
+ blk.column\[0\].row\[9\].yc/uin[1] blk.column\[0\].row\[8\].yc/hempty blk.column\[0\].row\[8\].yc/hempty2
+ blk.column\[0\].row\[8\].yc/lempty blk.column\[0\].row\[8\].yc/lin[0] blk.column\[0\].row\[8\].yc/lin[1]
+ blk.column\[1\].row\[8\].yc/rin[0] blk.column\[1\].row\[8\].yc/rin[1] _443_/HI blk.column\[0\].row\[8\].yc/reset
+ blk.column\[0\].row\[9\].yc/reset _507_/LO _508_/LO blk.column\[0\].row\[8\].yc/rout[0]
+ blk.column\[0\].row\[8\].yc/rout[1] blk.column\[0\].row\[8\].yc/uempty blk.column\[0\].row\[8\].yc/uin[0]
+ blk.column\[0\].row\[8\].yc/uin[1] blk.column\[0\].row\[7\].yc/din[0] blk.column\[0\].row\[7\].yc/din[1]
+ blk.column\[0\].row\[7\].yc/dempty blk.column\[0\].row\[9\].yc/uempty VPWR VGND
+ ycell
XPHY_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_360_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_402_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_495_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_428_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_389_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_712_ VGND VGND VPWR VPWR _712_/HI la_data_out[96] sky130_fd_sc_hd__conb_1
XPHY_7177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_643_ VGND VGND VPWR VPWR _643_/HI io_out[17] sky130_fd_sc_hd__conb_1
XPHY_6487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_574_ VGND VGND VPWR VPWR _574_/HI _574_/LO sky130_fd_sc_hd__conb_1
XPHY_5797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_396_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_508_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_507_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xblk.column\[14\].row\[1\].yc blk.column\[14\].row\[1\].yc/cbitin blk.column\[14\].row\[2\].yc/cbitin
+ blk.column\[14\].row\[1\].yc/confclk blk.column\[14\].row\[2\].yc/confclk blk.column\[14\].row\[1\].yc/dempty
+ blk.column\[14\].row\[1\].yc/din[0] blk.column\[14\].row\[1\].yc/din[1] blk.column\[14\].row\[2\].yc/uin[0]
+ blk.column\[14\].row\[2\].yc/uin[1] blk.column\[14\].row\[1\].yc/hempty blk.column\[13\].row\[1\].yc/lempty
+ blk.column\[14\].row\[1\].yc/lempty blk.column\[14\].row\[1\].yc/lin[0] blk.column\[14\].row\[1\].yc/lin[1]
+ blk.column\[15\].row\[1\].yc/rin[0] blk.column\[15\].row\[1\].yc/rin[1] blk.column\[13\].row\[1\].yc/hempty
+ blk.column\[14\].row\[1\].yc/reset blk.column\[14\].row\[2\].yc/reset blk.column\[14\].row\[1\].yc/rin[0]
+ blk.column\[14\].row\[1\].yc/rin[1] blk.column\[13\].row\[1\].yc/lin[0] blk.column\[13\].row\[1\].yc/lin[1]
+ blk.column\[14\].row\[1\].yc/uempty blk.column\[14\].row\[1\].yc/uin[0] blk.column\[14\].row\[1\].yc/uin[1]
+ blk.column\[14\].row\[0\].yc/din[0] blk.column\[14\].row\[0\].yc/din[1] blk.column\[14\].row\[0\].yc/dempty
+ blk.column\[14\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_286_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[13\].yc blk.column\[15\].row\[13\].yc/cbitin blk.column\[15\].row\[14\].yc/cbitin
+ blk.column\[15\].row\[13\].yc/confclk blk.column\[15\].row\[14\].yc/confclk blk.column\[15\].row\[13\].yc/dempty
+ blk.column\[15\].row\[13\].yc/din[0] blk.column\[15\].row\[13\].yc/din[1] blk.column\[15\].row\[14\].yc/uin[0]
+ blk.column\[15\].row\[14\].yc/uin[1] blk.column\[15\].row\[13\].yc/hempty blk.column\[14\].row\[13\].yc/lempty
+ _454_/HI _535_/LO _536_/LO blk.column\[15\].row\[13\].yc/lout[0] blk.column\[15\].row\[13\].yc/lout[1]
+ blk.column\[14\].row\[13\].yc/hempty blk.column\[15\].row\[13\].yc/reset blk.column\[15\].row\[14\].yc/reset
+ blk.column\[15\].row\[13\].yc/rin[0] blk.column\[15\].row\[13\].yc/rin[1] blk.column\[14\].row\[13\].yc/lin[0]
+ blk.column\[14\].row\[13\].yc/lin[1] blk.column\[15\].row\[13\].yc/uempty blk.column\[15\].row\[13\].yc/uin[0]
+ blk.column\[15\].row\[13\].yc/uin[1] blk.column\[15\].row\[12\].yc/din[0] blk.column\[15\].row\[12\].yc/din[1]
+ blk.column\[15\].row\[12\].yc/dempty blk.column\[15\].row\[14\].yc/uempty VPWR VGND
+ ycell
XFILLER_149_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_428_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[2\].yc blk.column\[5\].row\[2\].yc/cbitin blk.column\[5\].row\[3\].yc/cbitin
+ blk.column\[5\].row\[2\].yc/confclk blk.column\[5\].row\[3\].yc/confclk blk.column\[5\].row\[2\].yc/dempty
+ blk.column\[5\].row\[2\].yc/din[0] blk.column\[5\].row\[2\].yc/din[1] blk.column\[5\].row\[3\].yc/uin[0]
+ blk.column\[5\].row\[3\].yc/uin[1] blk.column\[5\].row\[2\].yc/hempty blk.column\[4\].row\[2\].yc/lempty
+ blk.column\[5\].row\[2\].yc/lempty blk.column\[5\].row\[2\].yc/lin[0] blk.column\[5\].row\[2\].yc/lin[1]
+ blk.column\[6\].row\[2\].yc/rin[0] blk.column\[6\].row\[2\].yc/rin[1] blk.column\[4\].row\[2\].yc/hempty
+ blk.column\[5\].row\[2\].yc/reset blk.column\[5\].row\[3\].yc/reset blk.column\[5\].row\[2\].yc/rin[0]
+ blk.column\[5\].row\[2\].yc/rin[1] blk.column\[4\].row\[2\].yc/lin[0] blk.column\[4\].row\[2\].yc/lin[1]
+ blk.column\[5\].row\[2\].yc/uempty blk.column\[5\].row\[2\].yc/uin[0] blk.column\[5\].row\[2\].yc/uin[1]
+ blk.column\[5\].row\[1\].yc/din[0] blk.column\[5\].row\[1\].yc/din[1] blk.column\[5\].row\[1\].yc/dempty
+ blk.column\[5\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_503_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_514_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_423_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_402_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_213_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_328_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_626_ VGND VGND VPWR VPWR _626_/HI io_out[0] sky130_fd_sc_hd__conb_1
XFILLER_480_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_378_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_504_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_557_ VGND VGND VPWR VPWR _557_/HI _557_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_488_ VGND VGND VPWR VPWR _488_/HI _488_/LO sky130_fd_sc_hd__conb_1
XFILLER_294_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_439_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_267_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_347_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_411_ _405_/X wbs_dat_o[11] _795_/Q _410_/X VGND VGND VPWR VPWR _411_/X sky130_fd_sc_hd__o22a_4
XFILLER_19_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_262_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_342_ _790_/Q VGND VGND VPWR VPWR _342_/Y sky130_fd_sc_hd__inv_2
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_457_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_441_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_609_ VGND VGND VPWR VPWR _609_/HI io_oeb[21] sky130_fd_sc_hd__conb_1
XFILLER_523_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[9\].yc blk.column\[10\].row\[9\].yc/cbitin blk.column\[10\].row\[9\].yc/cbitout
+ blk.column\[10\].row\[9\].yc/confclk blk.column\[10\].row\[9\].yc/confclko blk.column\[10\].row\[9\].yc/dempty
+ blk.column\[10\].row\[9\].yc/din[0] blk.column\[10\].row\[9\].yc/din[1] blk.column\[10\].row\[9\].yc/dout[0]
+ blk.column\[10\].row\[9\].yc/dout[1] blk.column\[10\].row\[9\].yc/hempty blk.column\[9\].row\[9\].yc/lempty
+ blk.column\[10\].row\[9\].yc/lempty blk.column\[10\].row\[9\].yc/lin[0] blk.column\[10\].row\[9\].yc/lin[1]
+ blk.column\[11\].row\[9\].yc/rin[0] blk.column\[11\].row\[9\].yc/rin[1] blk.column\[9\].row\[9\].yc/hempty
+ blk.column\[10\].row\[9\].yc/reset blk.column\[10\].row\[9\].yc/reseto blk.column\[9\].row\[9\].yc/lout[0]
+ blk.column\[9\].row\[9\].yc/lout[1] blk.column\[9\].row\[9\].yc/lin[0] blk.column\[9\].row\[9\].yc/lin[1]
+ blk.column\[10\].row\[9\].yc/uempty blk.column\[10\].row\[9\].yc/uin[0] blk.column\[10\].row\[9\].yc/uin[1]
+ blk.column\[10\].row\[8\].yc/din[0] blk.column\[10\].row\[8\].yc/din[1] blk.column\[10\].row\[8\].yc/dempty
+ blk.column\[10\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_14_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_517_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_487_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_485_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_270_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xblk.column\[3\].row\[12\].yc blk.column\[3\].row\[12\].yc/cbitin blk.column\[3\].row\[13\].yc/cbitin
+ blk.column\[3\].row\[12\].yc/confclk blk.column\[3\].row\[13\].yc/confclk blk.column\[3\].row\[12\].yc/dempty
+ blk.column\[3\].row\[12\].yc/din[0] blk.column\[3\].row\[12\].yc/din[1] blk.column\[3\].row\[13\].yc/uin[0]
+ blk.column\[3\].row\[13\].yc/uin[1] blk.column\[3\].row\[12\].yc/hempty blk.column\[2\].row\[12\].yc/lempty
+ blk.column\[3\].row\[12\].yc/lempty blk.column\[3\].row\[12\].yc/lin[0] blk.column\[3\].row\[12\].yc/lin[1]
+ blk.column\[4\].row\[12\].yc/rin[0] blk.column\[4\].row\[12\].yc/rin[1] blk.column\[2\].row\[12\].yc/hempty
+ blk.column\[3\].row\[12\].yc/reset blk.column\[3\].row\[13\].yc/reset blk.column\[3\].row\[12\].yc/rin[0]
+ blk.column\[3\].row\[12\].yc/rin[1] blk.column\[2\].row\[12\].yc/lin[0] blk.column\[2\].row\[12\].yc/lin[1]
+ blk.column\[3\].row\[12\].yc/uempty blk.column\[3\].row\[12\].yc/uin[0] blk.column\[3\].row\[12\].yc/uin[1]
+ blk.column\[3\].row\[11\].yc/din[0] blk.column\[3\].row\[11\].yc/din[1] blk.column\[3\].row\[11\].yc/dempty
+ blk.column\[3\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_522_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_502_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_454_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_429_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_483_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_360_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_395_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_375_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_325_ _323_/Y _319_/X wbs_dat_i[13] _324_/X VGND VGND VPWR VPWR _797_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_436_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xblk.column\[15\].row\[3\].yc blk.column\[15\].row\[3\].yc/cbitin blk.column\[15\].row\[4\].yc/cbitin
+ blk.column\[15\].row\[3\].yc/confclk blk.column\[15\].row\[4\].yc/confclk blk.column\[15\].row\[3\].yc/dempty
+ blk.column\[15\].row\[3\].yc/din[0] blk.column\[15\].row\[3\].yc/din[1] blk.column\[15\].row\[4\].yc/uin[0]
+ blk.column\[15\].row\[4\].yc/uin[1] blk.column\[15\].row\[3\].yc/hempty blk.column\[14\].row\[3\].yc/lempty
+ _460_/HI _547_/LO _548_/LO blk.column\[15\].row\[3\].yc/lout[0] blk.column\[15\].row\[3\].yc/lout[1]
+ blk.column\[14\].row\[3\].yc/hempty blk.column\[15\].row\[3\].yc/reset blk.column\[15\].row\[4\].yc/reset
+ blk.column\[15\].row\[3\].yc/rin[0] blk.column\[15\].row\[3\].yc/rin[1] blk.column\[14\].row\[3\].yc/lin[0]
+ blk.column\[14\].row\[3\].yc/lin[1] blk.column\[15\].row\[3\].yc/uempty blk.column\[15\].row\[3\].yc/uin[0]
+ blk.column\[15\].row\[3\].yc/uin[1] blk.column\[15\].row\[2\].yc/din[0] blk.column\[15\].row\[2\].yc/din[1]
+ blk.column\[15\].row\[2\].yc/dempty blk.column\[15\].row\[4\].yc/uempty VPWR VGND
+ ycell
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[6\].row\[4\].yc blk.column\[6\].row\[4\].yc/cbitin blk.column\[6\].row\[5\].yc/cbitin
+ blk.column\[6\].row\[4\].yc/confclk blk.column\[6\].row\[5\].yc/confclk blk.column\[6\].row\[4\].yc/dempty
+ blk.column\[6\].row\[4\].yc/din[0] blk.column\[6\].row\[4\].yc/din[1] blk.column\[6\].row\[5\].yc/uin[0]
+ blk.column\[6\].row\[5\].yc/uin[1] blk.column\[6\].row\[4\].yc/hempty blk.column\[5\].row\[4\].yc/lempty
+ blk.column\[6\].row\[4\].yc/lempty blk.column\[6\].row\[4\].yc/lin[0] blk.column\[6\].row\[4\].yc/lin[1]
+ blk.column\[7\].row\[4\].yc/rin[0] blk.column\[7\].row\[4\].yc/rin[1] blk.column\[5\].row\[4\].yc/hempty
+ blk.column\[6\].row\[4\].yc/reset blk.column\[6\].row\[5\].yc/reset blk.column\[6\].row\[4\].yc/rin[0]
+ blk.column\[6\].row\[4\].yc/rin[1] blk.column\[5\].row\[4\].yc/lin[0] blk.column\[5\].row\[4\].yc/lin[1]
+ blk.column\[6\].row\[4\].yc/uempty blk.column\[6\].row\[4\].yc/uin[0] blk.column\[6\].row\[4\].yc/uin[1]
+ blk.column\[6\].row\[3\].yc/din[0] blk.column\[6\].row\[3\].yc/din[1] blk.column\[6\].row\[3\].yc/dempty
+ blk.column\[6\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_438_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_476_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_436_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_383_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_417_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_502_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_297_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_528_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_327_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_332_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_442_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_520_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_308_ _307_/Y _303_/X wbs_dat_i[3] _303_/X VGND VGND VPWR VPWR _308_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_363_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[14\].yc blk.column\[10\].row\[14\].yc/cbitin blk.column\[10\].row\[15\].yc/cbitin
+ blk.column\[10\].row\[14\].yc/confclk blk.column\[10\].row\[15\].yc/confclk blk.column\[10\].row\[14\].yc/dempty
+ blk.column\[10\].row\[14\].yc/din[0] blk.column\[10\].row\[14\].yc/din[1] blk.column\[10\].row\[15\].yc/uin[0]
+ blk.column\[10\].row\[15\].yc/uin[1] blk.column\[10\].row\[14\].yc/hempty blk.column\[9\].row\[14\].yc/lempty
+ blk.column\[10\].row\[14\].yc/lempty blk.column\[10\].row\[14\].yc/lin[0] blk.column\[10\].row\[14\].yc/lin[1]
+ blk.column\[11\].row\[14\].yc/rin[0] blk.column\[11\].row\[14\].yc/rin[1] blk.column\[9\].row\[14\].yc/hempty
+ blk.column\[10\].row\[14\].yc/reset blk.column\[10\].row\[15\].yc/reset blk.column\[9\].row\[14\].yc/lout[0]
+ blk.column\[9\].row\[14\].yc/lout[1] blk.column\[9\].row\[14\].yc/lin[0] blk.column\[9\].row\[14\].yc/lin[1]
+ blk.column\[10\].row\[14\].yc/uempty blk.column\[10\].row\[14\].yc/uin[0] blk.column\[10\].row\[14\].yc/uin[1]
+ blk.column\[10\].row\[13\].yc/din[0] blk.column\[10\].row\[13\].yc/din[1] blk.column\[10\].row\[13\].yc/dempty
+ blk.column\[10\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_304_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_373_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_216_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_417_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_590_ VGND VGND VPWR VPWR _590_/HI io_oeb[2] sky130_fd_sc_hd__conb_1
XFILLER_524_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_521_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_298_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_788_ wb_clk_i _788_/D VGND VGND VPWR VPWR _347_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_56_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_490_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[15\].yc blk.column\[7\].row\[15\].yc/cbitin la_data_out[39]
+ blk.column\[7\].row\[15\].yc/confclk blk.column\[7\].row\[15\].yc/confclko _473_/HI
+ _580_/LO _581_/LO blk.column\[7\].row\[15\].yc/dout[0] blk.column\[7\].row\[15\].yc/dout[1]
+ blk.column\[7\].row\[15\].yc/hempty blk.column\[6\].row\[15\].yc/lempty blk.column\[7\].row\[15\].yc/lempty
+ blk.column\[7\].row\[15\].yc/lin[0] blk.column\[7\].row\[15\].yc/lin[1] blk.column\[8\].row\[15\].yc/rin[0]
+ blk.column\[8\].row\[15\].yc/rin[1] blk.column\[6\].row\[15\].yc/hempty blk.column\[7\].row\[15\].yc/reset
+ blk.column\[7\].row\[15\].yc/reseto blk.column\[7\].row\[15\].yc/rin[0] blk.column\[7\].row\[15\].yc/rin[1]
+ blk.column\[6\].row\[15\].yc/lin[0] blk.column\[6\].row\[15\].yc/lin[1] blk.column\[7\].row\[15\].yc/uempty
+ blk.column\[7\].row\[15\].yc/uin[0] blk.column\[7\].row\[15\].yc/uin[1] blk.column\[7\].row\[14\].yc/din[0]
+ blk.column\[7\].row\[14\].yc/din[1] blk.column\[7\].row\[14\].yc/dempty blk.column\[7\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_154_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_525_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_525_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_428_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_711_ VGND VGND VPWR VPWR _711_/HI la_data_out[95] sky130_fd_sc_hd__conb_1
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_460_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_642_ VGND VGND VPWR VPWR _642_/HI io_out[16] sky130_fd_sc_hd__conb_1
XPHY_6466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_360_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_573_ VGND VGND VPWR VPWR _573_/HI _573_/LO sky130_fd_sc_hd__conb_1
XFILLER_504_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_358_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_535_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_523_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[6\].yc blk.column\[7\].row\[6\].yc/cbitin blk.column\[7\].row\[7\].yc/cbitin
+ blk.column\[7\].row\[6\].yc/confclk blk.column\[7\].row\[7\].yc/confclk blk.column\[7\].row\[6\].yc/dempty
+ blk.column\[7\].row\[6\].yc/din[0] blk.column\[7\].row\[6\].yc/din[1] blk.column\[7\].row\[7\].yc/uin[0]
+ blk.column\[7\].row\[7\].yc/uin[1] blk.column\[7\].row\[6\].yc/hempty blk.column\[6\].row\[6\].yc/lempty
+ blk.column\[7\].row\[6\].yc/lempty blk.column\[7\].row\[6\].yc/lin[0] blk.column\[7\].row\[6\].yc/lin[1]
+ blk.column\[8\].row\[6\].yc/rin[0] blk.column\[8\].row\[6\].yc/rin[1] blk.column\[6\].row\[6\].yc/hempty
+ blk.column\[7\].row\[6\].yc/reset blk.column\[7\].row\[7\].yc/reset blk.column\[7\].row\[6\].yc/rin[0]
+ blk.column\[7\].row\[6\].yc/rin[1] blk.column\[6\].row\[6\].yc/lin[0] blk.column\[6\].row\[6\].yc/lin[1]
+ blk.column\[7\].row\[6\].yc/uempty blk.column\[7\].row\[6\].yc/uin[0] blk.column\[7\].row\[6\].yc/uin[1]
+ blk.column\[7\].row\[5\].yc/din[0] blk.column\[7\].row\[5\].yc/din[1] blk.column\[7\].row\[5\].yc/dempty
+ blk.column\[7\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_531_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_329_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_370_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_485_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_379_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_537_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_288_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_490_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_505_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_393_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_276_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_370_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_497_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_457_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_625_ VGND VGND VPWR VPWR _625_/HI io_oeb[37] sky130_fd_sc_hd__conb_1
XPHY_6296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_343_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_556_ VGND VGND VPWR VPWR _556_/HI _556_/LO sky130_fd_sc_hd__conb_1
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_487_ VGND VGND VPWR VPWR _487_/HI _487_/LO sky130_fd_sc_hd__conb_1
XFILLER_496_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_227_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_522_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_410_ wb_rst_i VGND VGND VPWR VPWR _410_/X sky130_fd_sc_hd__buf_2
XPHY_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_341_ _337_/Y _340_/X wbs_dat_i[23] _340_/X VGND VGND VPWR VPWR _791_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_319_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_534_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[10\].yc blk.column\[9\].row\[9\].yc/cbitout blk.column\[9\].row\[11\].yc/cbitin
+ blk.column\[9\].row\[9\].yc/confclko blk.column\[9\].row\[11\].yc/confclk blk.column\[9\].row\[10\].yc/dempty
+ blk.column\[9\].row\[10\].yc/din[0] blk.column\[9\].row\[10\].yc/din[1] blk.column\[9\].row\[11\].yc/uin[0]
+ blk.column\[9\].row\[11\].yc/uin[1] blk.column\[9\].row\[10\].yc/hempty blk.column\[8\].row\[10\].yc/lempty
+ blk.column\[9\].row\[10\].yc/lempty blk.column\[9\].row\[10\].yc/lin[0] blk.column\[9\].row\[10\].yc/lin[1]
+ blk.column\[9\].row\[10\].yc/lout[0] blk.column\[9\].row\[10\].yc/lout[1] blk.column\[8\].row\[10\].yc/hempty
+ blk.column\[9\].row\[9\].yc/reseto blk.column\[9\].row\[11\].yc/reset blk.column\[9\].row\[10\].yc/rin[0]
+ blk.column\[9\].row\[10\].yc/rin[1] blk.column\[8\].row\[10\].yc/lin[0] blk.column\[8\].row\[10\].yc/lin[1]
+ blk.column\[9\].row\[9\].yc/vempty2 blk.column\[9\].row\[9\].yc/dout[0] blk.column\[9\].row\[9\].yc/dout[1]
+ blk.column\[9\].row\[9\].yc/din[0] blk.column\[9\].row\[9\].yc/din[1] blk.column\[9\].row\[9\].yc/dempty
+ blk.column\[9\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_519_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_457_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_504_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_608_ VGND VGND VPWR VPWR _608_/HI io_oeb[20] sky130_fd_sc_hd__conb_1
XFILLER_441_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_539_ VGND VGND VPWR VPWR _539_/HI _539_/LO sky130_fd_sc_hd__conb_1
XFILLER_378_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_302_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_528_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_540_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_369_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_377_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_500_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_314_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_321_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ _319_/A VGND VGND VPWR VPWR _324_/X sky130_fd_sc_hd__buf_2
XFILLER_15_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[8\].row\[8\].yc blk.column\[8\].row\[8\].yc/cbitin blk.column\[8\].row\[9\].yc/cbitin
+ blk.column\[8\].row\[8\].yc/confclk blk.column\[8\].row\[9\].yc/confclk blk.column\[8\].row\[8\].yc/dempty
+ blk.column\[8\].row\[8\].yc/din[0] blk.column\[8\].row\[8\].yc/din[1] blk.column\[8\].row\[9\].yc/uin[0]
+ blk.column\[8\].row\[9\].yc/uin[1] blk.column\[8\].row\[8\].yc/hempty blk.column\[7\].row\[8\].yc/lempty
+ blk.column\[8\].row\[8\].yc/lempty blk.column\[8\].row\[8\].yc/lin[0] blk.column\[8\].row\[8\].yc/lin[1]
+ blk.column\[9\].row\[8\].yc/rin[0] blk.column\[9\].row\[8\].yc/rin[1] blk.column\[7\].row\[8\].yc/hempty
+ blk.column\[8\].row\[8\].yc/reset blk.column\[8\].row\[9\].yc/reset blk.column\[8\].row\[8\].yc/rin[0]
+ blk.column\[8\].row\[8\].yc/rin[1] blk.column\[7\].row\[8\].yc/lin[0] blk.column\[7\].row\[8\].yc/lin[1]
+ blk.column\[8\].row\[8\].yc/uempty blk.column\[8\].row\[8\].yc/uin[0] blk.column\[8\].row\[8\].yc/uin[1]
+ blk.column\[8\].row\[7\].yc/din[0] blk.column\[8\].row\[7\].yc/din[1] blk.column\[8\].row\[7\].yc/dempty
+ blk.column\[8\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_477_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_316_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_346_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_398_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_529_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_296_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_520_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_309_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_498_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_244_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_297_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_528_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_390_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_507_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_3039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_507_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_395_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_379_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_536_2109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_307_ _307_/A VGND VGND VPWR VPWR _307_/Y sky130_fd_sc_hd__inv_2
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_536_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_531_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[0\].yc la_data_in[108] blk.column\[12\].row\[1\].yc/cbitin
+ la_data_in[112] blk.column\[12\].row\[1\].yc/confclk blk.column\[12\].row\[0\].yc/dempty
+ blk.column\[12\].row\[0\].yc/din[0] blk.column\[12\].row\[0\].yc/din[1] blk.column\[12\].row\[1\].yc/uin[0]
+ blk.column\[12\].row\[1\].yc/uin[1] blk.column\[12\].row\[0\].yc/hempty blk.column\[11\].row\[0\].yc/lempty
+ blk.column\[12\].row\[0\].yc/lempty blk.column\[12\].row\[0\].yc/lin[0] blk.column\[12\].row\[0\].yc/lin[1]
+ blk.column\[13\].row\[0\].yc/rin[0] blk.column\[13\].row\[0\].yc/rin[1] blk.column\[11\].row\[0\].yc/hempty
+ la_data_in[113] blk.column\[12\].row\[1\].yc/reset blk.column\[12\].row\[0\].yc/rin[0]
+ blk.column\[12\].row\[0\].yc/rin[1] blk.column\[11\].row\[0\].yc/lin[0] blk.column\[11\].row\[0\].yc/lin[1]
+ _517_/LO la_data_in[88] la_data_in[89] la_data_out[24] la_data_out[25] blk.column\[12\].row\[0\].yc/vempty
+ blk.column\[12\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_178_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_339_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_493_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_335_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[1\].yc blk.column\[3\].row\[1\].yc/cbitin blk.column\[3\].row\[2\].yc/cbitin
+ blk.column\[3\].row\[1\].yc/confclk blk.column\[3\].row\[2\].yc/confclk blk.column\[3\].row\[1\].yc/dempty
+ blk.column\[3\].row\[1\].yc/din[0] blk.column\[3\].row\[1\].yc/din[1] blk.column\[3\].row\[2\].yc/uin[0]
+ blk.column\[3\].row\[2\].yc/uin[1] blk.column\[3\].row\[1\].yc/hempty blk.column\[2\].row\[1\].yc/lempty
+ blk.column\[3\].row\[1\].yc/lempty blk.column\[3\].row\[1\].yc/lin[0] blk.column\[3\].row\[1\].yc/lin[1]
+ blk.column\[4\].row\[1\].yc/rin[0] blk.column\[4\].row\[1\].yc/rin[1] blk.column\[2\].row\[1\].yc/hempty
+ blk.column\[3\].row\[1\].yc/reset blk.column\[3\].row\[2\].yc/reset blk.column\[3\].row\[1\].yc/rin[0]
+ blk.column\[3\].row\[1\].yc/rin[1] blk.column\[2\].row\[1\].yc/lin[0] blk.column\[2\].row\[1\].yc/lin[1]
+ blk.column\[3\].row\[1\].yc/uempty blk.column\[3\].row\[1\].yc/uin[0] blk.column\[3\].row\[1\].yc/uin[1]
+ blk.column\[3\].row\[0\].yc/din[0] blk.column\[3\].row\[0\].yc/din[1] blk.column\[3\].row\[0\].yc/dempty
+ blk.column\[3\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_510_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_322_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_420_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_298_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_458_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_472_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_531_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_526_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_787_ wb_clk_i _787_/D VGND VGND VPWR VPWR _349_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_1_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_514_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_345_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_421_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_538_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_497_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_513_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_710_ VGND VGND VPWR VPWR _710_/HI la_data_out[94] sky130_fd_sc_hd__conb_1
XPHY_6423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_641_ VGND VGND VPWR VPWR _641_/HI io_out[15] sky130_fd_sc_hd__conb_1
XPHY_6456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_572_ VGND VGND VPWR VPWR _572_/HI _572_/LO sky130_fd_sc_hd__conb_1
XPHY_5766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_353_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[11\].yc blk.column\[4\].row\[11\].yc/cbitin blk.column\[4\].row\[12\].yc/cbitin
+ blk.column\[4\].row\[11\].yc/confclk blk.column\[4\].row\[12\].yc/confclk blk.column\[4\].row\[11\].yc/dempty
+ blk.column\[4\].row\[11\].yc/din[0] blk.column\[4\].row\[11\].yc/din[1] blk.column\[4\].row\[12\].yc/uin[0]
+ blk.column\[4\].row\[12\].yc/uin[1] blk.column\[4\].row\[11\].yc/hempty blk.column\[3\].row\[11\].yc/lempty
+ blk.column\[4\].row\[11\].yc/lempty blk.column\[4\].row\[11\].yc/lin[0] blk.column\[4\].row\[11\].yc/lin[1]
+ blk.column\[5\].row\[11\].yc/rin[0] blk.column\[5\].row\[11\].yc/rin[1] blk.column\[3\].row\[11\].yc/hempty
+ blk.column\[4\].row\[11\].yc/reset blk.column\[4\].row\[12\].yc/reset blk.column\[4\].row\[11\].yc/rin[0]
+ blk.column\[4\].row\[11\].yc/rin[1] blk.column\[3\].row\[11\].yc/lin[0] blk.column\[3\].row\[11\].yc/lin[1]
+ blk.column\[4\].row\[11\].yc/uempty blk.column\[4\].row\[11\].yc/uin[0] blk.column\[4\].row\[11\].yc/uin[1]
+ blk.column\[4\].row\[10\].yc/din[0] blk.column\[4\].row\[10\].yc/din[1] blk.column\[4\].row\[10\].yc/dempty
+ blk.column\[4\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_16_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_396_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_490_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_513_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_475_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_538_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_511_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_282_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_402_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_510_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_512_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_624_ VGND VGND VPWR VPWR _624_/HI io_oeb[36] sky130_fd_sc_hd__conb_1
XPHY_6297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_382_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_343_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_555_ VGND VGND VPWR VPWR _555_/HI _555_/LO sky130_fd_sc_hd__conb_1
XFILLER_144_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_486_ VGND VGND VPWR VPWR _486_/HI _486_/LO sky130_fd_sc_hd__conb_1
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_536_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_533_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[2\].yc blk.column\[13\].row\[2\].yc/cbitin blk.column\[13\].row\[3\].yc/cbitin
+ blk.column\[13\].row\[2\].yc/confclk blk.column\[13\].row\[3\].yc/confclk blk.column\[13\].row\[2\].yc/dempty
+ blk.column\[13\].row\[2\].yc/din[0] blk.column\[13\].row\[2\].yc/din[1] blk.column\[13\].row\[3\].yc/uin[0]
+ blk.column\[13\].row\[3\].yc/uin[1] blk.column\[13\].row\[2\].yc/hempty blk.column\[12\].row\[2\].yc/lempty
+ blk.column\[13\].row\[2\].yc/lempty blk.column\[13\].row\[2\].yc/lin[0] blk.column\[13\].row\[2\].yc/lin[1]
+ blk.column\[14\].row\[2\].yc/rin[0] blk.column\[14\].row\[2\].yc/rin[1] blk.column\[12\].row\[2\].yc/hempty
+ blk.column\[13\].row\[2\].yc/reset blk.column\[13\].row\[3\].yc/reset blk.column\[13\].row\[2\].yc/rin[0]
+ blk.column\[13\].row\[2\].yc/rin[1] blk.column\[12\].row\[2\].yc/lin[0] blk.column\[12\].row\[2\].yc/lin[1]
+ blk.column\[13\].row\[2\].yc/uempty blk.column\[13\].row\[2\].yc/uin[0] blk.column\[13\].row\[2\].yc/uin[1]
+ blk.column\[13\].row\[1\].yc/din[0] blk.column\[13\].row\[1\].yc/din[1] blk.column\[13\].row\[1\].yc/dempty
+ blk.column\[13\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_416_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_541_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[3\].yc blk.column\[4\].row\[3\].yc/cbitin blk.column\[4\].row\[4\].yc/cbitin
+ blk.column\[4\].row\[3\].yc/confclk blk.column\[4\].row\[4\].yc/confclk blk.column\[4\].row\[3\].yc/dempty
+ blk.column\[4\].row\[3\].yc/din[0] blk.column\[4\].row\[3\].yc/din[1] blk.column\[4\].row\[4\].yc/uin[0]
+ blk.column\[4\].row\[4\].yc/uin[1] blk.column\[4\].row\[3\].yc/hempty blk.column\[3\].row\[3\].yc/lempty
+ blk.column\[4\].row\[3\].yc/lempty blk.column\[4\].row\[3\].yc/lin[0] blk.column\[4\].row\[3\].yc/lin[1]
+ blk.column\[5\].row\[3\].yc/rin[0] blk.column\[5\].row\[3\].yc/rin[1] blk.column\[3\].row\[3\].yc/hempty
+ blk.column\[4\].row\[3\].yc/reset blk.column\[4\].row\[4\].yc/reset blk.column\[4\].row\[3\].yc/rin[0]
+ blk.column\[4\].row\[3\].yc/rin[1] blk.column\[3\].row\[3\].yc/lin[0] blk.column\[3\].row\[3\].yc/lin[1]
+ blk.column\[4\].row\[3\].yc/uempty blk.column\[4\].row\[3\].yc/uin[0] blk.column\[4\].row\[3\].yc/uin[1]
+ blk.column\[4\].row\[2\].yc/din[0] blk.column\[4\].row\[2\].yc/din[1] blk.column\[4\].row\[2\].yc/dempty
+ blk.column\[4\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_527_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xblk.column\[11\].row\[13\].yc blk.column\[11\].row\[13\].yc/cbitin blk.column\[11\].row\[14\].yc/cbitin
+ blk.column\[11\].row\[13\].yc/confclk blk.column\[11\].row\[14\].yc/confclk blk.column\[11\].row\[13\].yc/dempty
+ blk.column\[11\].row\[13\].yc/din[0] blk.column\[11\].row\[13\].yc/din[1] blk.column\[11\].row\[14\].yc/uin[0]
+ blk.column\[11\].row\[14\].yc/uin[1] blk.column\[11\].row\[13\].yc/hempty blk.column\[10\].row\[13\].yc/lempty
+ blk.column\[11\].row\[13\].yc/lempty blk.column\[11\].row\[13\].yc/lin[0] blk.column\[11\].row\[13\].yc/lin[1]
+ blk.column\[12\].row\[13\].yc/rin[0] blk.column\[12\].row\[13\].yc/rin[1] blk.column\[10\].row\[13\].yc/hempty
+ blk.column\[11\].row\[13\].yc/reset blk.column\[11\].row\[14\].yc/reset blk.column\[11\].row\[13\].yc/rin[0]
+ blk.column\[11\].row\[13\].yc/rin[1] blk.column\[10\].row\[13\].yc/lin[0] blk.column\[10\].row\[13\].yc/lin[1]
+ blk.column\[11\].row\[13\].yc/uempty blk.column\[11\].row\[13\].yc/uin[0] blk.column\[11\].row\[13\].yc/uin[1]
+ blk.column\[11\].row\[12\].yc/din[0] blk.column\[11\].row\[12\].yc/din[1] blk.column\[11\].row\[12\].yc/dempty
+ blk.column\[11\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_514_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_527_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_340_ _339_/X VGND VGND VPWR VPWR _340_/X sky130_fd_sc_hd__buf_2
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_430_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_319_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_516_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_491_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_457_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_326_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_607_ VGND VGND VPWR VPWR _607_/HI io_oeb[19] sky130_fd_sc_hd__conb_1
XPHY_5382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_476_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_538_ VGND VGND VPWR VPWR _538_/HI _538_/LO sky130_fd_sc_hd__conb_1
XPHY_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_469_ VGND VGND VPWR VPWR _469_/HI _469_/LO sky130_fd_sc_hd__conb_1
XFILLER_259_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_278_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_524_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_530_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_389_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_383_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_266_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_320_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_457_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_539_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_492_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_238_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[14\].yc blk.column\[8\].row\[14\].yc/cbitin blk.column\[8\].row\[15\].yc/cbitin
+ blk.column\[8\].row\[14\].yc/confclk blk.column\[8\].row\[15\].yc/confclk blk.column\[8\].row\[14\].yc/dempty
+ blk.column\[8\].row\[14\].yc/din[0] blk.column\[8\].row\[14\].yc/din[1] blk.column\[8\].row\[15\].yc/uin[0]
+ blk.column\[8\].row\[15\].yc/uin[1] blk.column\[8\].row\[14\].yc/hempty blk.column\[7\].row\[14\].yc/lempty
+ blk.column\[8\].row\[14\].yc/lempty blk.column\[8\].row\[14\].yc/lin[0] blk.column\[8\].row\[14\].yc/lin[1]
+ blk.column\[9\].row\[14\].yc/rin[0] blk.column\[9\].row\[14\].yc/rin[1] blk.column\[7\].row\[14\].yc/hempty
+ blk.column\[8\].row\[14\].yc/reset blk.column\[8\].row\[15\].yc/reset blk.column\[8\].row\[14\].yc/rin[0]
+ blk.column\[8\].row\[14\].yc/rin[1] blk.column\[7\].row\[14\].yc/lin[0] blk.column\[7\].row\[14\].yc/lin[1]
+ blk.column\[8\].row\[14\].yc/uempty blk.column\[8\].row\[14\].yc/uin[0] blk.column\[8\].row\[14\].yc/uin[1]
+ blk.column\[8\].row\[13\].yc/din[0] blk.column\[8\].row\[13\].yc/din[1] blk.column\[8\].row\[13\].yc/dempty
+ blk.column\[8\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_191_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_533_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_413_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_323_ _323_/A VGND VGND VPWR VPWR _323_/Y sky130_fd_sc_hd__inv_2
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_375_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_534_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_322_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_297_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_400_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_528_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_542_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_520_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_519_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_306_ _305_/Y _303_/X wbs_dat_i[4] _303_/X VGND VGND VPWR VPWR _306_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_493_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_533_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_236_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[4\].yc blk.column\[14\].row\[4\].yc/cbitin blk.column\[14\].row\[5\].yc/cbitin
+ blk.column\[14\].row\[4\].yc/confclk blk.column\[14\].row\[5\].yc/confclk blk.column\[14\].row\[4\].yc/dempty
+ blk.column\[14\].row\[4\].yc/din[0] blk.column\[14\].row\[4\].yc/din[1] blk.column\[14\].row\[5\].yc/uin[0]
+ blk.column\[14\].row\[5\].yc/uin[1] blk.column\[14\].row\[4\].yc/hempty blk.column\[13\].row\[4\].yc/lempty
+ blk.column\[14\].row\[4\].yc/lempty blk.column\[14\].row\[4\].yc/lin[0] blk.column\[14\].row\[4\].yc/lin[1]
+ blk.column\[15\].row\[4\].yc/rin[0] blk.column\[15\].row\[4\].yc/rin[1] blk.column\[13\].row\[4\].yc/hempty
+ blk.column\[14\].row\[4\].yc/reset blk.column\[14\].row\[5\].yc/reset blk.column\[14\].row\[4\].yc/rin[0]
+ blk.column\[14\].row\[4\].yc/rin[1] blk.column\[13\].row\[4\].yc/lin[0] blk.column\[13\].row\[4\].yc/lin[1]
+ blk.column\[14\].row\[4\].yc/uempty blk.column\[14\].row\[4\].yc/uin[0] blk.column\[14\].row\[4\].yc/uin[1]
+ blk.column\[14\].row\[3\].yc/din[0] blk.column\[14\].row\[3\].yc/din[1] blk.column\[14\].row\[3\].yc/dempty
+ blk.column\[14\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_530_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_512_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_458_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_386_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_466_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_473_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_304_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[5\].yc blk.column\[5\].row\[5\].yc/cbitin blk.column\[5\].row\[6\].yc/cbitin
+ blk.column\[5\].row\[5\].yc/confclk blk.column\[5\].row\[6\].yc/confclk blk.column\[5\].row\[5\].yc/dempty
+ blk.column\[5\].row\[5\].yc/din[0] blk.column\[5\].row\[5\].yc/din[1] blk.column\[5\].row\[6\].yc/uin[0]
+ blk.column\[5\].row\[6\].yc/uin[1] blk.column\[5\].row\[5\].yc/hempty blk.column\[4\].row\[5\].yc/lempty
+ blk.column\[5\].row\[5\].yc/lempty blk.column\[5\].row\[5\].yc/lin[0] blk.column\[5\].row\[5\].yc/lin[1]
+ blk.column\[6\].row\[5\].yc/rin[0] blk.column\[6\].row\[5\].yc/rin[1] blk.column\[4\].row\[5\].yc/hempty
+ blk.column\[5\].row\[5\].yc/reset blk.column\[5\].row\[6\].yc/reset blk.column\[5\].row\[5\].yc/rin[0]
+ blk.column\[5\].row\[5\].yc/rin[1] blk.column\[4\].row\[5\].yc/lin[0] blk.column\[4\].row\[5\].yc/lin[1]
+ blk.column\[5\].row\[5\].yc/uempty blk.column\[5\].row\[5\].yc/uin[0] blk.column\[5\].row\[5\].yc/uin[1]
+ blk.column\[5\].row\[4\].yc/din[0] blk.column\[5\].row\[4\].yc/din[1] blk.column\[5\].row\[4\].yc/dempty
+ blk.column\[5\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_225_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_499_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_536_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_497_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_350_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_311_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_417_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_420_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_279_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_474_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_515_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_531_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_507_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_786_ wb_clk_i _786_/D VGND VGND VPWR VPWR _786_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_423_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_336_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_536_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_317_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_392_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_488_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_380_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_495_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_508_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_444_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_640_ VGND VGND VPWR VPWR _640_/HI io_out[14] sky130_fd_sc_hd__conb_1
XFILLER_492_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_571_ VGND VGND VPWR VPWR _571_/HI _571_/LO sky130_fd_sc_hd__conb_1
XFILLER_404_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_474_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_469_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_487_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_507_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_769_ wb_clk_i _769_/D VGND VGND VPWR VPWR wbs_dat_o[25] sky130_fd_sc_hd__dfxtp_4
XFILLER_250_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_451_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_522_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_434_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[15\].yc blk.column\[3\].row\[15\].yc/cbitin la_data_out[35]
+ blk.column\[3\].row\[15\].yc/confclk blk.column\[3\].row\[15\].yc/confclko _469_/HI
+ _568_/LO _569_/LO blk.column\[3\].row\[15\].yc/dout[0] blk.column\[3\].row\[15\].yc/dout[1]
+ blk.column\[3\].row\[15\].yc/hempty blk.column\[2\].row\[15\].yc/lempty blk.column\[3\].row\[15\].yc/lempty
+ blk.column\[3\].row\[15\].yc/lin[0] blk.column\[3\].row\[15\].yc/lin[1] blk.column\[4\].row\[15\].yc/rin[0]
+ blk.column\[4\].row\[15\].yc/rin[1] blk.column\[2\].row\[15\].yc/hempty blk.column\[3\].row\[15\].yc/reset
+ blk.column\[3\].row\[15\].yc/reseto blk.column\[3\].row\[15\].yc/rin[0] blk.column\[3\].row\[15\].yc/rin[1]
+ blk.column\[2\].row\[15\].yc/lin[0] blk.column\[2\].row\[15\].yc/lin[1] blk.column\[3\].row\[15\].yc/uempty
+ blk.column\[3\].row\[15\].yc/uin[0] blk.column\[3\].row\[15\].yc/uin[1] blk.column\[3\].row\[14\].yc/din[0]
+ blk.column\[3\].row\[14\].yc/din[1] blk.column\[3\].row\[14\].yc/dempty blk.column\[3\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_510_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_10913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_623_ VGND VGND VPWR VPWR _623_/HI io_oeb[35] sky130_fd_sc_hd__conb_1
XPHY_6276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_382_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_554_ VGND VGND VPWR VPWR _554_/HI _554_/LO sky130_fd_sc_hd__conb_1
XPHY_5597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_485_ VGND VGND VPWR VPWR _485_/HI _485_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_496_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[6\].yc blk.column\[15\].row\[6\].yc/cbitin blk.column\[15\].row\[7\].yc/cbitin
+ blk.column\[15\].row\[6\].yc/confclk blk.column\[15\].row\[7\].yc/confclk blk.column\[15\].row\[6\].yc/dempty
+ blk.column\[15\].row\[6\].yc/din[0] blk.column\[15\].row\[6\].yc/din[1] blk.column\[15\].row\[7\].yc/uin[0]
+ blk.column\[15\].row\[7\].yc/uin[1] blk.column\[15\].row\[6\].yc/hempty blk.column\[14\].row\[6\].yc/lempty
+ _463_/HI _553_/LO _554_/LO blk.column\[15\].row\[6\].yc/lout[0] blk.column\[15\].row\[6\].yc/lout[1]
+ blk.column\[14\].row\[6\].yc/hempty blk.column\[15\].row\[6\].yc/reset blk.column\[15\].row\[7\].yc/reset
+ blk.column\[15\].row\[6\].yc/rin[0] blk.column\[15\].row\[6\].yc/rin[1] blk.column\[14\].row\[6\].yc/lin[0]
+ blk.column\[14\].row\[6\].yc/lin[1] blk.column\[15\].row\[6\].yc/uempty blk.column\[15\].row\[6\].yc/uin[0]
+ blk.column\[15\].row\[6\].yc/uin[1] blk.column\[15\].row\[5\].yc/din[0] blk.column\[15\].row\[5\].yc/din[1]
+ blk.column\[15\].row\[5\].yc/dempty blk.column\[15\].row\[7\].yc/uempty VPWR VGND
+ ycell
XFILLER_197_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_302_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[7\].yc blk.column\[6\].row\[7\].yc/cbitin blk.column\[6\].row\[8\].yc/cbitin
+ blk.column\[6\].row\[7\].yc/confclk blk.column\[6\].row\[8\].yc/confclk blk.column\[6\].row\[7\].yc/dempty
+ blk.column\[6\].row\[7\].yc/din[0] blk.column\[6\].row\[7\].yc/din[1] blk.column\[6\].row\[8\].yc/uin[0]
+ blk.column\[6\].row\[8\].yc/uin[1] blk.column\[6\].row\[7\].yc/hempty blk.column\[5\].row\[7\].yc/lempty
+ blk.column\[6\].row\[7\].yc/lempty blk.column\[6\].row\[7\].yc/lin[0] blk.column\[6\].row\[7\].yc/lin[1]
+ blk.column\[7\].row\[7\].yc/rin[0] blk.column\[7\].row\[7\].yc/rin[1] blk.column\[5\].row\[7\].yc/hempty
+ blk.column\[6\].row\[7\].yc/reset blk.column\[6\].row\[8\].yc/reset blk.column\[6\].row\[7\].yc/rin[0]
+ blk.column\[6\].row\[7\].yc/rin[1] blk.column\[5\].row\[7\].yc/lin[0] blk.column\[5\].row\[7\].yc/lin[1]
+ blk.column\[6\].row\[7\].yc/uempty blk.column\[6\].row\[7\].yc/uin[0] blk.column\[6\].row\[7\].yc/uin[1]
+ blk.column\[6\].row\[6\].yc/din[0] blk.column\[6\].row\[6\].yc/din[1] blk.column\[6\].row\[6\].yc/dempty
+ blk.column\[6\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_500_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_503_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_492_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_466_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_447_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_430_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_516_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_413_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_606_ VGND VGND VPWR VPWR _606_/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XPHY_5361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_232_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_537_ VGND VGND VPWR VPWR _537_/HI _537_/LO sky130_fd_sc_hd__conb_1
XPHY_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_501_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_468_ VGND VGND VPWR VPWR _468_/HI _468_/LO sky130_fd_sc_hd__conb_1
XFILLER_14_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_399_ _398_/X wbs_dat_o[20] _347_/A _396_/X VGND VGND VPWR VPWR _764_/D sky130_fd_sc_hd__o22a_4
XFILLER_509_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_534_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_429_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_215_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_326_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_498_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_457_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_413_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[0\].yc la_data_in[97] blk.column\[1\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[1\].row\[1\].yc/confclk blk.column\[1\].row\[0\].yc/dempty blk.column\[1\].row\[0\].yc/din[0]
+ blk.column\[1\].row\[0\].yc/din[1] blk.column\[1\].row\[1\].yc/uin[0] blk.column\[1\].row\[1\].yc/uin[1]
+ blk.column\[1\].row\[0\].yc/hempty blk.column\[0\].row\[0\].yc/lempty blk.column\[1\].row\[0\].yc/lempty
+ blk.column\[1\].row\[0\].yc/lin[0] blk.column\[1\].row\[0\].yc/lin[1] blk.column\[2\].row\[0\].yc/rin[0]
+ blk.column\[2\].row\[0\].yc/rin[1] blk.column\[0\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[1\].row\[1\].yc/reset blk.column\[1\].row\[0\].yc/rin[0] blk.column\[1\].row\[0\].yc/rin[1]
+ blk.column\[0\].row\[0\].yc/lin[0] blk.column\[0\].row\[0\].yc/lin[1] _561_/LO la_data_in[66]
+ la_data_in[67] la_data_out[2] la_data_out[3] blk.column\[1\].row\[0\].yc/vempty
+ blk.column\[1\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_497_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_322_ _321_/Y _319_/X wbs_dat_i[14] _319_/X VGND VGND VPWR VPWR _798_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[10\].yc blk.column\[5\].row\[9\].yc/cbitout blk.column\[5\].row\[11\].yc/cbitin
+ blk.column\[5\].row\[9\].yc/confclko blk.column\[5\].row\[11\].yc/confclk blk.column\[5\].row\[10\].yc/dempty
+ blk.column\[5\].row\[10\].yc/din[0] blk.column\[5\].row\[10\].yc/din[1] blk.column\[5\].row\[11\].yc/uin[0]
+ blk.column\[5\].row\[11\].yc/uin[1] blk.column\[5\].row\[10\].yc/hempty blk.column\[4\].row\[10\].yc/lempty
+ blk.column\[5\].row\[10\].yc/lempty blk.column\[5\].row\[10\].yc/lin[0] blk.column\[5\].row\[10\].yc/lin[1]
+ blk.column\[6\].row\[10\].yc/rin[0] blk.column\[6\].row\[10\].yc/rin[1] blk.column\[4\].row\[10\].yc/hempty
+ blk.column\[5\].row\[9\].yc/reseto blk.column\[5\].row\[11\].yc/reset blk.column\[5\].row\[10\].yc/rin[0]
+ blk.column\[5\].row\[10\].yc/rin[1] blk.column\[4\].row\[10\].yc/lin[0] blk.column\[4\].row\[10\].yc/lin[1]
+ blk.column\[5\].row\[9\].yc/vempty2 blk.column\[5\].row\[9\].yc/dout[0] blk.column\[5\].row\[9\].yc/dout[1]
+ blk.column\[5\].row\[9\].yc/din[0] blk.column\[5\].row\[9\].yc/din[1] blk.column\[5\].row\[9\].yc/dempty
+ blk.column\[5\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_453_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_356_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_532_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_476_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_528_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_481_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_498_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_300_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_355_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_527_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_483_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_507_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_2675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_2307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_540_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_505_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_520_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_305_ _305_/A VGND VGND VPWR VPWR _305_/Y sky130_fd_sc_hd__inv_2
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_256_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[9\].yc blk.column\[7\].row\[9\].yc/cbitin blk.column\[7\].row\[9\].yc/cbitout
+ blk.column\[7\].row\[9\].yc/confclk blk.column\[7\].row\[9\].yc/confclko blk.column\[7\].row\[9\].yc/dempty
+ blk.column\[7\].row\[9\].yc/din[0] blk.column\[7\].row\[9\].yc/din[1] blk.column\[7\].row\[9\].yc/dout[0]
+ blk.column\[7\].row\[9\].yc/dout[1] blk.column\[7\].row\[9\].yc/hempty blk.column\[6\].row\[9\].yc/lempty
+ blk.column\[7\].row\[9\].yc/lempty blk.column\[7\].row\[9\].yc/lin[0] blk.column\[7\].row\[9\].yc/lin[1]
+ blk.column\[8\].row\[9\].yc/rin[0] blk.column\[8\].row\[9\].yc/rin[1] blk.column\[6\].row\[9\].yc/hempty
+ blk.column\[7\].row\[9\].yc/reset blk.column\[7\].row\[9\].yc/reseto blk.column\[7\].row\[9\].yc/rin[0]
+ blk.column\[7\].row\[9\].yc/rin[1] blk.column\[6\].row\[9\].yc/lin[0] blk.column\[6\].row\[9\].yc/lin[1]
+ blk.column\[7\].row\[9\].yc/uempty blk.column\[7\].row\[9\].yc/uin[0] blk.column\[7\].row\[9\].yc/uin[1]
+ blk.column\[7\].row\[8\].yc/din[0] blk.column\[7\].row\[8\].yc/din[1] blk.column\[7\].row\[8\].yc/dempty
+ blk.column\[7\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_507_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_312_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_458_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_473_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_394_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_410_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_528_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_437_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_458_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[12\].yc blk.column\[12\].row\[12\].yc/cbitin blk.column\[12\].row\[13\].yc/cbitin
+ blk.column\[12\].row\[12\].yc/confclk blk.column\[12\].row\[13\].yc/confclk blk.column\[12\].row\[12\].yc/dempty
+ blk.column\[12\].row\[12\].yc/din[0] blk.column\[12\].row\[12\].yc/din[1] blk.column\[12\].row\[13\].yc/uin[0]
+ blk.column\[12\].row\[13\].yc/uin[1] blk.column\[12\].row\[12\].yc/hempty blk.column\[11\].row\[12\].yc/lempty
+ blk.column\[12\].row\[12\].yc/lempty blk.column\[12\].row\[12\].yc/lin[0] blk.column\[12\].row\[12\].yc/lin[1]
+ blk.column\[13\].row\[12\].yc/rin[0] blk.column\[13\].row\[12\].yc/rin[1] blk.column\[11\].row\[12\].yc/hempty
+ blk.column\[12\].row\[12\].yc/reset blk.column\[12\].row\[13\].yc/reset blk.column\[12\].row\[12\].yc/rin[0]
+ blk.column\[12\].row\[12\].yc/rin[1] blk.column\[11\].row\[12\].yc/lin[0] blk.column\[11\].row\[12\].yc/lin[1]
+ blk.column\[12\].row\[12\].yc/uempty blk.column\[12\].row\[12\].yc/uin[0] blk.column\[12\].row\[12\].yc/uin[1]
+ blk.column\[12\].row\[11\].yc/din[0] blk.column\[12\].row\[11\].yc/din[1] blk.column\[12\].row\[11\].yc/dempty
+ blk.column\[12\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_535_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_487_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_343_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_785_ wb_clk_i _355_/X VGND VGND VPWR VPWR _354_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_131_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_373_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_384_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_488_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_300_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_384_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_503_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_278_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_495_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[1\].yc blk.column\[11\].row\[1\].yc/cbitin blk.column\[11\].row\[2\].yc/cbitin
+ blk.column\[11\].row\[1\].yc/confclk blk.column\[11\].row\[2\].yc/confclk blk.column\[11\].row\[1\].yc/dempty
+ blk.column\[11\].row\[1\].yc/din[0] blk.column\[11\].row\[1\].yc/din[1] blk.column\[11\].row\[2\].yc/uin[0]
+ blk.column\[11\].row\[2\].yc/uin[1] blk.column\[11\].row\[1\].yc/hempty blk.column\[10\].row\[1\].yc/lempty
+ blk.column\[11\].row\[1\].yc/lempty blk.column\[11\].row\[1\].yc/lin[0] blk.column\[11\].row\[1\].yc/lin[1]
+ blk.column\[12\].row\[1\].yc/rin[0] blk.column\[12\].row\[1\].yc/rin[1] blk.column\[10\].row\[1\].yc/hempty
+ blk.column\[11\].row\[1\].yc/reset blk.column\[11\].row\[2\].yc/reset blk.column\[11\].row\[1\].yc/rin[0]
+ blk.column\[11\].row\[1\].yc/rin[1] blk.column\[10\].row\[1\].yc/lin[0] blk.column\[10\].row\[1\].yc/lin[1]
+ blk.column\[11\].row\[1\].yc/uempty blk.column\[11\].row\[1\].yc/uin[0] blk.column\[11\].row\[1\].yc/uin[1]
+ blk.column\[11\].row\[0\].yc/din[0] blk.column\[11\].row\[0\].yc/din[1] blk.column\[11\].row\[0\].yc/dempty
+ blk.column\[11\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_519_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_524_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[2\].row\[2\].yc blk.column\[2\].row\[2\].yc/cbitin blk.column\[2\].row\[3\].yc/cbitin
+ blk.column\[2\].row\[2\].yc/confclk blk.column\[2\].row\[3\].yc/confclk blk.column\[2\].row\[2\].yc/dempty
+ blk.column\[2\].row\[2\].yc/din[0] blk.column\[2\].row\[2\].yc/din[1] blk.column\[2\].row\[3\].yc/uin[0]
+ blk.column\[2\].row\[3\].yc/uin[1] blk.column\[2\].row\[2\].yc/hempty blk.column\[1\].row\[2\].yc/lempty
+ blk.column\[2\].row\[2\].yc/lempty blk.column\[2\].row\[2\].yc/lin[0] blk.column\[2\].row\[2\].yc/lin[1]
+ blk.column\[3\].row\[2\].yc/rin[0] blk.column\[3\].row\[2\].yc/rin[1] blk.column\[1\].row\[2\].yc/hempty
+ blk.column\[2\].row\[2\].yc/reset blk.column\[2\].row\[3\].yc/reset blk.column\[2\].row\[2\].yc/rin[0]
+ blk.column\[2\].row\[2\].yc/rin[1] blk.column\[1\].row\[2\].yc/lin[0] blk.column\[1\].row\[2\].yc/lin[1]
+ blk.column\[2\].row\[2\].yc/uempty blk.column\[2\].row\[2\].yc/uin[0] blk.column\[2\].row\[2\].yc/uin[1]
+ blk.column\[2\].row\[1\].yc/din[0] blk.column\[2\].row\[1\].yc/din[1] blk.column\[2\].row\[1\].yc/dempty
+ blk.column\[2\].row\[3\].yc/uempty VPWR VGND ycell
XPHY_6414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_570_ VGND VGND VPWR VPWR _570_/HI _570_/LO sky130_fd_sc_hd__conb_1
XFILLER_0_3070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_521_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_339_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[13\].yc blk.column\[9\].row\[13\].yc/cbitin blk.column\[9\].row\[14\].yc/cbitin
+ blk.column\[9\].row\[13\].yc/confclk blk.column\[9\].row\[14\].yc/confclk blk.column\[9\].row\[13\].yc/dempty
+ blk.column\[9\].row\[13\].yc/din[0] blk.column\[9\].row\[13\].yc/din[1] blk.column\[9\].row\[14\].yc/uin[0]
+ blk.column\[9\].row\[14\].yc/uin[1] blk.column\[9\].row\[13\].yc/hempty blk.column\[8\].row\[13\].yc/lempty
+ blk.column\[9\].row\[13\].yc/lempty blk.column\[9\].row\[13\].yc/lin[0] blk.column\[9\].row\[13\].yc/lin[1]
+ blk.column\[9\].row\[13\].yc/lout[0] blk.column\[9\].row\[13\].yc/lout[1] blk.column\[8\].row\[13\].yc/hempty
+ blk.column\[9\].row\[13\].yc/reset blk.column\[9\].row\[14\].yc/reset blk.column\[9\].row\[13\].yc/rin[0]
+ blk.column\[9\].row\[13\].yc/rin[1] blk.column\[8\].row\[13\].yc/lin[0] blk.column\[8\].row\[13\].yc/lin[1]
+ blk.column\[9\].row\[13\].yc/uempty blk.column\[9\].row\[13\].yc/uin[0] blk.column\[9\].row\[13\].yc/uin[1]
+ blk.column\[9\].row\[12\].yc/din[0] blk.column\[9\].row\[12\].yc/din[1] blk.column\[9\].row\[12\].yc/dempty
+ blk.column\[9\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_338_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_495_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_537_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_506_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_417_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_314_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_368_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_434_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_303_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_529_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_768_ wb_clk_i _768_/D VGND VGND VPWR VPWR wbs_dat_o[24] sky130_fd_sc_hd__dfxtp_4
XFILLER_235_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_699_ VGND VGND VPWR VPWR _699_/HI la_data_out[83] sky130_fd_sc_hd__conb_1
XFILLER_1_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_506_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_280_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_430_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_399_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_510_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_622_ VGND VGND VPWR VPWR _622_/HI io_oeb[34] sky130_fd_sc_hd__conb_1
XFILLER_484_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_526_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_382_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_553_ VGND VGND VPWR VPWR _553_/HI _553_/LO sky130_fd_sc_hd__conb_1
XPHY_5587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_484_ VGND VGND VPWR VPWR _484_/HI _484_/LO sky130_fd_sc_hd__conb_1
XPHY_4886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_420_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_537_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_531_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[11\].yc blk.column\[0\].row\[11\].yc/cbitin blk.column\[0\].row\[12\].yc/cbitin
+ blk.column\[0\].row\[11\].yc/confclk blk.column\[0\].row\[12\].yc/confclk blk.column\[0\].row\[11\].yc/dempty
+ blk.column\[0\].row\[11\].yc/din[0] blk.column\[0\].row\[11\].yc/din[1] blk.column\[0\].row\[12\].yc/uin[0]
+ blk.column\[0\].row\[12\].yc/uin[1] blk.column\[0\].row\[11\].yc/hempty blk.column\[0\].row\[11\].yc/hempty2
+ blk.column\[0\].row\[11\].yc/lempty blk.column\[0\].row\[11\].yc/lin[0] blk.column\[0\].row\[11\].yc/lin[1]
+ blk.column\[1\].row\[11\].yc/rin[0] blk.column\[1\].row\[11\].yc/rin[1] _430_/HI
+ blk.column\[0\].row\[11\].yc/reset blk.column\[0\].row\[12\].yc/reset _481_/LO _482_/LO
+ blk.column\[0\].row\[11\].yc/rout[0] blk.column\[0\].row\[11\].yc/rout[1] blk.column\[0\].row\[11\].yc/uempty
+ blk.column\[0\].row\[11\].yc/uin[0] blk.column\[0\].row\[11\].yc/uin[1] blk.column\[0\].row\[10\].yc/din[0]
+ blk.column\[0\].row\[10\].yc/din[1] blk.column\[0\].row\[10\].yc/dempty blk.column\[0\].row\[12\].yc/uempty
+ VPWR VGND ycell
XFILLER_302_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_531_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_416_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_381_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_503_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_457_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_447_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_527_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_480_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_401_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_351_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_406_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_605_ VGND VGND VPWR VPWR _605_/HI io_oeb[17] sky130_fd_sc_hd__conb_1
XPHY_5362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_536_ VGND VGND VPWR VPWR _536_/HI _536_/LO sky130_fd_sc_hd__conb_1
XPHY_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_467_ VGND VGND VPWR VPWR _467_/HI _467_/LO sky130_fd_sc_hd__conb_1
XPHY_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_535_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_398_ _419_/A VGND VGND VPWR VPWR _398_/X sky130_fd_sc_hd__buf_2
XFILLER_491_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[3\].yc blk.column\[12\].row\[3\].yc/cbitin blk.column\[12\].row\[4\].yc/cbitin
+ blk.column\[12\].row\[3\].yc/confclk blk.column\[12\].row\[4\].yc/confclk blk.column\[12\].row\[3\].yc/dempty
+ blk.column\[12\].row\[3\].yc/din[0] blk.column\[12\].row\[3\].yc/din[1] blk.column\[12\].row\[4\].yc/uin[0]
+ blk.column\[12\].row\[4\].yc/uin[1] blk.column\[12\].row\[3\].yc/hempty blk.column\[11\].row\[3\].yc/lempty
+ blk.column\[12\].row\[3\].yc/lempty blk.column\[12\].row\[3\].yc/lin[0] blk.column\[12\].row\[3\].yc/lin[1]
+ blk.column\[13\].row\[3\].yc/rin[0] blk.column\[13\].row\[3\].yc/rin[1] blk.column\[11\].row\[3\].yc/hempty
+ blk.column\[12\].row\[3\].yc/reset blk.column\[12\].row\[4\].yc/reset blk.column\[12\].row\[3\].yc/rin[0]
+ blk.column\[12\].row\[3\].yc/rin[1] blk.column\[11\].row\[3\].yc/lin[0] blk.column\[11\].row\[3\].yc/lin[1]
+ blk.column\[12\].row\[3\].yc/uempty blk.column\[12\].row\[3\].yc/uin[0] blk.column\[12\].row\[3\].yc/uin[1]
+ blk.column\[12\].row\[2\].yc/din[0] blk.column\[12\].row\[2\].yc/din[1] blk.column\[12\].row\[2\].yc/dempty
+ blk.column\[12\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_526_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_384_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_496_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[4\].yc blk.column\[3\].row\[4\].yc/cbitin blk.column\[3\].row\[5\].yc/cbitin
+ blk.column\[3\].row\[4\].yc/confclk blk.column\[3\].row\[5\].yc/confclk blk.column\[3\].row\[4\].yc/dempty
+ blk.column\[3\].row\[4\].yc/din[0] blk.column\[3\].row\[4\].yc/din[1] blk.column\[3\].row\[5\].yc/uin[0]
+ blk.column\[3\].row\[5\].yc/uin[1] blk.column\[3\].row\[4\].yc/hempty blk.column\[2\].row\[4\].yc/lempty
+ blk.column\[3\].row\[4\].yc/lempty blk.column\[3\].row\[4\].yc/lin[0] blk.column\[3\].row\[4\].yc/lin[1]
+ blk.column\[4\].row\[4\].yc/rin[0] blk.column\[4\].row\[4\].yc/rin[1] blk.column\[2\].row\[4\].yc/hempty
+ blk.column\[3\].row\[4\].yc/reset blk.column\[3\].row\[5\].yc/reset blk.column\[3\].row\[4\].yc/rin[0]
+ blk.column\[3\].row\[4\].yc/rin[1] blk.column\[2\].row\[4\].yc/lin[0] blk.column\[2\].row\[4\].yc/lin[1]
+ blk.column\[3\].row\[4\].yc/uempty blk.column\[3\].row\[4\].yc/uin[0] blk.column\[3\].row\[4\].yc/uin[1]
+ blk.column\[3\].row\[3\].yc/din[0] blk.column\[3\].row\[3\].yc/din[1] blk.column\[3\].row\[3\].yc/dempty
+ blk.column\[3\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_318_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_491_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_527_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_325_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_401_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_321_ _321_/A VGND VGND VPWR VPWR _321_/Y sky130_fd_sc_hd__inv_2
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_420_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_368_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_383_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_311_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_519_ VGND VGND VPWR VPWR _519_/HI _519_/LO sky130_fd_sc_hd__conb_1
XFILLER_366_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_2805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_256_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_528_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_221_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_459_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_251_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_300_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_365_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_510_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[14\].yc blk.column\[4\].row\[14\].yc/cbitin blk.column\[4\].row\[15\].yc/cbitin
+ blk.column\[4\].row\[14\].yc/confclk blk.column\[4\].row\[15\].yc/confclk blk.column\[4\].row\[14\].yc/dempty
+ blk.column\[4\].row\[14\].yc/din[0] blk.column\[4\].row\[14\].yc/din[1] blk.column\[4\].row\[15\].yc/uin[0]
+ blk.column\[4\].row\[15\].yc/uin[1] blk.column\[4\].row\[14\].yc/hempty blk.column\[3\].row\[14\].yc/lempty
+ blk.column\[4\].row\[14\].yc/lempty blk.column\[4\].row\[14\].yc/lin[0] blk.column\[4\].row\[14\].yc/lin[1]
+ blk.column\[5\].row\[14\].yc/rin[0] blk.column\[5\].row\[14\].yc/rin[1] blk.column\[3\].row\[14\].yc/hempty
+ blk.column\[4\].row\[14\].yc/reset blk.column\[4\].row\[15\].yc/reset blk.column\[4\].row\[14\].yc/rin[0]
+ blk.column\[4\].row\[14\].yc/rin[1] blk.column\[3\].row\[14\].yc/lin[0] blk.column\[3\].row\[14\].yc/lin[1]
+ blk.column\[4\].row\[14\].yc/uempty blk.column\[4\].row\[14\].yc/uin[0] blk.column\[4\].row\[14\].yc/uin[1]
+ blk.column\[4\].row\[13\].yc/din[0] blk.column\[4\].row\[13\].yc/din[1] blk.column\[4\].row\[13\].yc/dempty
+ blk.column\[4\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_262_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_399_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_304_ _302_/Y _298_/X wbs_dat_i[5] _303_/X VGND VGND VPWR VPWR _304_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_490_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_488_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_523_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_380_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_536_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_274_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_410_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_353_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_784_ wb_clk_i _784_/D VGND VGND VPWR VPWR _356_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_483_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_368_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_537_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[5\].yc blk.column\[13\].row\[5\].yc/cbitin blk.column\[13\].row\[6\].yc/cbitin
+ blk.column\[13\].row\[5\].yc/confclk blk.column\[13\].row\[6\].yc/confclk blk.column\[13\].row\[5\].yc/dempty
+ blk.column\[13\].row\[5\].yc/din[0] blk.column\[13\].row\[5\].yc/din[1] blk.column\[13\].row\[6\].yc/uin[0]
+ blk.column\[13\].row\[6\].yc/uin[1] blk.column\[13\].row\[5\].yc/hempty blk.column\[12\].row\[5\].yc/lempty
+ blk.column\[13\].row\[5\].yc/lempty blk.column\[13\].row\[5\].yc/lin[0] blk.column\[13\].row\[5\].yc/lin[1]
+ blk.column\[14\].row\[5\].yc/rin[0] blk.column\[14\].row\[5\].yc/rin[1] blk.column\[12\].row\[5\].yc/hempty
+ blk.column\[13\].row\[5\].yc/reset blk.column\[13\].row\[6\].yc/reset blk.column\[13\].row\[5\].yc/rin[0]
+ blk.column\[13\].row\[5\].yc/rin[1] blk.column\[12\].row\[5\].yc/lin[0] blk.column\[12\].row\[5\].yc/lin[1]
+ blk.column\[13\].row\[5\].yc/uempty blk.column\[13\].row\[5\].yc/uin[0] blk.column\[13\].row\[5\].yc/uin[1]
+ blk.column\[13\].row\[4\].yc/din[0] blk.column\[13\].row\[4\].yc/din[1] blk.column\[13\].row\[4\].yc/dempty
+ blk.column\[13\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_446_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_525_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[6\].yc blk.column\[4\].row\[6\].yc/cbitin blk.column\[4\].row\[7\].yc/cbitin
+ blk.column\[4\].row\[6\].yc/confclk blk.column\[4\].row\[7\].yc/confclk blk.column\[4\].row\[6\].yc/dempty
+ blk.column\[4\].row\[6\].yc/din[0] blk.column\[4\].row\[6\].yc/din[1] blk.column\[4\].row\[7\].yc/uin[0]
+ blk.column\[4\].row\[7\].yc/uin[1] blk.column\[4\].row\[6\].yc/hempty blk.column\[3\].row\[6\].yc/lempty
+ blk.column\[4\].row\[6\].yc/lempty blk.column\[4\].row\[6\].yc/lin[0] blk.column\[4\].row\[6\].yc/lin[1]
+ blk.column\[5\].row\[6\].yc/rin[0] blk.column\[5\].row\[6\].yc/rin[1] blk.column\[3\].row\[6\].yc/hempty
+ blk.column\[4\].row\[6\].yc/reset blk.column\[4\].row\[7\].yc/reset blk.column\[4\].row\[6\].yc/rin[0]
+ blk.column\[4\].row\[6\].yc/rin[1] blk.column\[3\].row\[6\].yc/lin[0] blk.column\[3\].row\[6\].yc/lin[1]
+ blk.column\[4\].row\[6\].yc/uempty blk.column\[4\].row\[6\].yc/uin[0] blk.column\[4\].row\[6\].yc/uin[1]
+ blk.column\[4\].row\[5\].yc/din[0] blk.column\[4\].row\[5\].yc/din[1] blk.column\[4\].row\[5\].yc/dempty
+ blk.column\[4\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_503_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_308_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_536_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_524_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_530_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_350_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_449_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_437_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_488_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_767_ wb_clk_i _394_/X VGND VGND VPWR VPWR wbs_dat_o[23] sky130_fd_sc_hd__dfxtp_4
XFILLER_483_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_450_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_507_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_507_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_698_ VGND VGND VPWR VPWR _698_/HI la_data_out[82] sky130_fd_sc_hd__conb_1
XFILLER_250_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_494_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_507_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_536_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_455_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[0\].yc la_data_in[105] blk.column\[9\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[9\].row\[1\].yc/confclk blk.column\[9\].row\[0\].yc/dempty blk.column\[9\].row\[0\].yc/din[0]
+ blk.column\[9\].row\[0\].yc/din[1] blk.column\[9\].row\[1\].yc/uin[0] blk.column\[9\].row\[1\].yc/uin[1]
+ blk.column\[9\].row\[0\].yc/hempty blk.column\[8\].row\[0\].yc/lempty blk.column\[9\].row\[0\].yc/lempty
+ blk.column\[9\].row\[0\].yc/lin[0] blk.column\[9\].row\[0\].yc/lin[1] blk.column\[9\].row\[0\].yc/lout[0]
+ blk.column\[9\].row\[0\].yc/lout[1] blk.column\[8\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[9\].row\[1\].yc/reset blk.column\[9\].row\[0\].yc/rin[0] blk.column\[9\].row\[0\].yc/rin[1]
+ blk.column\[8\].row\[0\].yc/lin[0] blk.column\[8\].row\[0\].yc/lin[1] _585_/LO la_data_in[82]
+ la_data_in[83] la_data_out[18] la_data_out[19] blk.column\[9\].row\[0\].yc/vempty
+ blk.column\[9\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_451_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_518_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_497_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_439_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_538_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_469_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_382_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_621_ VGND VGND VPWR VPWR _621_/HI io_oeb[33] sky130_fd_sc_hd__conb_1
XFILLER_523_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_504_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_552_ VGND VGND VPWR VPWR _552_/HI _552_/LO sky130_fd_sc_hd__conb_1
XFILLER_183_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_351_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_483_ VGND VGND VPWR VPWR _483_/HI _483_/LO sky130_fd_sc_hd__conb_1
XPHY_4887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_386_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_349_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_537_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_534_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_485_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_496_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_511_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_407_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_538_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_358_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_492_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_482_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_604_ VGND VGND VPWR VPWR _604_/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XPHY_6086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_535_ VGND VGND VPWR VPWR _535_/HI _535_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_466_ VGND VGND VPWR VPWR _466_/HI _466_/LO sky130_fd_sc_hd__conb_1
XPHY_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[11\].yc blk.column\[13\].row\[11\].yc/cbitin blk.column\[13\].row\[12\].yc/cbitin
+ blk.column\[13\].row\[11\].yc/confclk blk.column\[13\].row\[12\].yc/confclk blk.column\[13\].row\[11\].yc/dempty
+ blk.column\[13\].row\[11\].yc/din[0] blk.column\[13\].row\[11\].yc/din[1] blk.column\[13\].row\[12\].yc/uin[0]
+ blk.column\[13\].row\[12\].yc/uin[1] blk.column\[13\].row\[11\].yc/hempty blk.column\[12\].row\[11\].yc/lempty
+ blk.column\[13\].row\[11\].yc/lempty blk.column\[13\].row\[11\].yc/lin[0] blk.column\[13\].row\[11\].yc/lin[1]
+ blk.column\[14\].row\[11\].yc/rin[0] blk.column\[14\].row\[11\].yc/rin[1] blk.column\[12\].row\[11\].yc/hempty
+ blk.column\[13\].row\[11\].yc/reset blk.column\[13\].row\[12\].yc/reset blk.column\[13\].row\[11\].yc/rin[0]
+ blk.column\[13\].row\[11\].yc/rin[1] blk.column\[12\].row\[11\].yc/lin[0] blk.column\[12\].row\[11\].yc/lin[1]
+ blk.column\[13\].row\[11\].yc/uempty blk.column\[13\].row\[11\].yc/uin[0] blk.column\[13\].row\[11\].yc/uin[1]
+ blk.column\[13\].row\[10\].yc/din[0] blk.column\[13\].row\[10\].yc/din[1] blk.column\[13\].row\[10\].yc/dempty
+ blk.column\[13\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_397_ _391_/X wbs_dat_o[21] _344_/A _396_/X VGND VGND VPWR VPWR _397_/X sky130_fd_sc_hd__o22a_4
XFILLER_536_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[7\].yc blk.column\[14\].row\[7\].yc/cbitin blk.column\[14\].row\[8\].yc/cbitin
+ blk.column\[14\].row\[7\].yc/confclk blk.column\[14\].row\[8\].yc/confclk blk.column\[14\].row\[7\].yc/dempty
+ blk.column\[14\].row\[7\].yc/din[0] blk.column\[14\].row\[7\].yc/din[1] blk.column\[14\].row\[8\].yc/uin[0]
+ blk.column\[14\].row\[8\].yc/uin[1] blk.column\[14\].row\[7\].yc/hempty blk.column\[13\].row\[7\].yc/lempty
+ blk.column\[14\].row\[7\].yc/lempty blk.column\[14\].row\[7\].yc/lin[0] blk.column\[14\].row\[7\].yc/lin[1]
+ blk.column\[15\].row\[7\].yc/rin[0] blk.column\[15\].row\[7\].yc/rin[1] blk.column\[13\].row\[7\].yc/hempty
+ blk.column\[14\].row\[7\].yc/reset blk.column\[14\].row\[8\].yc/reset blk.column\[14\].row\[7\].yc/rin[0]
+ blk.column\[14\].row\[7\].yc/rin[1] blk.column\[13\].row\[7\].yc/lin[0] blk.column\[13\].row\[7\].yc/lin[1]
+ blk.column\[14\].row\[7\].yc/uempty blk.column\[14\].row\[7\].yc/uin[0] blk.column\[14\].row\[7\].yc/uin[1]
+ blk.column\[14\].row\[6\].yc/din[0] blk.column\[14\].row\[6\].yc/din[1] blk.column\[14\].row\[6\].yc/dempty
+ blk.column\[14\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_526_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_334_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_429_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[8\].yc blk.column\[5\].row\[8\].yc/cbitin blk.column\[5\].row\[9\].yc/cbitin
+ blk.column\[5\].row\[8\].yc/confclk blk.column\[5\].row\[9\].yc/confclk blk.column\[5\].row\[8\].yc/dempty
+ blk.column\[5\].row\[8\].yc/din[0] blk.column\[5\].row\[8\].yc/din[1] blk.column\[5\].row\[9\].yc/uin[0]
+ blk.column\[5\].row\[9\].yc/uin[1] blk.column\[5\].row\[8\].yc/hempty blk.column\[4\].row\[8\].yc/lempty
+ blk.column\[5\].row\[8\].yc/lempty blk.column\[5\].row\[8\].yc/lin[0] blk.column\[5\].row\[8\].yc/lin[1]
+ blk.column\[6\].row\[8\].yc/rin[0] blk.column\[6\].row\[8\].yc/rin[1] blk.column\[4\].row\[8\].yc/hempty
+ blk.column\[5\].row\[8\].yc/reset blk.column\[5\].row\[9\].yc/reset blk.column\[5\].row\[8\].yc/rin[0]
+ blk.column\[5\].row\[8\].yc/rin[1] blk.column\[4\].row\[8\].yc/lin[0] blk.column\[4\].row\[8\].yc/lin[1]
+ blk.column\[5\].row\[8\].yc/uempty blk.column\[5\].row\[8\].yc/uin[0] blk.column\[5\].row\[8\].yc/uin[1]
+ blk.column\[5\].row\[7\].yc/din[0] blk.column\[5\].row\[7\].yc/din[1] blk.column\[5\].row\[7\].yc/dempty
+ blk.column\[5\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_485_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_270_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_527_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_436_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_353_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_516_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_320_ _316_/Y _319_/X wbs_dat_i[15] _319_/X VGND VGND VPWR VPWR _320_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_401_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_505_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_346_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_316_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_237_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_518_ VGND VGND VPWR VPWR _518_/HI _518_/LO sky130_fd_sc_hd__conb_1
XFILLER_504_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_454_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_449_ VGND VGND VPWR VPWR _449_/HI _449_/LO sky130_fd_sc_hd__conb_1
XFILLER_337_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_493_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_436_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_512_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_524_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_432_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_492_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_515_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_251_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_530_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_303_ _298_/A VGND VGND VPWR VPWR _303_/X sky130_fd_sc_hd__buf_2
XFILLER_125_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_540_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[0\].row\[1\].yc blk.column\[0\].row\[1\].yc/cbitin blk.column\[0\].row\[2\].yc/cbitin
+ blk.column\[0\].row\[1\].yc/confclk blk.column\[0\].row\[2\].yc/confclk blk.column\[0\].row\[1\].yc/dempty
+ blk.column\[0\].row\[1\].yc/din[0] blk.column\[0\].row\[1\].yc/din[1] blk.column\[0\].row\[2\].yc/uin[0]
+ blk.column\[0\].row\[2\].yc/uin[1] blk.column\[0\].row\[1\].yc/hempty blk.column\[0\].row\[1\].yc/hempty2
+ blk.column\[0\].row\[1\].yc/lempty blk.column\[0\].row\[1\].yc/lin[0] blk.column\[0\].row\[1\].yc/lin[1]
+ blk.column\[1\].row\[1\].yc/rin[0] blk.column\[1\].row\[1\].yc/rin[1] _436_/HI blk.column\[0\].row\[1\].yc/reset
+ blk.column\[0\].row\[2\].yc/reset _493_/LO _494_/LO blk.column\[0\].row\[1\].yc/rout[0]
+ blk.column\[0\].row\[1\].yc/rout[1] blk.column\[0\].row\[1\].yc/uempty blk.column\[0\].row\[1\].yc/uin[0]
+ blk.column\[0\].row\[1\].yc/uin[1] blk.column\[0\].row\[0\].yc/din[0] blk.column\[0\].row\[0\].yc/din[1]
+ blk.column\[0\].row\[0\].yc/dempty blk.column\[0\].row\[2\].yc/uempty VPWR VGND
+ ycell
XFILLER_295_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_505_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_274_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_517_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[10\].yc blk.column\[1\].row\[9\].yc/cbitout blk.column\[1\].row\[11\].yc/cbitin
+ blk.column\[1\].row\[9\].yc/confclko blk.column\[1\].row\[11\].yc/confclk blk.column\[1\].row\[10\].yc/dempty
+ blk.column\[1\].row\[10\].yc/din[0] blk.column\[1\].row\[10\].yc/din[1] blk.column\[1\].row\[11\].yc/uin[0]
+ blk.column\[1\].row\[11\].yc/uin[1] blk.column\[1\].row\[10\].yc/hempty blk.column\[0\].row\[10\].yc/lempty
+ blk.column\[1\].row\[10\].yc/lempty blk.column\[1\].row\[10\].yc/lin[0] blk.column\[1\].row\[10\].yc/lin[1]
+ blk.column\[2\].row\[10\].yc/rin[0] blk.column\[2\].row\[10\].yc/rin[1] blk.column\[0\].row\[10\].yc/hempty
+ blk.column\[1\].row\[9\].yc/reseto blk.column\[1\].row\[11\].yc/reset blk.column\[1\].row\[10\].yc/rin[0]
+ blk.column\[1\].row\[10\].yc/rin[1] blk.column\[0\].row\[10\].yc/lin[0] blk.column\[0\].row\[10\].yc/lin[1]
+ blk.column\[1\].row\[9\].yc/vempty2 blk.column\[1\].row\[9\].yc/dout[0] blk.column\[1\].row\[9\].yc/dout[1]
+ blk.column\[1\].row\[9\].yc/din[0] blk.column\[1\].row\[9\].yc/din[1] blk.column\[1\].row\[9\].yc/dempty
+ blk.column\[1\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_170_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_410_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_417_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_437_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_538_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_542_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_531_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_535_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_783_ wb_clk_i _362_/X VGND VGND VPWR VPWR _358_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_147_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[9\].yc blk.column\[15\].row\[9\].yc/cbitin blk.column\[15\].row\[9\].yc/cbitout
+ blk.column\[15\].row\[9\].yc/confclk blk.column\[15\].row\[9\].yc/confclko blk.column\[15\].row\[9\].yc/dempty
+ blk.column\[15\].row\[9\].yc/din[0] blk.column\[15\].row\[9\].yc/din[1] blk.column\[15\].row\[9\].yc/dout[0]
+ blk.column\[15\].row\[9\].yc/dout[1] blk.column\[15\].row\[9\].yc/hempty blk.column\[14\].row\[9\].yc/lempty
+ _466_/HI _559_/LO _560_/LO blk.column\[15\].row\[9\].yc/lout[0] blk.column\[15\].row\[9\].yc/lout[1]
+ blk.column\[14\].row\[9\].yc/hempty blk.column\[15\].row\[9\].yc/reset blk.column\[15\].row\[9\].yc/reseto
+ blk.column\[15\].row\[9\].yc/rin[0] blk.column\[15\].row\[9\].yc/rin[1] blk.column\[14\].row\[9\].yc/lin[0]
+ blk.column\[14\].row\[9\].yc/lin[1] blk.column\[15\].row\[9\].yc/uempty blk.column\[15\].row\[9\].yc/uin[0]
+ blk.column\[15\].row\[9\].yc/uin[1] blk.column\[15\].row\[8\].yc/din[0] blk.column\[15\].row\[8\].yc/din[1]
+ blk.column\[15\].row\[8\].yc/dempty blk.column\[15\].row\[9\].yc/vempty2 VPWR VGND
+ ycell
XFILLER_215_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_490_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_534_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_534_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_317_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_265_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_514_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_444_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_530_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_460_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_437_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_488_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_531_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_507_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_766_ wb_clk_i _395_/X VGND VGND VPWR VPWR wbs_dat_o[22] sky130_fd_sc_hd__dfxtp_4
XFILLER_526_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_697_ VGND VGND VPWR VPWR _697_/HI la_data_out[81] sky130_fd_sc_hd__conb_1
XFILLER_379_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_531_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_514_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[2\].yc blk.column\[10\].row\[2\].yc/cbitin blk.column\[10\].row\[3\].yc/cbitin
+ blk.column\[10\].row\[2\].yc/confclk blk.column\[10\].row\[3\].yc/confclk blk.column\[10\].row\[2\].yc/dempty
+ blk.column\[10\].row\[2\].yc/din[0] blk.column\[10\].row\[2\].yc/din[1] blk.column\[10\].row\[3\].yc/uin[0]
+ blk.column\[10\].row\[3\].yc/uin[1] blk.column\[10\].row\[2\].yc/hempty blk.column\[9\].row\[2\].yc/lempty
+ blk.column\[10\].row\[2\].yc/lempty blk.column\[10\].row\[2\].yc/lin[0] blk.column\[10\].row\[2\].yc/lin[1]
+ blk.column\[11\].row\[2\].yc/rin[0] blk.column\[11\].row\[2\].yc/rin[1] blk.column\[9\].row\[2\].yc/hempty
+ blk.column\[10\].row\[2\].yc/reset blk.column\[10\].row\[3\].yc/reset blk.column\[9\].row\[2\].yc/lout[0]
+ blk.column\[9\].row\[2\].yc/lout[1] blk.column\[9\].row\[2\].yc/lin[0] blk.column\[9\].row\[2\].yc/lin[1]
+ blk.column\[10\].row\[2\].yc/uempty blk.column\[10\].row\[2\].yc/uin[0] blk.column\[10\].row\[2\].yc/uin[1]
+ blk.column\[10\].row\[1\].yc/din[0] blk.column\[10\].row\[1\].yc/din[1] blk.column\[10\].row\[1\].yc/dempty
+ blk.column\[10\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_85_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_323_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_489_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_620_ VGND VGND VPWR VPWR _620_/HI io_oeb[32] sky130_fd_sc_hd__conb_1
XPHY_6246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_527_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_382_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_523_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[1\].row\[3\].yc blk.column\[1\].row\[3\].yc/cbitin blk.column\[1\].row\[4\].yc/cbitin
+ blk.column\[1\].row\[3\].yc/confclk blk.column\[1\].row\[4\].yc/confclk blk.column\[1\].row\[3\].yc/dempty
+ blk.column\[1\].row\[3\].yc/din[0] blk.column\[1\].row\[3\].yc/din[1] blk.column\[1\].row\[4\].yc/uin[0]
+ blk.column\[1\].row\[4\].yc/uin[1] blk.column\[1\].row\[3\].yc/hempty blk.column\[0\].row\[3\].yc/lempty
+ blk.column\[1\].row\[3\].yc/lempty blk.column\[1\].row\[3\].yc/lin[0] blk.column\[1\].row\[3\].yc/lin[1]
+ blk.column\[2\].row\[3\].yc/rin[0] blk.column\[2\].row\[3\].yc/rin[1] blk.column\[0\].row\[3\].yc/hempty
+ blk.column\[1\].row\[3\].yc/reset blk.column\[1\].row\[4\].yc/reset blk.column\[1\].row\[3\].yc/rin[0]
+ blk.column\[1\].row\[3\].yc/rin[1] blk.column\[0\].row\[3\].yc/lin[0] blk.column\[0\].row\[3\].yc/lin[1]
+ blk.column\[1\].row\[3\].yc/uempty blk.column\[1\].row\[3\].yc/uin[0] blk.column\[1\].row\[3\].yc/uin[1]
+ blk.column\[1\].row\[2\].yc/din[0] blk.column\[1\].row\[2\].yc/din[1] blk.column\[1\].row\[2\].yc/dempty
+ blk.column\[1\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_508_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_551_ VGND VGND VPWR VPWR _551_/HI _551_/LO sky130_fd_sc_hd__conb_1
XPHY_5567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_482_ VGND VGND VPWR VPWR _482_/HI _482_/LO sky130_fd_sc_hd__conb_1
XPHY_4866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_519_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_515_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[5\].row\[13\].yc blk.column\[5\].row\[13\].yc/cbitin blk.column\[5\].row\[14\].yc/cbitin
+ blk.column\[5\].row\[13\].yc/confclk blk.column\[5\].row\[14\].yc/confclk blk.column\[5\].row\[13\].yc/dempty
+ blk.column\[5\].row\[13\].yc/din[0] blk.column\[5\].row\[13\].yc/din[1] blk.column\[5\].row\[14\].yc/uin[0]
+ blk.column\[5\].row\[14\].yc/uin[1] blk.column\[5\].row\[13\].yc/hempty blk.column\[4\].row\[13\].yc/lempty
+ blk.column\[5\].row\[13\].yc/lempty blk.column\[5\].row\[13\].yc/lin[0] blk.column\[5\].row\[13\].yc/lin[1]
+ blk.column\[6\].row\[13\].yc/rin[0] blk.column\[6\].row\[13\].yc/rin[1] blk.column\[4\].row\[13\].yc/hempty
+ blk.column\[5\].row\[13\].yc/reset blk.column\[5\].row\[14\].yc/reset blk.column\[5\].row\[13\].yc/rin[0]
+ blk.column\[5\].row\[13\].yc/rin[1] blk.column\[4\].row\[13\].yc/lin[0] blk.column\[4\].row\[13\].yc/lin[1]
+ blk.column\[5\].row\[13\].yc/uempty blk.column\[5\].row\[13\].yc/uin[0] blk.column\[5\].row\[13\].yc/uin[1]
+ blk.column\[5\].row\[12\].yc/din[0] blk.column\[5\].row\[12\].yc/din[1] blk.column\[5\].row\[12\].yc/dempty
+ blk.column\[5\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_168_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_409_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_749_ wb_clk_i _420_/X VGND VGND VPWR VPWR wbs_dat_o[5] sky130_fd_sc_hd__dfxtp_4
XFILLER_526_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_520_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_507_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_526_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_275_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_522_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_459_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_440_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_397_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_311_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_351_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_603_ VGND VGND VPWR VPWR _603_/HI io_oeb[15] sky130_fd_sc_hd__conb_1
XPHY_6076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_534_ VGND VGND VPWR VPWR _534_/HI _534_/LO sky130_fd_sc_hd__conb_1
XPHY_5386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_217_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_465_ VGND VGND VPWR VPWR _465_/HI _465_/LO sky130_fd_sc_hd__conb_1
XPHY_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_396_ _382_/A VGND VGND VPWR VPWR _396_/X sky130_fd_sc_hd__buf_2
XFILLER_417_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_488_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_325_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_487_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_452_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_429_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_214_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_249_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_527_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_505_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[12\].row\[15\].yc blk.column\[12\].row\[15\].yc/cbitin la_data_out[44]
+ blk.column\[12\].row\[15\].yc/confclk blk.column\[12\].row\[15\].yc/confclko _447_/HI
+ _518_/LO _519_/LO blk.column\[12\].row\[15\].yc/dout[0] blk.column\[12\].row\[15\].yc/dout[1]
+ blk.column\[12\].row\[15\].yc/hempty blk.column\[11\].row\[15\].yc/lempty blk.column\[12\].row\[15\].yc/lempty
+ blk.column\[12\].row\[15\].yc/lin[0] blk.column\[12\].row\[15\].yc/lin[1] blk.column\[13\].row\[15\].yc/rin[0]
+ blk.column\[13\].row\[15\].yc/rin[1] blk.column\[11\].row\[15\].yc/hempty blk.column\[12\].row\[15\].yc/reset
+ blk.column\[12\].row\[15\].yc/reseto blk.column\[12\].row\[15\].yc/rin[0] blk.column\[12\].row\[15\].yc/rin[1]
+ blk.column\[11\].row\[15\].yc/lin[0] blk.column\[11\].row\[15\].yc/lin[1] blk.column\[12\].row\[15\].yc/uempty
+ blk.column\[12\].row\[15\].yc/uin[0] blk.column\[12\].row\[15\].yc/uin[1] blk.column\[12\].row\[14\].yc/din[0]
+ blk.column\[12\].row\[14\].yc/din[1] blk.column\[12\].row\[14\].yc/dempty blk.column\[12\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_401_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_503_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_534_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_362_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_438_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_517_ VGND VGND VPWR VPWR _517_/HI _517_/LO sky130_fd_sc_hd__conb_1
XPHY_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ VGND VGND VPWR VPWR _448_/HI _448_/LO sky130_fd_sc_hd__conb_1
XFILLER_366_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_337_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_537_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_347_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_379_ _295_/Y VGND VGND VPWR VPWR _419_/A sky130_fd_sc_hd__buf_2
XFILLER_122_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_485_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[11\].row\[4\].yc blk.column\[11\].row\[4\].yc/cbitin blk.column\[11\].row\[5\].yc/cbitin
+ blk.column\[11\].row\[4\].yc/confclk blk.column\[11\].row\[5\].yc/confclk blk.column\[11\].row\[4\].yc/dempty
+ blk.column\[11\].row\[4\].yc/din[0] blk.column\[11\].row\[4\].yc/din[1] blk.column\[11\].row\[5\].yc/uin[0]
+ blk.column\[11\].row\[5\].yc/uin[1] blk.column\[11\].row\[4\].yc/hempty blk.column\[10\].row\[4\].yc/lempty
+ blk.column\[11\].row\[4\].yc/lempty blk.column\[11\].row\[4\].yc/lin[0] blk.column\[11\].row\[4\].yc/lin[1]
+ blk.column\[12\].row\[4\].yc/rin[0] blk.column\[12\].row\[4\].yc/rin[1] blk.column\[10\].row\[4\].yc/hempty
+ blk.column\[11\].row\[4\].yc/reset blk.column\[11\].row\[5\].yc/reset blk.column\[11\].row\[4\].yc/rin[0]
+ blk.column\[11\].row\[4\].yc/rin[1] blk.column\[10\].row\[4\].yc/lin[0] blk.column\[10\].row\[4\].yc/lin[1]
+ blk.column\[11\].row\[4\].yc/uempty blk.column\[11\].row\[4\].yc/uin[0] blk.column\[11\].row\[4\].yc/uin[1]
+ blk.column\[11\].row\[3\].yc/din[0] blk.column\[11\].row\[3\].yc/din[1] blk.column\[11\].row\[3\].yc/dempty
+ blk.column\[11\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_522_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_321_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[5\].yc blk.column\[2\].row\[5\].yc/cbitin blk.column\[2\].row\[6\].yc/cbitin
+ blk.column\[2\].row\[5\].yc/confclk blk.column\[2\].row\[6\].yc/confclk blk.column\[2\].row\[5\].yc/dempty
+ blk.column\[2\].row\[5\].yc/din[0] blk.column\[2\].row\[5\].yc/din[1] blk.column\[2\].row\[6\].yc/uin[0]
+ blk.column\[2\].row\[6\].yc/uin[1] blk.column\[2\].row\[5\].yc/hempty blk.column\[1\].row\[5\].yc/lempty
+ blk.column\[2\].row\[5\].yc/lempty blk.column\[2\].row\[5\].yc/lin[0] blk.column\[2\].row\[5\].yc/lin[1]
+ blk.column\[3\].row\[5\].yc/rin[0] blk.column\[3\].row\[5\].yc/rin[1] blk.column\[1\].row\[5\].yc/hempty
+ blk.column\[2\].row\[5\].yc/reset blk.column\[2\].row\[6\].yc/reset blk.column\[2\].row\[5\].yc/rin[0]
+ blk.column\[2\].row\[5\].yc/rin[1] blk.column\[1\].row\[5\].yc/lin[0] blk.column\[1\].row\[5\].yc/lin[1]
+ blk.column\[2\].row\[5\].yc/uempty blk.column\[2\].row\[5\].yc/uin[0] blk.column\[2\].row\[5\].yc/uin[1]
+ blk.column\[2\].row\[4\].yc/din[0] blk.column\[2\].row\[4\].yc/din[1] blk.column\[2\].row\[4\].yc/dempty
+ blk.column\[2\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_483_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_522_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ _805_/Q VGND VGND VPWR VPWR _302_/Y sky130_fd_sc_hd__inv_2
XFILLER_518_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_371_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_506_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_398_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_508_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_385_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_407_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_327_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_782_ wb_clk_i _782_/D VGND VGND VPWR VPWR _363_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_112_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_374_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_507_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_520_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_414_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[14\].yc blk.column\[0\].row\[14\].yc/cbitin blk.column\[0\].row\[15\].yc/cbitin
+ blk.column\[0\].row\[14\].yc/confclk blk.column\[0\].row\[15\].yc/confclk blk.column\[0\].row\[14\].yc/dempty
+ blk.column\[0\].row\[14\].yc/din[0] blk.column\[0\].row\[14\].yc/din[1] blk.column\[0\].row\[15\].yc/uin[0]
+ blk.column\[0\].row\[15\].yc/uin[1] blk.column\[0\].row\[14\].yc/hempty blk.column\[0\].row\[14\].yc/hempty2
+ blk.column\[0\].row\[14\].yc/lempty blk.column\[0\].row\[14\].yc/lin[0] blk.column\[0\].row\[14\].yc/lin[1]
+ blk.column\[1\].row\[14\].yc/rin[0] blk.column\[1\].row\[14\].yc/rin[1] _433_/HI
+ blk.column\[0\].row\[14\].yc/reset blk.column\[0\].row\[15\].yc/reset _487_/LO _488_/LO
+ blk.column\[0\].row\[14\].yc/rout[0] blk.column\[0\].row\[14\].yc/rout[1] blk.column\[0\].row\[14\].yc/uempty
+ blk.column\[0\].row\[14\].yc/uin[0] blk.column\[0\].row\[14\].yc/uin[1] blk.column\[0\].row\[13\].yc/din[0]
+ blk.column\[0\].row\[13\].yc/din[1] blk.column\[0\].row\[13\].yc/dempty blk.column\[0\].row\[15\].yc/uempty
+ VPWR VGND ycell
XFILLER_332_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_488_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_484_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_345_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[10\].yc blk.column\[14\].row\[9\].yc/cbitout blk.column\[14\].row\[11\].yc/cbitin
+ blk.column\[14\].row\[9\].yc/confclko blk.column\[14\].row\[11\].yc/confclk blk.column\[14\].row\[10\].yc/dempty
+ blk.column\[14\].row\[10\].yc/din[0] blk.column\[14\].row\[10\].yc/din[1] blk.column\[14\].row\[11\].yc/uin[0]
+ blk.column\[14\].row\[11\].yc/uin[1] blk.column\[14\].row\[10\].yc/hempty blk.column\[13\].row\[10\].yc/lempty
+ blk.column\[14\].row\[10\].yc/lempty blk.column\[14\].row\[10\].yc/lin[0] blk.column\[14\].row\[10\].yc/lin[1]
+ blk.column\[15\].row\[10\].yc/rin[0] blk.column\[15\].row\[10\].yc/rin[1] blk.column\[13\].row\[10\].yc/hempty
+ blk.column\[14\].row\[9\].yc/reseto blk.column\[14\].row\[11\].yc/reset blk.column\[14\].row\[10\].yc/rin[0]
+ blk.column\[14\].row\[10\].yc/rin[1] blk.column\[13\].row\[10\].yc/lin[0] blk.column\[13\].row\[10\].yc/lin[1]
+ blk.column\[14\].row\[9\].yc/vempty2 blk.column\[14\].row\[9\].yc/dout[0] blk.column\[14\].row\[9\].yc/dout[1]
+ blk.column\[14\].row\[9\].yc/din[0] blk.column\[14\].row\[9\].yc/din[1] blk.column\[14\].row\[9\].yc/dempty
+ blk.column\[14\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_147_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_536_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_525_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_460_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_488_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_531_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_352_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_765_ wb_clk_i _397_/X VGND VGND VPWR VPWR wbs_dat_o[21] sky130_fd_sc_hd__dfxtp_4
XPHY_6973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_450_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_696_ VGND VGND VPWR VPWR _696_/HI la_data_out[80] sky130_fd_sc_hd__conb_1
XFILLER_235_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_483_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_250_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[6\].yc blk.column\[12\].row\[6\].yc/cbitin blk.column\[12\].row\[7\].yc/cbitin
+ blk.column\[12\].row\[6\].yc/confclk blk.column\[12\].row\[7\].yc/confclk blk.column\[12\].row\[6\].yc/dempty
+ blk.column\[12\].row\[6\].yc/din[0] blk.column\[12\].row\[6\].yc/din[1] blk.column\[12\].row\[7\].yc/uin[0]
+ blk.column\[12\].row\[7\].yc/uin[1] blk.column\[12\].row\[6\].yc/hempty blk.column\[11\].row\[6\].yc/lempty
+ blk.column\[12\].row\[6\].yc/lempty blk.column\[12\].row\[6\].yc/lin[0] blk.column\[12\].row\[6\].yc/lin[1]
+ blk.column\[13\].row\[6\].yc/rin[0] blk.column\[13\].row\[6\].yc/rin[1] blk.column\[11\].row\[6\].yc/hempty
+ blk.column\[12\].row\[6\].yc/reset blk.column\[12\].row\[7\].yc/reset blk.column\[12\].row\[6\].yc/rin[0]
+ blk.column\[12\].row\[6\].yc/rin[1] blk.column\[11\].row\[6\].yc/lin[0] blk.column\[11\].row\[6\].yc/lin[1]
+ blk.column\[12\].row\[6\].yc/uempty blk.column\[12\].row\[6\].yc/uin[0] blk.column\[12\].row\[6\].yc/uin[1]
+ blk.column\[12\].row\[5\].yc/din[0] blk.column\[12\].row\[5\].yc/din[1] blk.column\[12\].row\[5\].yc/dempty
+ blk.column\[12\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_503_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_323_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_542_3194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_395_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_499_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[7\].yc blk.column\[3\].row\[7\].yc/cbitin blk.column\[3\].row\[8\].yc/cbitin
+ blk.column\[3\].row\[7\].yc/confclk blk.column\[3\].row\[8\].yc/confclk blk.column\[3\].row\[7\].yc/dempty
+ blk.column\[3\].row\[7\].yc/din[0] blk.column\[3\].row\[7\].yc/din[1] blk.column\[3\].row\[8\].yc/uin[0]
+ blk.column\[3\].row\[8\].yc/uin[1] blk.column\[3\].row\[7\].yc/hempty blk.column\[2\].row\[7\].yc/lempty
+ blk.column\[3\].row\[7\].yc/lempty blk.column\[3\].row\[7\].yc/lin[0] blk.column\[3\].row\[7\].yc/lin[1]
+ blk.column\[4\].row\[7\].yc/rin[0] blk.column\[4\].row\[7\].yc/rin[1] blk.column\[2\].row\[7\].yc/hempty
+ blk.column\[3\].row\[7\].yc/reset blk.column\[3\].row\[8\].yc/reset blk.column\[3\].row\[7\].yc/rin[0]
+ blk.column\[3\].row\[7\].yc/rin[1] blk.column\[2\].row\[7\].yc/lin[0] blk.column\[2\].row\[7\].yc/lin[1]
+ blk.column\[3\].row\[7\].yc/uempty blk.column\[3\].row\[7\].yc/uin[0] blk.column\[3\].row\[7\].yc/uin[1]
+ blk.column\[3\].row\[6\].yc/din[0] blk.column\[3\].row\[6\].yc/din[1] blk.column\[3\].row\[6\].yc/dempty
+ blk.column\[3\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_536_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_516_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_10906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_248_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_508_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_328_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_480_2547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_550_ VGND VGND VPWR VPWR _550_/HI _550_/LO sky130_fd_sc_hd__conb_1
XFILLER_480_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_398_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_481_ VGND VGND VPWR VPWR _481_/HI _481_/LO sky130_fd_sc_hd__conb_1
XPHY_4856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_491_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_485_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_748_ wb_clk_i _748_/D VGND VGND VPWR VPWR wbs_dat_o[4] sky130_fd_sc_hd__dfxtp_4
XFILLER_162_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_542_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_679_ VGND VGND VPWR VPWR _679_/HI la_data_out[63] sky130_fd_sc_hd__conb_1
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_345_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[1\].yc blk.column\[8\].row\[1\].yc/cbitin blk.column\[8\].row\[2\].yc/cbitin
+ blk.column\[8\].row\[1\].yc/confclk blk.column\[8\].row\[2\].yc/confclk blk.column\[8\].row\[1\].yc/dempty
+ blk.column\[8\].row\[1\].yc/din[0] blk.column\[8\].row\[1\].yc/din[1] blk.column\[8\].row\[2\].yc/uin[0]
+ blk.column\[8\].row\[2\].yc/uin[1] blk.column\[8\].row\[1\].yc/hempty blk.column\[7\].row\[1\].yc/lempty
+ blk.column\[8\].row\[1\].yc/lempty blk.column\[8\].row\[1\].yc/lin[0] blk.column\[8\].row\[1\].yc/lin[1]
+ blk.column\[9\].row\[1\].yc/rin[0] blk.column\[9\].row\[1\].yc/rin[1] blk.column\[7\].row\[1\].yc/hempty
+ blk.column\[8\].row\[1\].yc/reset blk.column\[8\].row\[2\].yc/reset blk.column\[8\].row\[1\].yc/rin[0]
+ blk.column\[8\].row\[1\].yc/rin[1] blk.column\[7\].row\[1\].yc/lin[0] blk.column\[7\].row\[1\].yc/lin[1]
+ blk.column\[8\].row\[1\].yc/uempty blk.column\[8\].row\[1\].yc/uin[0] blk.column\[8\].row\[1\].yc/uin[1]
+ blk.column\[8\].row\[0\].yc/din[0] blk.column\[8\].row\[0\].yc/din[1] blk.column\[8\].row\[0\].yc/dempty
+ blk.column\[8\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_208_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_488_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_509_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_360_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_397_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_538_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_541_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_602_ VGND VGND VPWR VPWR _602_/HI io_oeb[14] sky130_fd_sc_hd__conb_1
XFILLER_431_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_533_ VGND VGND VPWR VPWR _533_/HI _533_/LO sky130_fd_sc_hd__conb_1
XPHY_5387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_359_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_464_ VGND VGND VPWR VPWR _464_/HI _464_/LO sky130_fd_sc_hd__conb_1
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_374_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_395_ _391_/X wbs_dat_o[22] _790_/Q _389_/X VGND VGND VPWR VPWR _395_/X sky130_fd_sc_hd__o22a_4
XPHY_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_489_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_341_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_498_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_517_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_533_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_511_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_251_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_509_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_403_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_475_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_436_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_512_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_309_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_343_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_516_ VGND VGND VPWR VPWR _516_/HI _516_/LO sky130_fd_sc_hd__conb_1
XFILLER_260_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_447_ VGND VGND VPWR VPWR _447_/HI _447_/LO sky130_fd_sc_hd__conb_1
XPHY_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_378_ _377_/Y _373_/X wbs_dat_i[24] _361_/A VGND VGND VPWR VPWR _378_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_374_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[8\].yc blk.column\[13\].row\[8\].yc/cbitin blk.column\[13\].row\[9\].yc/cbitin
+ blk.column\[13\].row\[8\].yc/confclk blk.column\[13\].row\[9\].yc/confclk blk.column\[13\].row\[8\].yc/dempty
+ blk.column\[13\].row\[8\].yc/din[0] blk.column\[13\].row\[8\].yc/din[1] blk.column\[13\].row\[9\].yc/uin[0]
+ blk.column\[13\].row\[9\].yc/uin[1] blk.column\[13\].row\[8\].yc/hempty blk.column\[12\].row\[8\].yc/lempty
+ blk.column\[13\].row\[8\].yc/lempty blk.column\[13\].row\[8\].yc/lin[0] blk.column\[13\].row\[8\].yc/lin[1]
+ blk.column\[14\].row\[8\].yc/rin[0] blk.column\[14\].row\[8\].yc/rin[1] blk.column\[12\].row\[8\].yc/hempty
+ blk.column\[13\].row\[8\].yc/reset blk.column\[13\].row\[9\].yc/reset blk.column\[13\].row\[8\].yc/rin[0]
+ blk.column\[13\].row\[8\].yc/rin[1] blk.column\[12\].row\[8\].yc/lin[0] blk.column\[12\].row\[8\].yc/lin[1]
+ blk.column\[13\].row\[8\].yc/uempty blk.column\[13\].row\[8\].yc/uin[0] blk.column\[13\].row\[8\].yc/uin[1]
+ blk.column\[13\].row\[7\].yc/din[0] blk.column\[13\].row\[7\].yc/din[1] blk.column\[13\].row\[7\].yc/dempty
+ blk.column\[13\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_512_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[9\].yc blk.column\[4\].row\[9\].yc/cbitin blk.column\[4\].row\[9\].yc/cbitout
+ blk.column\[4\].row\[9\].yc/confclk blk.column\[4\].row\[9\].yc/confclko blk.column\[4\].row\[9\].yc/dempty
+ blk.column\[4\].row\[9\].yc/din[0] blk.column\[4\].row\[9\].yc/din[1] blk.column\[4\].row\[9\].yc/dout[0]
+ blk.column\[4\].row\[9\].yc/dout[1] blk.column\[4\].row\[9\].yc/hempty blk.column\[3\].row\[9\].yc/lempty
+ blk.column\[4\].row\[9\].yc/lempty blk.column\[4\].row\[9\].yc/lin[0] blk.column\[4\].row\[9\].yc/lin[1]
+ blk.column\[5\].row\[9\].yc/rin[0] blk.column\[5\].row\[9\].yc/rin[1] blk.column\[3\].row\[9\].yc/hempty
+ blk.column\[4\].row\[9\].yc/reset blk.column\[4\].row\[9\].yc/reseto blk.column\[4\].row\[9\].yc/rin[0]
+ blk.column\[4\].row\[9\].yc/rin[1] blk.column\[3\].row\[9\].yc/lin[0] blk.column\[3\].row\[9\].yc/lin[1]
+ blk.column\[4\].row\[9\].yc/uempty blk.column\[4\].row\[9\].yc/uin[0] blk.column\[4\].row\[9\].yc/uin[1]
+ blk.column\[4\].row\[8\].yc/din[0] blk.column\[4\].row\[8\].yc/din[1] blk.column\[4\].row\[8\].yc/dempty
+ blk.column\[4\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_541_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_528_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_495_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_2635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_505_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_301_ _300_/Y _298_/X wbs_dat_i[6] _298_/X VGND VGND VPWR VPWR _806_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_479_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_497_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_417_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_537_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[9\].row\[3\].yc blk.column\[9\].row\[3\].yc/cbitin blk.column\[9\].row\[4\].yc/cbitin
+ blk.column\[9\].row\[3\].yc/confclk blk.column\[9\].row\[4\].yc/confclk blk.column\[9\].row\[3\].yc/dempty
+ blk.column\[9\].row\[3\].yc/din[0] blk.column\[9\].row\[3\].yc/din[1] blk.column\[9\].row\[4\].yc/uin[0]
+ blk.column\[9\].row\[4\].yc/uin[1] blk.column\[9\].row\[3\].yc/hempty blk.column\[8\].row\[3\].yc/lempty
+ blk.column\[9\].row\[3\].yc/lempty blk.column\[9\].row\[3\].yc/lin[0] blk.column\[9\].row\[3\].yc/lin[1]
+ blk.column\[9\].row\[3\].yc/lout[0] blk.column\[9\].row\[3\].yc/lout[1] blk.column\[8\].row\[3\].yc/hempty
+ blk.column\[9\].row\[3\].yc/reset blk.column\[9\].row\[4\].yc/reset blk.column\[9\].row\[3\].yc/rin[0]
+ blk.column\[9\].row\[3\].yc/rin[1] blk.column\[8\].row\[3\].yc/lin[0] blk.column\[8\].row\[3\].yc/lin[1]
+ blk.column\[9\].row\[3\].yc/uempty blk.column\[9\].row\[3\].yc/uin[0] blk.column\[9\].row\[3\].yc/uin[1]
+ blk.column\[9\].row\[2\].yc/din[0] blk.column\[9\].row\[2\].yc/din[1] blk.column\[9\].row\[2\].yc/dempty
+ blk.column\[9\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_18_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_493_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_350_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[12\].yc blk.column\[6\].row\[12\].yc/cbitin blk.column\[6\].row\[13\].yc/cbitin
+ blk.column\[6\].row\[12\].yc/confclk blk.column\[6\].row\[13\].yc/confclk blk.column\[6\].row\[12\].yc/dempty
+ blk.column\[6\].row\[12\].yc/din[0] blk.column\[6\].row\[12\].yc/din[1] blk.column\[6\].row\[13\].yc/uin[0]
+ blk.column\[6\].row\[13\].yc/uin[1] blk.column\[6\].row\[12\].yc/hempty blk.column\[5\].row\[12\].yc/lempty
+ blk.column\[6\].row\[12\].yc/lempty blk.column\[6\].row\[12\].yc/lin[0] blk.column\[6\].row\[12\].yc/lin[1]
+ blk.column\[7\].row\[12\].yc/rin[0] blk.column\[7\].row\[12\].yc/rin[1] blk.column\[5\].row\[12\].yc/hempty
+ blk.column\[6\].row\[12\].yc/reset blk.column\[6\].row\[13\].yc/reset blk.column\[6\].row\[12\].yc/rin[0]
+ blk.column\[6\].row\[12\].yc/rin[1] blk.column\[5\].row\[12\].yc/lin[0] blk.column\[5\].row\[12\].yc/lin[1]
+ blk.column\[6\].row\[12\].yc/uempty blk.column\[6\].row\[12\].yc/uin[0] blk.column\[6\].row\[12\].yc/uin[1]
+ blk.column\[6\].row\[11\].yc/din[0] blk.column\[6\].row\[11\].yc/din[1] blk.column\[6\].row\[11\].yc/dempty
+ blk.column\[6\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_5_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_481_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_502_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_476_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_498_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_494_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_538_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_517_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_407_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_327_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_781_ wb_clk_i _781_/D VGND VGND VPWR VPWR _365_/A sky130_fd_sc_hd__dfxtp_4
XPHY_7867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_540_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_519_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_518_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_448_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_418_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_530_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_454_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_345_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_520_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_536_2402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_367_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_358_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_512_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_326_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_420_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_396_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_292_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_352_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_764_ wb_clk_i _764_/D VGND VGND VPWR VPWR wbs_dat_o[20] sky130_fd_sc_hd__dfxtp_4
XPHY_7697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_451_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_695_ VGND VGND VPWR VPWR _695_/HI la_data_out[79] sky130_fd_sc_hd__conb_1
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[14\].yc blk.column\[13\].row\[14\].yc/cbitin blk.column\[13\].row\[15\].yc/cbitin
+ blk.column\[13\].row\[14\].yc/confclk blk.column\[13\].row\[15\].yc/confclk blk.column\[13\].row\[14\].yc/dempty
+ blk.column\[13\].row\[14\].yc/din[0] blk.column\[13\].row\[14\].yc/din[1] blk.column\[13\].row\[15\].yc/uin[0]
+ blk.column\[13\].row\[15\].yc/uin[1] blk.column\[13\].row\[14\].yc/hempty blk.column\[12\].row\[14\].yc/lempty
+ blk.column\[13\].row\[14\].yc/lempty blk.column\[13\].row\[14\].yc/lin[0] blk.column\[13\].row\[14\].yc/lin[1]
+ blk.column\[14\].row\[14\].yc/rin[0] blk.column\[14\].row\[14\].yc/rin[1] blk.column\[12\].row\[14\].yc/hempty
+ blk.column\[13\].row\[14\].yc/reset blk.column\[13\].row\[15\].yc/reset blk.column\[13\].row\[14\].yc/rin[0]
+ blk.column\[13\].row\[14\].yc/rin[1] blk.column\[12\].row\[14\].yc/lin[0] blk.column\[12\].row\[14\].yc/lin[1]
+ blk.column\[13\].row\[14\].yc/uempty blk.column\[13\].row\[14\].yc/uin[0] blk.column\[13\].row\[14\].yc/uin[1]
+ blk.column\[13\].row\[13\].yc/din[0] blk.column\[13\].row\[13\].yc/din[1] blk.column\[13\].row\[13\].yc/dempty
+ blk.column\[13\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_379_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_305_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_522_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_521_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_479_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_434_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_455_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_252_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_418_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_480_ VGND VGND VPWR VPWR _480_/HI _480_/LO sky130_fd_sc_hd__conb_1
XPHY_4857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_478_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_346_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_335_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_513_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_747_ wb_clk_i _747_/D VGND VGND VPWR VPWR wbs_dat_o[3] sky130_fd_sc_hd__dfxtp_4
XPHY_6782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_678_ VGND VGND VPWR VPWR _678_/HI la_data_out[62] sky130_fd_sc_hd__conb_1
XFILLER_524_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_339_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_397_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_473_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_328_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_293_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_532_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_330_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_601_ VGND VGND VPWR VPWR _601_/HI io_oeb[13] sky130_fd_sc_hd__conb_1
XPHY_6056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_532_ VGND VGND VPWR VPWR _532_/HI _532_/LO sky130_fd_sc_hd__conb_1
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_463_ VGND VGND VPWR VPWR _463_/HI _463_/LO sky130_fd_sc_hd__conb_1
XPHY_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[0\].row\[4\].yc blk.column\[0\].row\[4\].yc/cbitin blk.column\[0\].row\[5\].yc/cbitin
+ blk.column\[0\].row\[4\].yc/confclk blk.column\[0\].row\[5\].yc/confclk blk.column\[0\].row\[4\].yc/dempty
+ blk.column\[0\].row\[4\].yc/din[0] blk.column\[0\].row\[4\].yc/din[1] blk.column\[0\].row\[5\].yc/uin[0]
+ blk.column\[0\].row\[5\].yc/uin[1] blk.column\[0\].row\[4\].yc/hempty blk.column\[0\].row\[4\].yc/hempty2
+ blk.column\[0\].row\[4\].yc/lempty blk.column\[0\].row\[4\].yc/lin[0] blk.column\[0\].row\[4\].yc/lin[1]
+ blk.column\[1\].row\[4\].yc/rin[0] blk.column\[1\].row\[4\].yc/rin[1] _439_/HI blk.column\[0\].row\[4\].yc/reset
+ blk.column\[0\].row\[5\].yc/reset _499_/LO _500_/LO blk.column\[0\].row\[4\].yc/rout[0]
+ blk.column\[0\].row\[4\].yc/rout[1] blk.column\[0\].row\[4\].yc/uempty blk.column\[0\].row\[4\].yc/uin[0]
+ blk.column\[0\].row\[4\].yc/uin[1] blk.column\[0\].row\[3\].yc/din[0] blk.column\[0\].row\[3\].yc/din[1]
+ blk.column\[0\].row\[4\].yc/vempty blk.column\[0\].row\[5\].yc/uempty VPWR VGND
+ ycell
XPHY_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_359_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_394_ _391_/X wbs_dat_o[23] _337_/A _389_/X VGND VGND VPWR VPWR _394_/X sky130_fd_sc_hd__o22a_4
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_417_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_392_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_469_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_500_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_485_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_238_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_318_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[13\].yc blk.column\[1\].row\[13\].yc/cbitin blk.column\[1\].row\[14\].yc/cbitin
+ blk.column\[1\].row\[13\].yc/confclk blk.column\[1\].row\[14\].yc/confclk blk.column\[1\].row\[13\].yc/dempty
+ blk.column\[1\].row\[13\].yc/din[0] blk.column\[1\].row\[13\].yc/din[1] blk.column\[1\].row\[14\].yc/uin[0]
+ blk.column\[1\].row\[14\].yc/uin[1] blk.column\[1\].row\[13\].yc/hempty blk.column\[0\].row\[13\].yc/lempty
+ blk.column\[1\].row\[13\].yc/lempty blk.column\[1\].row\[13\].yc/lin[0] blk.column\[1\].row\[13\].yc/lin[1]
+ blk.column\[2\].row\[13\].yc/rin[0] blk.column\[2\].row\[13\].yc/rin[1] blk.column\[0\].row\[13\].yc/hempty
+ blk.column\[1\].row\[13\].yc/reset blk.column\[1\].row\[14\].yc/reset blk.column\[1\].row\[13\].yc/rin[0]
+ blk.column\[1\].row\[13\].yc/rin[1] blk.column\[0\].row\[13\].yc/lin[0] blk.column\[0\].row\[13\].yc/lin[1]
+ blk.column\[1\].row\[13\].yc/uempty blk.column\[1\].row\[13\].yc/uin[0] blk.column\[1\].row\[13\].yc/uin[1]
+ blk.column\[1\].row\[12\].yc/din[0] blk.column\[1\].row\[12\].yc/din[1] blk.column\[1\].row\[12\].yc/dempty
+ blk.column\[1\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_380_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_388_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_540_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_470_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_403_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_477_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_356_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_516_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_296_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_397_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_382_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_486_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_515_ VGND VGND VPWR VPWR _515_/HI _515_/LO sky130_fd_sc_hd__conb_1
XFILLER_480_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_446_ VGND VGND VPWR VPWR _446_/HI _446_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_376_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_395_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_377_ _776_/Q VGND VGND VPWR VPWR _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_536_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_347_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_436_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_313_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_506_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_504_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_527_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_300_ _806_/Q VGND VGND VPWR VPWR _300_/Y sky130_fd_sc_hd__inv_2
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_295_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_371_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_516_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_542_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_488_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_473_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_527_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_507_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_343_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_419_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_429_ VGND VGND VPWR VPWR _429_/HI _429_/LO sky130_fd_sc_hd__conb_1
XFILLER_15_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_2639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_315_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_432_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[5\].yc blk.column\[10\].row\[5\].yc/cbitin blk.column\[10\].row\[6\].yc/cbitin
+ blk.column\[10\].row\[5\].yc/confclk blk.column\[10\].row\[6\].yc/confclk blk.column\[10\].row\[5\].yc/dempty
+ blk.column\[10\].row\[5\].yc/din[0] blk.column\[10\].row\[5\].yc/din[1] blk.column\[10\].row\[6\].yc/uin[0]
+ blk.column\[10\].row\[6\].yc/uin[1] blk.column\[10\].row\[5\].yc/hempty blk.column\[9\].row\[5\].yc/lempty
+ blk.column\[10\].row\[5\].yc/lempty blk.column\[10\].row\[5\].yc/lin[0] blk.column\[10\].row\[5\].yc/lin[1]
+ blk.column\[11\].row\[5\].yc/rin[0] blk.column\[11\].row\[5\].yc/rin[1] blk.column\[9\].row\[5\].yc/hempty
+ blk.column\[10\].row\[5\].yc/reset blk.column\[10\].row\[6\].yc/reset blk.column\[9\].row\[5\].yc/lout[0]
+ blk.column\[9\].row\[5\].yc/lout[1] blk.column\[9\].row\[5\].yc/lin[0] blk.column\[9\].row\[5\].yc/lin[1]
+ blk.column\[10\].row\[5\].yc/uempty blk.column\[10\].row\[5\].yc/uin[0] blk.column\[10\].row\[5\].yc/uin[1]
+ blk.column\[10\].row\[4\].yc/din[0] blk.column\[10\].row\[4\].yc/din[1] blk.column\[10\].row\[4\].yc/dempty
+ blk.column\[10\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_535_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_326_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_257_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_257_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_419_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_780_ wb_clk_i _369_/X VGND VGND VPWR VPWR _780_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_5_2444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[6\].yc blk.column\[1\].row\[6\].yc/cbitin blk.column\[1\].row\[7\].yc/cbitin
+ blk.column\[1\].row\[6\].yc/confclk blk.column\[1\].row\[7\].yc/confclk blk.column\[1\].row\[6\].yc/dempty
+ blk.column\[1\].row\[6\].yc/din[0] blk.column\[1\].row\[6\].yc/din[1] blk.column\[1\].row\[7\].yc/uin[0]
+ blk.column\[1\].row\[7\].yc/uin[1] blk.column\[1\].row\[6\].yc/hempty blk.column\[0\].row\[6\].yc/lempty
+ blk.column\[1\].row\[6\].yc/lempty blk.column\[1\].row\[6\].yc/lin[0] blk.column\[1\].row\[6\].yc/lin[1]
+ blk.column\[2\].row\[6\].yc/rin[0] blk.column\[2\].row\[6\].yc/rin[1] blk.column\[0\].row\[6\].yc/hempty
+ blk.column\[1\].row\[6\].yc/reset blk.column\[1\].row\[7\].yc/reset blk.column\[1\].row\[6\].yc/rin[0]
+ blk.column\[1\].row\[6\].yc/rin[1] blk.column\[0\].row\[6\].yc/lin[0] blk.column\[0\].row\[6\].yc/lin[1]
+ blk.column\[1\].row\[6\].yc/uempty blk.column\[1\].row\[6\].yc/uin[0] blk.column\[1\].row\[6\].yc/uin[1]
+ blk.column\[1\].row\[5\].yc/din[0] blk.column\[1\].row\[5\].yc/din[1] blk.column\[1\].row\[5\].yc/dempty
+ blk.column\[1\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_491_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_2499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_373_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_497_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_384_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_238_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_460_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_335_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_493_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_239_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[0\].yc la_data_in[102] blk.column\[6\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[6\].row\[1\].yc/confclk blk.column\[6\].row\[0\].yc/dempty blk.column\[6\].row\[0\].yc/din[0]
+ blk.column\[6\].row\[0\].yc/din[1] blk.column\[6\].row\[1\].yc/uin[0] blk.column\[6\].row\[1\].yc/uin[1]
+ blk.column\[6\].row\[0\].yc/hempty blk.column\[5\].row\[0\].yc/lempty blk.column\[6\].row\[0\].yc/lempty
+ blk.column\[6\].row\[0\].yc/lin[0] blk.column\[6\].row\[0\].yc/lin[1] blk.column\[7\].row\[0\].yc/rin[0]
+ blk.column\[7\].row\[0\].yc/rin[1] blk.column\[5\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[6\].row\[1\].yc/reset blk.column\[6\].row\[0\].yc/rin[0] blk.column\[6\].row\[0\].yc/rin[1]
+ blk.column\[5\].row\[0\].yc/lin[0] blk.column\[5\].row\[0\].yc/lin[1] _576_/LO la_data_in[76]
+ la_data_in[77] la_data_out[12] la_data_out[13] blk.column\[6\].row\[0\].yc/vempty
+ blk.column\[6\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_181_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_358_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_292_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_763_ wb_clk_i _400_/X VGND VGND VPWR VPWR wbs_dat_o[19] sky130_fd_sc_hd__dfxtp_4
XFILLER_153_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_694_ VGND VGND VPWR VPWR _694_/HI la_data_out[78] sky130_fd_sc_hd__conb_1
XFILLER_21_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_526_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_340_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_317_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_514_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_522_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_482_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_507_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_410_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_540_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[10\].yc blk.column\[10\].row\[9\].yc/cbitout blk.column\[10\].row\[11\].yc/cbitin
+ blk.column\[10\].row\[9\].yc/confclko blk.column\[10\].row\[11\].yc/confclk blk.column\[10\].row\[10\].yc/dempty
+ blk.column\[10\].row\[10\].yc/din[0] blk.column\[10\].row\[10\].yc/din[1] blk.column\[10\].row\[11\].yc/uin[0]
+ blk.column\[10\].row\[11\].yc/uin[1] blk.column\[10\].row\[10\].yc/hempty blk.column\[9\].row\[10\].yc/lempty
+ blk.column\[10\].row\[10\].yc/lempty blk.column\[10\].row\[10\].yc/lin[0] blk.column\[10\].row\[10\].yc/lin[1]
+ blk.column\[11\].row\[10\].yc/rin[0] blk.column\[11\].row\[10\].yc/rin[1] blk.column\[9\].row\[10\].yc/hempty
+ blk.column\[10\].row\[9\].yc/reseto blk.column\[10\].row\[11\].yc/reset blk.column\[9\].row\[10\].yc/lout[0]
+ blk.column\[9\].row\[10\].yc/lout[1] blk.column\[9\].row\[10\].yc/lin[0] blk.column\[9\].row\[10\].yc/lin[1]
+ blk.column\[10\].row\[9\].yc/vempty2 blk.column\[10\].row\[9\].yc/dout[0] blk.column\[10\].row\[9\].yc/dout[1]
+ blk.column\[10\].row\[9\].yc/din[0] blk.column\[10\].row\[9\].yc/din[1] blk.column\[10\].row\[9\].yc/dempty
+ blk.column\[10\].row\[11\].yc/uempty VPWR VGND ycell
XPHY_10908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_478_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_294_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_746_ wb_clk_i _423_/X VGND VGND VPWR VPWR wbs_dat_o[2] sky130_fd_sc_hd__dfxtp_4
XPHY_6783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_677_ VGND VGND VPWR VPWR _677_/HI la_data_out[61] sky130_fd_sc_hd__conb_1
XFILLER_1_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_520_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_486_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_490_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_488_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[7\].yc blk.column\[11\].row\[7\].yc/cbitin blk.column\[11\].row\[8\].yc/cbitin
+ blk.column\[11\].row\[7\].yc/confclk blk.column\[11\].row\[8\].yc/confclk blk.column\[11\].row\[7\].yc/dempty
+ blk.column\[11\].row\[7\].yc/din[0] blk.column\[11\].row\[7\].yc/din[1] blk.column\[11\].row\[8\].yc/uin[0]
+ blk.column\[11\].row\[8\].yc/uin[1] blk.column\[11\].row\[7\].yc/hempty blk.column\[10\].row\[7\].yc/lempty
+ blk.column\[11\].row\[7\].yc/lempty blk.column\[11\].row\[7\].yc/lin[0] blk.column\[11\].row\[7\].yc/lin[1]
+ blk.column\[12\].row\[7\].yc/rin[0] blk.column\[12\].row\[7\].yc/rin[1] blk.column\[10\].row\[7\].yc/hempty
+ blk.column\[11\].row\[7\].yc/reset blk.column\[11\].row\[8\].yc/reset blk.column\[11\].row\[7\].yc/rin[0]
+ blk.column\[11\].row\[7\].yc/rin[1] blk.column\[10\].row\[7\].yc/lin[0] blk.column\[10\].row\[7\].yc/lin[1]
+ blk.column\[11\].row\[7\].yc/uempty blk.column\[11\].row\[7\].yc/uin[0] blk.column\[11\].row\[7\].yc/uin[1]
+ blk.column\[11\].row\[6\].yc/din[0] blk.column\[11\].row\[6\].yc/din[1] blk.column\[11\].row\[6\].yc/dempty
+ blk.column\[11\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_397_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_538_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_513_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_334_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[8\].yc blk.column\[2\].row\[8\].yc/cbitin blk.column\[2\].row\[9\].yc/cbitin
+ blk.column\[2\].row\[8\].yc/confclk blk.column\[2\].row\[9\].yc/confclk blk.column\[2\].row\[8\].yc/dempty
+ blk.column\[2\].row\[8\].yc/din[0] blk.column\[2\].row\[8\].yc/din[1] blk.column\[2\].row\[9\].yc/uin[0]
+ blk.column\[2\].row\[9\].yc/uin[1] blk.column\[2\].row\[8\].yc/hempty blk.column\[1\].row\[8\].yc/lempty
+ blk.column\[2\].row\[8\].yc/lempty blk.column\[2\].row\[8\].yc/lin[0] blk.column\[2\].row\[8\].yc/lin[1]
+ blk.column\[3\].row\[8\].yc/rin[0] blk.column\[3\].row\[8\].yc/rin[1] blk.column\[1\].row\[8\].yc/hempty
+ blk.column\[2\].row\[8\].yc/reset blk.column\[2\].row\[9\].yc/reset blk.column\[2\].row\[8\].yc/rin[0]
+ blk.column\[2\].row\[8\].yc/rin[1] blk.column\[1\].row\[8\].yc/lin[0] blk.column\[1\].row\[8\].yc/lin[1]
+ blk.column\[2\].row\[8\].yc/uempty blk.column\[2\].row\[8\].yc/uin[0] blk.column\[2\].row\[8\].yc/uin[1]
+ blk.column\[2\].row\[7\].yc/din[0] blk.column\[2\].row\[7\].yc/din[1] blk.column\[2\].row\[7\].yc/dempty
+ blk.column\[2\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_330_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_497_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[11\].yc blk.column\[7\].row\[11\].yc/cbitin blk.column\[7\].row\[12\].yc/cbitin
+ blk.column\[7\].row\[11\].yc/confclk blk.column\[7\].row\[12\].yc/confclk blk.column\[7\].row\[11\].yc/dempty
+ blk.column\[7\].row\[11\].yc/din[0] blk.column\[7\].row\[11\].yc/din[1] blk.column\[7\].row\[12\].yc/uin[0]
+ blk.column\[7\].row\[12\].yc/uin[1] blk.column\[7\].row\[11\].yc/hempty blk.column\[6\].row\[11\].yc/lempty
+ blk.column\[7\].row\[11\].yc/lempty blk.column\[7\].row\[11\].yc/lin[0] blk.column\[7\].row\[11\].yc/lin[1]
+ blk.column\[8\].row\[11\].yc/rin[0] blk.column\[8\].row\[11\].yc/rin[1] blk.column\[6\].row\[11\].yc/hempty
+ blk.column\[7\].row\[11\].yc/reset blk.column\[7\].row\[12\].yc/reset blk.column\[7\].row\[11\].yc/rin[0]
+ blk.column\[7\].row\[11\].yc/rin[1] blk.column\[6\].row\[11\].yc/lin[0] blk.column\[6\].row\[11\].yc/lin[1]
+ blk.column\[7\].row\[11\].yc/uempty blk.column\[7\].row\[11\].yc/uin[0] blk.column\[7\].row\[11\].yc/uin[1]
+ blk.column\[7\].row\[10\].yc/din[0] blk.column\[7\].row\[10\].yc/din[1] blk.column\[7\].row\[10\].yc/dempty
+ blk.column\[7\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_600_ VGND VGND VPWR VPWR _600_/HI io_oeb[12] sky130_fd_sc_hd__conb_1
XFILLER_480_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_531_ VGND VGND VPWR VPWR _531_/HI _531_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_378_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_462_ VGND VGND VPWR VPWR _462_/HI _462_/LO sky130_fd_sc_hd__conb_1
XPHY_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_359_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_393_ _391_/X wbs_dat_o[24] _776_/Q _389_/X VGND VGND VPWR VPWR _768_/D sky130_fd_sc_hd__o22a_4
XPHY_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_300_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_504_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_526_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_729_ VGND VGND VPWR VPWR _729_/HI la_data_out[113] sky130_fd_sc_hd__conb_1
XFILLER_500_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_406_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_520_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xblk.column\[7\].row\[2\].yc blk.column\[7\].row\[2\].yc/cbitin blk.column\[7\].row\[3\].yc/cbitin
+ blk.column\[7\].row\[2\].yc/confclk blk.column\[7\].row\[3\].yc/confclk blk.column\[7\].row\[2\].yc/dempty
+ blk.column\[7\].row\[2\].yc/din[0] blk.column\[7\].row\[2\].yc/din[1] blk.column\[7\].row\[3\].yc/uin[0]
+ blk.column\[7\].row\[3\].yc/uin[1] blk.column\[7\].row\[2\].yc/hempty blk.column\[6\].row\[2\].yc/lempty
+ blk.column\[7\].row\[2\].yc/lempty blk.column\[7\].row\[2\].yc/lin[0] blk.column\[7\].row\[2\].yc/lin[1]
+ blk.column\[8\].row\[2\].yc/rin[0] blk.column\[8\].row\[2\].yc/rin[1] blk.column\[6\].row\[2\].yc/hempty
+ blk.column\[7\].row\[2\].yc/reset blk.column\[7\].row\[3\].yc/reset blk.column\[7\].row\[2\].yc/rin[0]
+ blk.column\[7\].row\[2\].yc/rin[1] blk.column\[6\].row\[2\].yc/lin[0] blk.column\[6\].row\[2\].yc/lin[1]
+ blk.column\[7\].row\[2\].yc/uempty blk.column\[7\].row\[2\].yc/uin[0] blk.column\[7\].row\[2\].yc/uin[1]
+ blk.column\[7\].row\[1\].yc/din[0] blk.column\[7\].row\[1\].yc/din[1] blk.column\[7\].row\[1\].yc/dempty
+ blk.column\[7\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_325_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_440_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_383_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_412_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_284_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_514_ VGND VGND VPWR VPWR _514_/HI _514_/LO sky130_fd_sc_hd__conb_1
XPHY_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_325_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_445_ VGND VGND VPWR VPWR _445_/HI _445_/LO sky130_fd_sc_hd__conb_1
XFILLER_387_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_376_ _375_/Y _373_/X wbs_dat_i[25] _373_/X VGND VGND VPWR VPWR _777_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[13\].yc blk.column\[14\].row\[13\].yc/cbitin blk.column\[14\].row\[14\].yc/cbitin
+ blk.column\[14\].row\[13\].yc/confclk blk.column\[14\].row\[14\].yc/confclk blk.column\[14\].row\[13\].yc/dempty
+ blk.column\[14\].row\[13\].yc/din[0] blk.column\[14\].row\[13\].yc/din[1] blk.column\[14\].row\[14\].yc/uin[0]
+ blk.column\[14\].row\[14\].yc/uin[1] blk.column\[14\].row\[13\].yc/hempty blk.column\[13\].row\[13\].yc/lempty
+ blk.column\[14\].row\[13\].yc/lempty blk.column\[14\].row\[13\].yc/lin[0] blk.column\[14\].row\[13\].yc/lin[1]
+ blk.column\[15\].row\[13\].yc/rin[0] blk.column\[15\].row\[13\].yc/rin[1] blk.column\[13\].row\[13\].yc/hempty
+ blk.column\[14\].row\[13\].yc/reset blk.column\[14\].row\[14\].yc/reset blk.column\[14\].row\[13\].yc/rin[0]
+ blk.column\[14\].row\[13\].yc/rin[1] blk.column\[13\].row\[13\].yc/lin[0] blk.column\[13\].row\[13\].yc/lin[1]
+ blk.column\[14\].row\[13\].yc/uempty blk.column\[14\].row\[13\].yc/uin[0] blk.column\[14\].row\[13\].yc/uin[1]
+ blk.column\[14\].row\[12\].yc/din[0] blk.column\[14\].row\[12\].yc/din[1] blk.column\[14\].row\[12\].yc/dempty
+ blk.column\[14\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_506_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_486_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_459_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_375_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_379_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_428_ VGND VGND VPWR VPWR _428_/HI _428_/LO sky130_fd_sc_hd__conb_1
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_359_ _295_/Y wbs_we_i wbs_sel_i[3] VGND VGND VPWR VPWR _359_/X sky130_fd_sc_hd__and3_4
XFILLER_536_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_493_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_530_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[9\].yc blk.column\[12\].row\[9\].yc/cbitin blk.column\[12\].row\[9\].yc/cbitout
+ blk.column\[12\].row\[9\].yc/confclk blk.column\[12\].row\[9\].yc/confclko blk.column\[12\].row\[9\].yc/dempty
+ blk.column\[12\].row\[9\].yc/din[0] blk.column\[12\].row\[9\].yc/din[1] blk.column\[12\].row\[9\].yc/dout[0]
+ blk.column\[12\].row\[9\].yc/dout[1] blk.column\[12\].row\[9\].yc/hempty blk.column\[11\].row\[9\].yc/lempty
+ blk.column\[12\].row\[9\].yc/lempty blk.column\[12\].row\[9\].yc/lin[0] blk.column\[12\].row\[9\].yc/lin[1]
+ blk.column\[13\].row\[9\].yc/rin[0] blk.column\[13\].row\[9\].yc/rin[1] blk.column\[11\].row\[9\].yc/hempty
+ blk.column\[12\].row\[9\].yc/reset blk.column\[12\].row\[9\].yc/reseto blk.column\[12\].row\[9\].yc/rin[0]
+ blk.column\[12\].row\[9\].yc/rin[1] blk.column\[11\].row\[9\].yc/lin[0] blk.column\[11\].row\[9\].yc/lin[1]
+ blk.column\[12\].row\[9\].yc/uempty blk.column\[12\].row\[9\].yc/uin[0] blk.column\[12\].row\[9\].yc/uin[1]
+ blk.column\[12\].row\[8\].yc/din[0] blk.column\[12\].row\[8\].yc/din[1] blk.column\[12\].row\[8\].yc/dempty
+ blk.column\[12\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_9_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_541_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_498_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_539_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_315_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_491_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_524_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_255_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_242_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_422_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_373_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_418_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_234_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_487_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[4\].yc blk.column\[8\].row\[4\].yc/cbitin blk.column\[8\].row\[5\].yc/cbitin
+ blk.column\[8\].row\[4\].yc/confclk blk.column\[8\].row\[5\].yc/confclk blk.column\[8\].row\[4\].yc/dempty
+ blk.column\[8\].row\[4\].yc/din[0] blk.column\[8\].row\[4\].yc/din[1] blk.column\[8\].row\[5\].yc/uin[0]
+ blk.column\[8\].row\[5\].yc/uin[1] blk.column\[8\].row\[4\].yc/hempty blk.column\[7\].row\[4\].yc/lempty
+ blk.column\[8\].row\[4\].yc/lempty blk.column\[8\].row\[4\].yc/lin[0] blk.column\[8\].row\[4\].yc/lin[1]
+ blk.column\[9\].row\[4\].yc/rin[0] blk.column\[9\].row\[4\].yc/rin[1] blk.column\[7\].row\[4\].yc/hempty
+ blk.column\[8\].row\[4\].yc/reset blk.column\[8\].row\[5\].yc/reset blk.column\[8\].row\[4\].yc/rin[0]
+ blk.column\[8\].row\[4\].yc/rin[1] blk.column\[7\].row\[4\].yc/lin[0] blk.column\[7\].row\[4\].yc/lin[1]
+ blk.column\[8\].row\[4\].yc/uempty blk.column\[8\].row\[4\].yc/uin[0] blk.column\[8\].row\[4\].yc/uin[1]
+ blk.column\[8\].row\[3\].yc/din[0] blk.column\[8\].row\[3\].yc/din[1] blk.column\[8\].row\[3\].yc/dempty
+ blk.column\[8\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_525_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_484_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_243_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_498_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_358_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_539_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_516_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[12\].yc blk.column\[2\].row\[12\].yc/cbitin blk.column\[2\].row\[13\].yc/cbitin
+ blk.column\[2\].row\[12\].yc/confclk blk.column\[2\].row\[13\].yc/confclk blk.column\[2\].row\[12\].yc/dempty
+ blk.column\[2\].row\[12\].yc/din[0] blk.column\[2\].row\[12\].yc/din[1] blk.column\[2\].row\[13\].yc/uin[0]
+ blk.column\[2\].row\[13\].yc/uin[1] blk.column\[2\].row\[12\].yc/hempty blk.column\[1\].row\[12\].yc/lempty
+ blk.column\[2\].row\[12\].yc/lempty blk.column\[2\].row\[12\].yc/lin[0] blk.column\[2\].row\[12\].yc/lin[1]
+ blk.column\[3\].row\[12\].yc/rin[0] blk.column\[3\].row\[12\].yc/rin[1] blk.column\[1\].row\[12\].yc/hempty
+ blk.column\[2\].row\[12\].yc/reset blk.column\[2\].row\[13\].yc/reset blk.column\[2\].row\[12\].yc/rin[0]
+ blk.column\[2\].row\[12\].yc/rin[1] blk.column\[1\].row\[12\].yc/lin[0] blk.column\[1\].row\[12\].yc/lin[1]
+ blk.column\[2\].row\[12\].yc/uempty blk.column\[2\].row\[12\].yc/uin[0] blk.column\[2\].row\[12\].yc/uin[1]
+ blk.column\[2\].row\[11\].yc/din[0] blk.column\[2\].row\[11\].yc/din[1] blk.column\[2\].row\[11\].yc/dempty
+ blk.column\[2\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_296_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_513_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_762_ wb_clk_i _762_/D VGND VGND VPWR VPWR wbs_dat_o[18] sky130_fd_sc_hd__dfxtp_4
XPHY_7677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_372_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_507_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_693_ VGND VGND VPWR VPWR _693_/HI la_data_out[77] sky130_fd_sc_hd__conb_1
XFILLER_5_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_451_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_531_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_372_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_332_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_269_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_474_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_293_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_409_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_503_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_356_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_489_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_484_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_462_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_541_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_314_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_745_ wb_clk_i _745_/D VGND VGND VPWR VPWR wbs_dat_o[1] sky130_fd_sc_hd__dfxtp_4
XFILLER_208_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_676_ VGND VGND VPWR VPWR _676_/HI la_data_out[60] sky130_fd_sc_hd__conb_1
XFILLER_542_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_539_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_294_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_316_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_381_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_526_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_541_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_438_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_453_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_530_ VGND VGND VPWR VPWR _530_/HI _530_/LO sky130_fd_sc_hd__conb_1
XFILLER_272_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_461_ VGND VGND VPWR VPWR _461_/HI _461_/LO sky130_fd_sc_hd__conb_1
XFILLER_521_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_376_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_392_ _391_/X wbs_dat_o[25] _375_/A _389_/X VGND VGND VPWR VPWR _769_/D sky130_fd_sc_hd__o22a_4
XPHY_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_386_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_319_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_310_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_485_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_541_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_526_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_728_ VGND VGND VPWR VPWR _728_/HI la_data_out[112] sky130_fd_sc_hd__conb_1
XFILLER_127_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_326_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_659_ VGND VGND VPWR VPWR _659_/HI io_out[33] sky130_fd_sc_hd__conb_1
XFILLER_281_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[6\].yc blk.column\[9\].row\[6\].yc/cbitin blk.column\[9\].row\[7\].yc/cbitin
+ blk.column\[9\].row\[6\].yc/confclk blk.column\[9\].row\[7\].yc/confclk blk.column\[9\].row\[6\].yc/dempty
+ blk.column\[9\].row\[6\].yc/din[0] blk.column\[9\].row\[6\].yc/din[1] blk.column\[9\].row\[7\].yc/uin[0]
+ blk.column\[9\].row\[7\].yc/uin[1] blk.column\[9\].row\[6\].yc/hempty blk.column\[8\].row\[6\].yc/lempty
+ blk.column\[9\].row\[6\].yc/lempty blk.column\[9\].row\[6\].yc/lin[0] blk.column\[9\].row\[6\].yc/lin[1]
+ blk.column\[9\].row\[6\].yc/lout[0] blk.column\[9\].row\[6\].yc/lout[1] blk.column\[8\].row\[6\].yc/hempty
+ blk.column\[9\].row\[6\].yc/reset blk.column\[9\].row\[7\].yc/reset blk.column\[9\].row\[6\].yc/rin[0]
+ blk.column\[9\].row\[6\].yc/rin[1] blk.column\[8\].row\[6\].yc/lin[0] blk.column\[8\].row\[6\].yc/lin[1]
+ blk.column\[9\].row\[6\].yc/uempty blk.column\[9\].row\[6\].yc/uin[0] blk.column\[9\].row\[6\].yc/uin[1]
+ blk.column\[9\].row\[5\].yc/din[0] blk.column\[9\].row\[5\].yc/din[1] blk.column\[9\].row\[5\].yc/dempty
+ blk.column\[9\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_457_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[15\].yc blk.column\[6\].row\[15\].yc/cbitin la_data_out[38]
+ blk.column\[6\].row\[15\].yc/confclk blk.column\[6\].row\[15\].yc/confclko _472_/HI
+ _577_/LO _578_/LO blk.column\[6\].row\[15\].yc/dout[0] blk.column\[6\].row\[15\].yc/dout[1]
+ blk.column\[6\].row\[15\].yc/hempty blk.column\[5\].row\[15\].yc/lempty blk.column\[6\].row\[15\].yc/lempty
+ blk.column\[6\].row\[15\].yc/lin[0] blk.column\[6\].row\[15\].yc/lin[1] blk.column\[7\].row\[15\].yc/rin[0]
+ blk.column\[7\].row\[15\].yc/rin[1] blk.column\[5\].row\[15\].yc/hempty blk.column\[6\].row\[15\].yc/reset
+ blk.column\[6\].row\[15\].yc/reseto blk.column\[6\].row\[15\].yc/rin[0] blk.column\[6\].row\[15\].yc/rin[1]
+ blk.column\[5\].row\[15\].yc/lin[0] blk.column\[5\].row\[15\].yc/lin[1] blk.column\[6\].row\[15\].yc/uempty
+ blk.column\[6\].row\[15\].yc/uin[0] blk.column\[6\].row\[15\].yc/uin[1] blk.column\[6\].row\[14\].yc/din[0]
+ blk.column\[6\].row\[14\].yc/din[1] blk.column\[6\].row\[14\].yc/dempty blk.column\[6\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_487_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_491_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_368_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_411_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_538_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_277_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_438_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_513_ VGND VGND VPWR VPWR _513_/HI _513_/LO sky130_fd_sc_hd__conb_1
XPHY_5176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_444_ VGND VGND VPWR VPWR _444_/HI _444_/LO sky130_fd_sc_hd__conb_1
XFILLER_260_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_375_ _375_/A VGND VGND VPWR VPWR _375_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_517_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_387_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_506_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_488_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_459_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_355_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_218_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_527_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_508_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_379_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_427_ _391_/A wbs_stb_i wbs_cyc_i _426_/Y VGND VGND VPWR VPWR _808_/D sky130_fd_sc_hd__and4_4
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_394_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_358_ _358_/A VGND VGND VPWR VPWR _358_/Y sky130_fd_sc_hd__inv_2
XFILLER_534_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_533_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_541_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_385_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_317_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_415_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_273_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[10\].yc blk.column\[8\].row\[9\].yc/cbitout blk.column\[8\].row\[11\].yc/cbitin
+ blk.column\[8\].row\[9\].yc/confclko blk.column\[8\].row\[11\].yc/confclk blk.column\[8\].row\[10\].yc/dempty
+ blk.column\[8\].row\[10\].yc/din[0] blk.column\[8\].row\[10\].yc/din[1] blk.column\[8\].row\[11\].yc/uin[0]
+ blk.column\[8\].row\[11\].yc/uin[1] blk.column\[8\].row\[10\].yc/hempty blk.column\[7\].row\[10\].yc/lempty
+ blk.column\[8\].row\[10\].yc/lempty blk.column\[8\].row\[10\].yc/lin[0] blk.column\[8\].row\[10\].yc/lin[1]
+ blk.column\[9\].row\[10\].yc/rin[0] blk.column\[9\].row\[10\].yc/rin[1] blk.column\[7\].row\[10\].yc/hempty
+ blk.column\[8\].row\[9\].yc/reseto blk.column\[8\].row\[11\].yc/reset blk.column\[8\].row\[10\].yc/rin[0]
+ blk.column\[8\].row\[10\].yc/rin[1] blk.column\[7\].row\[10\].yc/lin[0] blk.column\[7\].row\[10\].yc/lin[1]
+ blk.column\[8\].row\[9\].yc/vempty2 blk.column\[8\].row\[9\].yc/dout[0] blk.column\[8\].row\[9\].yc/dout[1]
+ blk.column\[8\].row\[9\].yc/din[0] blk.column\[8\].row\[9\].yc/din[1] blk.column\[8\].row\[9\].yc/dempty
+ blk.column\[8\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_234_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_534_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_525_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_358_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_532_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_434_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_761_ wb_clk_i _761_/D VGND VGND VPWR VPWR wbs_dat_o[17] sky130_fd_sc_hd__dfxtp_4
XFILLER_524_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_692_ VGND VGND VPWR VPWR _692_/HI la_data_out[76] sky130_fd_sc_hd__conb_1
XPHY_6977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[7\].yc blk.column\[0\].row\[7\].yc/cbitin blk.column\[0\].row\[8\].yc/cbitin
+ blk.column\[0\].row\[7\].yc/confclk blk.column\[0\].row\[8\].yc/confclk blk.column\[0\].row\[7\].yc/dempty
+ blk.column\[0\].row\[7\].yc/din[0] blk.column\[0\].row\[7\].yc/din[1] blk.column\[0\].row\[8\].yc/uin[0]
+ blk.column\[0\].row\[8\].yc/uin[1] blk.column\[0\].row\[7\].yc/hempty blk.column\[0\].row\[7\].yc/hempty2
+ blk.column\[0\].row\[7\].yc/lempty blk.column\[0\].row\[7\].yc/lin[0] blk.column\[0\].row\[7\].yc/lin[1]
+ blk.column\[1\].row\[7\].yc/rin[0] blk.column\[1\].row\[7\].yc/rin[1] _442_/HI blk.column\[0\].row\[7\].yc/reset
+ blk.column\[0\].row\[8\].yc/reset _505_/LO _506_/LO blk.column\[0\].row\[7\].yc/rout[0]
+ blk.column\[0\].row\[7\].yc/rout[1] blk.column\[0\].row\[7\].yc/uempty blk.column\[0\].row\[7\].yc/uin[0]
+ blk.column\[0\].row\[7\].yc/uin[1] blk.column\[0\].row\[6\].yc/din[0] blk.column\[0\].row\[6\].yc/din[1]
+ blk.column\[0\].row\[6\].yc/dempty blk.column\[0\].row\[8\].yc/uempty VPWR VGND
+ ycell
XFILLER_524_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_520_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_532_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_459_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_455_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_531_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_390_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_486_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_529_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_264_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_495_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_536_2268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_536_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_490_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_530_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[0\].yc la_data_in[110] blk.column\[14\].row\[1\].yc/cbitin
+ la_data_in[112] blk.column\[14\].row\[1\].yc/confclk blk.column\[14\].row\[0\].yc/dempty
+ blk.column\[14\].row\[0\].yc/din[0] blk.column\[14\].row\[0\].yc/din[1] blk.column\[14\].row\[1\].yc/uin[0]
+ blk.column\[14\].row\[1\].yc/uin[1] blk.column\[14\].row\[0\].yc/hempty blk.column\[13\].row\[0\].yc/lempty
+ blk.column\[14\].row\[0\].yc/lempty blk.column\[14\].row\[0\].yc/lin[0] blk.column\[14\].row\[0\].yc/lin[1]
+ blk.column\[15\].row\[0\].yc/rin[0] blk.column\[15\].row\[0\].yc/rin[1] blk.column\[13\].row\[0\].yc/hempty
+ la_data_in[113] blk.column\[14\].row\[1\].yc/reset blk.column\[14\].row\[0\].yc/rin[0]
+ blk.column\[14\].row\[0\].yc/rin[1] blk.column\[13\].row\[0\].yc/lin[0] blk.column\[13\].row\[0\].yc/lin[1]
+ _523_/LO la_data_in[92] la_data_in[93] la_data_out[28] la_data_out[29] blk.column\[14\].row\[0\].yc/vempty
+ blk.column\[14\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_276_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_367_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[15\].row\[12\].yc blk.column\[15\].row\[12\].yc/cbitin blk.column\[15\].row\[13\].yc/cbitin
+ blk.column\[15\].row\[12\].yc/confclk blk.column\[15\].row\[13\].yc/confclk blk.column\[15\].row\[12\].yc/dempty
+ blk.column\[15\].row\[12\].yc/din[0] blk.column\[15\].row\[12\].yc/din[1] blk.column\[15\].row\[13\].yc/uin[0]
+ blk.column\[15\].row\[13\].yc/uin[1] blk.column\[15\].row\[12\].yc/hempty blk.column\[14\].row\[12\].yc/lempty
+ _453_/HI _533_/LO _534_/LO blk.column\[15\].row\[12\].yc/lout[0] blk.column\[15\].row\[12\].yc/lout[1]
+ blk.column\[14\].row\[12\].yc/hempty blk.column\[15\].row\[12\].yc/reset blk.column\[15\].row\[13\].yc/reset
+ blk.column\[15\].row\[12\].yc/rin[0] blk.column\[15\].row\[12\].yc/rin[1] blk.column\[14\].row\[12\].yc/lin[0]
+ blk.column\[14\].row\[12\].yc/lin[1] blk.column\[15\].row\[12\].yc/uempty blk.column\[15\].row\[12\].yc/uin[0]
+ blk.column\[15\].row\[12\].yc/uin[1] blk.column\[15\].row\[11\].yc/din[0] blk.column\[15\].row\[11\].yc/din[1]
+ blk.column\[15\].row\[11\].yc/dempty blk.column\[15\].row\[13\].yc/uempty VPWR VGND
+ ycell
XFILLER_6_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_382_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_224_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_423_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_496_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[1\].yc blk.column\[5\].row\[1\].yc/cbitin blk.column\[5\].row\[2\].yc/cbitin
+ blk.column\[5\].row\[1\].yc/confclk blk.column\[5\].row\[2\].yc/confclk blk.column\[5\].row\[1\].yc/dempty
+ blk.column\[5\].row\[1\].yc/din[0] blk.column\[5\].row\[1\].yc/din[1] blk.column\[5\].row\[2\].yc/uin[0]
+ blk.column\[5\].row\[2\].yc/uin[1] blk.column\[5\].row\[1\].yc/hempty blk.column\[4\].row\[1\].yc/lempty
+ blk.column\[5\].row\[1\].yc/lempty blk.column\[5\].row\[1\].yc/lin[0] blk.column\[5\].row\[1\].yc/lin[1]
+ blk.column\[6\].row\[1\].yc/rin[0] blk.column\[6\].row\[1\].yc/rin[1] blk.column\[4\].row\[1\].yc/hempty
+ blk.column\[5\].row\[1\].yc/reset blk.column\[5\].row\[2\].yc/reset blk.column\[5\].row\[1\].yc/rin[0]
+ blk.column\[5\].row\[1\].yc/rin[1] blk.column\[4\].row\[1\].yc/lin[0] blk.column\[4\].row\[1\].yc/lin[1]
+ blk.column\[5\].row\[1\].yc/uempty blk.column\[5\].row\[1\].yc/uin[0] blk.column\[5\].row\[1\].yc/uin[1]
+ blk.column\[5\].row\[0\].yc/din[0] blk.column\[5\].row\[0\].yc/din[1] blk.column\[5\].row\[0\].yc/dempty
+ blk.column\[5\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_197_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_744_ wb_clk_i _425_/X VGND VGND VPWR VPWR wbs_dat_o[0] sky130_fd_sc_hd__dfxtp_4
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_675_ VGND VGND VPWR VPWR _675_/HI la_data_out[59] sky130_fd_sc_hd__conb_1
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_422_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_345_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_486_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_518_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_355_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_509_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_490_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_516_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_495_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_410_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_521_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_460_ VGND VGND VPWR VPWR _460_/HI _460_/LO sky130_fd_sc_hd__conb_1
XFILLER_128_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_391_ _391_/A VGND VGND VPWR VPWR _391_/X sky130_fd_sc_hd__buf_2
XPHY_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_376_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_259_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_469_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_727_ VGND VGND VPWR VPWR _727_/HI la_data_out[111] sky130_fd_sc_hd__conb_1
XFILLER_526_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_658_ VGND VGND VPWR VPWR _658_/HI io_out[32] sky130_fd_sc_hd__conb_1
XPHY_5881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_589_ VGND VGND VPWR VPWR _589_/HI io_oeb[1] sky130_fd_sc_hd__conb_1
XFILLER_504_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_353_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_392_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_481_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_401_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_411_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xblk.column\[10\].row\[8\].yc blk.column\[10\].row\[8\].yc/cbitin blk.column\[10\].row\[9\].yc/cbitin
+ blk.column\[10\].row\[8\].yc/confclk blk.column\[10\].row\[9\].yc/confclk blk.column\[10\].row\[8\].yc/dempty
+ blk.column\[10\].row\[8\].yc/din[0] blk.column\[10\].row\[8\].yc/din[1] blk.column\[10\].row\[9\].yc/uin[0]
+ blk.column\[10\].row\[9\].yc/uin[1] blk.column\[10\].row\[8\].yc/hempty blk.column\[9\].row\[8\].yc/lempty
+ blk.column\[10\].row\[8\].yc/lempty blk.column\[10\].row\[8\].yc/lin[0] blk.column\[10\].row\[8\].yc/lin[1]
+ blk.column\[11\].row\[8\].yc/rin[0] blk.column\[11\].row\[8\].yc/rin[1] blk.column\[9\].row\[8\].yc/hempty
+ blk.column\[10\].row\[8\].yc/reset blk.column\[10\].row\[9\].yc/reset blk.column\[9\].row\[8\].yc/lout[0]
+ blk.column\[9\].row\[8\].yc/lout[1] blk.column\[9\].row\[8\].yc/lin[0] blk.column\[9\].row\[8\].yc/lin[1]
+ blk.column\[10\].row\[8\].yc/uempty blk.column\[10\].row\[8\].yc/uin[0] blk.column\[10\].row\[8\].yc/uin[1]
+ blk.column\[10\].row\[7\].yc/din[0] blk.column\[10\].row\[7\].yc/din[1] blk.column\[10\].row\[7\].yc/dempty
+ blk.column\[10\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_500_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_426_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[9\].yc blk.column\[1\].row\[9\].yc/cbitin blk.column\[1\].row\[9\].yc/cbitout
+ blk.column\[1\].row\[9\].yc/confclk blk.column\[1\].row\[9\].yc/confclko blk.column\[1\].row\[9\].yc/dempty
+ blk.column\[1\].row\[9\].yc/din[0] blk.column\[1\].row\[9\].yc/din[1] blk.column\[1\].row\[9\].yc/dout[0]
+ blk.column\[1\].row\[9\].yc/dout[1] blk.column\[1\].row\[9\].yc/hempty blk.column\[0\].row\[9\].yc/lempty
+ blk.column\[1\].row\[9\].yc/lempty blk.column\[1\].row\[9\].yc/lin[0] blk.column\[1\].row\[9\].yc/lin[1]
+ blk.column\[2\].row\[9\].yc/rin[0] blk.column\[2\].row\[9\].yc/rin[1] blk.column\[0\].row\[9\].yc/hempty
+ blk.column\[1\].row\[9\].yc/reset blk.column\[1\].row\[9\].yc/reseto blk.column\[1\].row\[9\].yc/rin[0]
+ blk.column\[1\].row\[9\].yc/rin[1] blk.column\[0\].row\[9\].yc/lin[0] blk.column\[0\].row\[9\].yc/lin[1]
+ blk.column\[1\].row\[9\].yc/uempty blk.column\[1\].row\[9\].yc/uin[0] blk.column\[1\].row\[9\].yc/uin[1]
+ blk.column\[1\].row\[8\].yc/din[0] blk.column\[1\].row\[8\].yc/din[1] blk.column\[1\].row\[8\].yc/dempty
+ blk.column\[1\].row\[9\].yc/vempty2 VPWR VGND ycell
XPHY_10526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_512_ VGND VGND VPWR VPWR _512_/HI _512_/LO sky130_fd_sc_hd__conb_1
XPHY_5166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_443_ VGND VGND VPWR VPWR _443_/HI _443_/LO sky130_fd_sc_hd__conb_1
XPHY_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_374_ _372_/Y _373_/X wbs_dat_i[26] _373_/X VGND VGND VPWR VPWR _778_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[11\].yc blk.column\[3\].row\[11\].yc/cbitin blk.column\[3\].row\[12\].yc/cbitin
+ blk.column\[3\].row\[11\].yc/confclk blk.column\[3\].row\[12\].yc/confclk blk.column\[3\].row\[11\].yc/dempty
+ blk.column\[3\].row\[11\].yc/din[0] blk.column\[3\].row\[11\].yc/din[1] blk.column\[3\].row\[12\].yc/uin[0]
+ blk.column\[3\].row\[12\].yc/uin[1] blk.column\[3\].row\[11\].yc/hempty blk.column\[2\].row\[11\].yc/lempty
+ blk.column\[3\].row\[11\].yc/lempty blk.column\[3\].row\[11\].yc/lin[0] blk.column\[3\].row\[11\].yc/lin[1]
+ blk.column\[4\].row\[11\].yc/rin[0] blk.column\[4\].row\[11\].yc/rin[1] blk.column\[2\].row\[11\].yc/hempty
+ blk.column\[3\].row\[11\].yc/reset blk.column\[3\].row\[12\].yc/reset blk.column\[3\].row\[11\].yc/rin[0]
+ blk.column\[3\].row\[11\].yc/rin[1] blk.column\[2\].row\[11\].yc/lin[0] blk.column\[2\].row\[11\].yc/lin[1]
+ blk.column\[3\].row\[11\].yc/uempty blk.column\[3\].row\[11\].yc/uin[0] blk.column\[3\].row\[11\].yc/uin[1]
+ blk.column\[3\].row\[10\].yc/din[0] blk.column\[3\].row\[10\].yc/din[1] blk.column\[3\].row\[10\].yc/dempty
+ blk.column\[3\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_14_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_467_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_456_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_505_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_515_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_283_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_440_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_500_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[2\].yc blk.column\[15\].row\[2\].yc/cbitin blk.column\[15\].row\[3\].yc/cbitin
+ blk.column\[15\].row\[2\].yc/confclk blk.column\[15\].row\[3\].yc/confclk blk.column\[15\].row\[2\].yc/dempty
+ blk.column\[15\].row\[2\].yc/din[0] blk.column\[15\].row\[2\].yc/din[1] blk.column\[15\].row\[3\].yc/uin[0]
+ blk.column\[15\].row\[3\].yc/uin[1] blk.column\[15\].row\[2\].yc/hempty blk.column\[14\].row\[2\].yc/lempty
+ _459_/HI _545_/LO _546_/LO blk.column\[15\].row\[2\].yc/lout[0] blk.column\[15\].row\[2\].yc/lout[1]
+ blk.column\[14\].row\[2\].yc/hempty blk.column\[15\].row\[2\].yc/reset blk.column\[15\].row\[3\].yc/reset
+ blk.column\[15\].row\[2\].yc/rin[0] blk.column\[15\].row\[2\].yc/rin[1] blk.column\[14\].row\[2\].yc/lin[0]
+ blk.column\[14\].row\[2\].yc/lin[1] blk.column\[15\].row\[2\].yc/uempty blk.column\[15\].row\[2\].yc/uin[0]
+ blk.column\[15\].row\[2\].yc/uin[1] blk.column\[15\].row\[1\].yc/din[0] blk.column\[15\].row\[1\].yc/din[1]
+ blk.column\[15\].row\[1\].yc/dempty blk.column\[15\].row\[3\].yc/uempty VPWR VGND
+ ycell
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_219_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_524_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[3\].yc blk.column\[6\].row\[3\].yc/cbitin blk.column\[6\].row\[4\].yc/cbitin
+ blk.column\[6\].row\[3\].yc/confclk blk.column\[6\].row\[4\].yc/confclk blk.column\[6\].row\[3\].yc/dempty
+ blk.column\[6\].row\[3\].yc/din[0] blk.column\[6\].row\[3\].yc/din[1] blk.column\[6\].row\[4\].yc/uin[0]
+ blk.column\[6\].row\[4\].yc/uin[1] blk.column\[6\].row\[3\].yc/hempty blk.column\[5\].row\[3\].yc/lempty
+ blk.column\[6\].row\[3\].yc/lempty blk.column\[6\].row\[3\].yc/lin[0] blk.column\[6\].row\[3\].yc/lin[1]
+ blk.column\[7\].row\[3\].yc/rin[0] blk.column\[7\].row\[3\].yc/rin[1] blk.column\[5\].row\[3\].yc/hempty
+ blk.column\[6\].row\[3\].yc/reset blk.column\[6\].row\[4\].yc/reset blk.column\[6\].row\[3\].yc/rin[0]
+ blk.column\[6\].row\[3\].yc/rin[1] blk.column\[5\].row\[3\].yc/lin[0] blk.column\[5\].row\[3\].yc/lin[1]
+ blk.column\[6\].row\[3\].yc/uempty blk.column\[6\].row\[3\].yc/uin[0] blk.column\[6\].row\[3\].yc/uin[1]
+ blk.column\[6\].row\[2\].yc/din[0] blk.column\[6\].row\[2\].yc/din[1] blk.column\[6\].row\[2\].yc/dempty
+ blk.column\[6\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_428_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_443_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_541_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_395_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_403_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_426_ wbs_ack_o VGND VGND VPWR VPWR _426_/Y sky130_fd_sc_hd__inv_2
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_537_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ _356_/Y _352_/X wbs_dat_i[16] _339_/X VGND VGND VPWR VPWR _784_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_361_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_228_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_425_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[13\].yc blk.column\[10\].row\[13\].yc/cbitin blk.column\[10\].row\[14\].yc/cbitin
+ blk.column\[10\].row\[13\].yc/confclk blk.column\[10\].row\[14\].yc/confclk blk.column\[10\].row\[13\].yc/dempty
+ blk.column\[10\].row\[13\].yc/din[0] blk.column\[10\].row\[13\].yc/din[1] blk.column\[10\].row\[14\].yc/uin[0]
+ blk.column\[10\].row\[14\].yc/uin[1] blk.column\[10\].row\[13\].yc/hempty blk.column\[9\].row\[13\].yc/lempty
+ blk.column\[10\].row\[13\].yc/lempty blk.column\[10\].row\[13\].yc/lin[0] blk.column\[10\].row\[13\].yc/lin[1]
+ blk.column\[11\].row\[13\].yc/rin[0] blk.column\[11\].row\[13\].yc/rin[1] blk.column\[9\].row\[13\].yc/hempty
+ blk.column\[10\].row\[13\].yc/reset blk.column\[10\].row\[14\].yc/reset blk.column\[9\].row\[13\].yc/lout[0]
+ blk.column\[9\].row\[13\].yc/lout[1] blk.column\[9\].row\[13\].yc/lin[0] blk.column\[9\].row\[13\].yc/lin[1]
+ blk.column\[10\].row\[13\].yc/uempty blk.column\[10\].row\[13\].yc/uin[0] blk.column\[10\].row\[13\].yc/uin[1]
+ blk.column\[10\].row\[12\].yc/din[0] blk.column\[10\].row\[12\].yc/din[1] blk.column\[10\].row\[12\].yc/dempty
+ blk.column\[10\].row\[14\].yc/uempty VPWR VGND ycell
XPHY_9218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_361_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_369_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_317_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_472_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_310_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_453_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_529_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_464_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_542_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_409_ _405_/X wbs_dat_o[12] _326_/A _403_/X VGND VGND VPWR VPWR _756_/D sky130_fd_sc_hd__o22a_4
XFILLER_159_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_493_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_520_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_487_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_506_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[14\].yc blk.column\[7\].row\[14\].yc/cbitin blk.column\[7\].row\[15\].yc/cbitin
+ blk.column\[7\].row\[14\].yc/confclk blk.column\[7\].row\[15\].yc/confclk blk.column\[7\].row\[14\].yc/dempty
+ blk.column\[7\].row\[14\].yc/din[0] blk.column\[7\].row\[14\].yc/din[1] blk.column\[7\].row\[15\].yc/uin[0]
+ blk.column\[7\].row\[15\].yc/uin[1] blk.column\[7\].row\[14\].yc/hempty blk.column\[6\].row\[14\].yc/lempty
+ blk.column\[7\].row\[14\].yc/lempty blk.column\[7\].row\[14\].yc/lin[0] blk.column\[7\].row\[14\].yc/lin[1]
+ blk.column\[8\].row\[14\].yc/rin[0] blk.column\[8\].row\[14\].yc/rin[1] blk.column\[6\].row\[14\].yc/hempty
+ blk.column\[7\].row\[14\].yc/reset blk.column\[7\].row\[15\].yc/reset blk.column\[7\].row\[14\].yc/rin[0]
+ blk.column\[7\].row\[14\].yc/rin[1] blk.column\[6\].row\[14\].yc/lin[0] blk.column\[6\].row\[14\].yc/lin[1]
+ blk.column\[7\].row\[14\].yc/uempty blk.column\[7\].row\[14\].yc/uin[0] blk.column\[7\].row\[14\].yc/uin[1]
+ blk.column\[7\].row\[13\].yc/din[0] blk.column\[7\].row\[13\].yc/din[1] blk.column\[7\].row\[13\].yc/dempty
+ blk.column\[7\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_192_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_434_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_760_ wb_clk_i _760_/D VGND VGND VPWR VPWR wbs_dat_o[16] sky130_fd_sc_hd__dfxtp_4
XPHY_6923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_450_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_235_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_691_ VGND VGND VPWR VPWR _691_/HI la_data_out[75] sky130_fd_sc_hd__conb_1
XFILLER_101_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_305_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_455_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_531_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_475_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_351_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_344_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_462_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_483_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_245_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_507_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_503_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_510_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_529_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_363_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_513_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[5\].yc blk.column\[7\].row\[5\].yc/cbitin blk.column\[7\].row\[6\].yc/cbitin
+ blk.column\[7\].row\[5\].yc/confclk blk.column\[7\].row\[6\].yc/confclk blk.column\[7\].row\[5\].yc/dempty
+ blk.column\[7\].row\[5\].yc/din[0] blk.column\[7\].row\[5\].yc/din[1] blk.column\[7\].row\[6\].yc/uin[0]
+ blk.column\[7\].row\[6\].yc/uin[1] blk.column\[7\].row\[5\].yc/hempty blk.column\[6\].row\[5\].yc/lempty
+ blk.column\[7\].row\[5\].yc/lempty blk.column\[7\].row\[5\].yc/lin[0] blk.column\[7\].row\[5\].yc/lin[1]
+ blk.column\[8\].row\[5\].yc/rin[0] blk.column\[8\].row\[5\].yc/rin[1] blk.column\[6\].row\[5\].yc/hempty
+ blk.column\[7\].row\[5\].yc/reset blk.column\[7\].row\[6\].yc/reset blk.column\[7\].row\[5\].yc/rin[0]
+ blk.column\[7\].row\[5\].yc/rin[1] blk.column\[6\].row\[5\].yc/lin[0] blk.column\[6\].row\[5\].yc/lin[1]
+ blk.column\[7\].row\[5\].yc/uempty blk.column\[7\].row\[5\].yc/uin[0] blk.column\[7\].row\[5\].yc/uin[1]
+ blk.column\[7\].row\[4\].yc/din[0] blk.column\[7\].row\[4\].yc/din[1] blk.column\[7\].row\[4\].yc/dempty
+ blk.column\[7\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_367_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_224_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_295_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_526_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_475_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_268_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_743_ VGND VGND VPWR VPWR _743_/HI la_data_out[127] sky130_fd_sc_hd__conb_1
XPHY_7487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_674_ VGND VGND VPWR VPWR _674_/HI la_data_out[58] sky130_fd_sc_hd__conb_1
XFILLER_2_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_524_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_439_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_439_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_392_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_433_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_294_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_515_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_258_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_371_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_265_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_380_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_390_ _384_/X wbs_dat_o[26] _778_/Q _389_/X VGND VGND VPWR VPWR _770_/D sky130_fd_sc_hd__o22a_4
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_386_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_515_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_254_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_726_ VGND VGND VPWR VPWR _726_/HI la_data_out[110] sky130_fd_sc_hd__conb_1
XPHY_6572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_657_ VGND VGND VPWR VPWR _657_/HI io_out[31] sky130_fd_sc_hd__conb_1
XFILLER_483_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_588_ VGND VGND VPWR VPWR _588_/HI io_oeb[0] sky130_fd_sc_hd__conb_1
XFILLER_537_3010 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_521_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_492_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_433_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_531_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_462_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_525_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_301_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_442_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_511_ VGND VGND VPWR VPWR _511_/HI _511_/LO sky130_fd_sc_hd__conb_1
XPHY_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_442_ VGND VGND VPWR VPWR _442_/HI _442_/LO sky130_fd_sc_hd__conb_1
XPHY_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_438_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_373_ _361_/A VGND VGND VPWR VPWR _373_/X sky130_fd_sc_hd__buf_2
XFILLER_15_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_515_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_709_ VGND VGND VPWR VPWR _709_/HI la_data_out[93] sky130_fd_sc_hd__conb_1
XFILLER_541_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_480_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[7\].yc blk.column\[8\].row\[7\].yc/cbitin blk.column\[8\].row\[8\].yc/cbitin
+ blk.column\[8\].row\[7\].yc/confclk blk.column\[8\].row\[8\].yc/confclk blk.column\[8\].row\[7\].yc/dempty
+ blk.column\[8\].row\[7\].yc/din[0] blk.column\[8\].row\[7\].yc/din[1] blk.column\[8\].row\[8\].yc/uin[0]
+ blk.column\[8\].row\[8\].yc/uin[1] blk.column\[8\].row\[7\].yc/hempty blk.column\[7\].row\[7\].yc/lempty
+ blk.column\[8\].row\[7\].yc/lempty blk.column\[8\].row\[7\].yc/lin[0] blk.column\[8\].row\[7\].yc/lin[1]
+ blk.column\[9\].row\[7\].yc/rin[0] blk.column\[9\].row\[7\].yc/rin[1] blk.column\[7\].row\[7\].yc/hempty
+ blk.column\[8\].row\[7\].yc/reset blk.column\[8\].row\[8\].yc/reset blk.column\[8\].row\[7\].yc/rin[0]
+ blk.column\[8\].row\[7\].yc/rin[1] blk.column\[7\].row\[7\].yc/lin[0] blk.column\[7\].row\[7\].yc/lin[1]
+ blk.column\[8\].row\[7\].yc/uempty blk.column\[8\].row\[7\].yc/uin[0] blk.column\[8\].row\[7\].yc/uin[1]
+ blk.column\[8\].row\[6\].yc/din[0] blk.column\[8\].row\[6\].yc/din[1] blk.column\[8\].row\[6\].yc/dempty
+ blk.column\[8\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_220_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_533_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_366_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_262_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_309_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_479_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[15\].yc blk.column\[2\].row\[15\].yc/cbitin la_data_out[34]
+ blk.column\[2\].row\[15\].yc/confclk blk.column\[2\].row\[15\].yc/confclko _468_/HI
+ _565_/LO _566_/LO blk.column\[2\].row\[15\].yc/dout[0] blk.column\[2\].row\[15\].yc/dout[1]
+ blk.column\[2\].row\[15\].yc/hempty blk.column\[1\].row\[15\].yc/lempty blk.column\[2\].row\[15\].yc/lempty
+ blk.column\[2\].row\[15\].yc/lin[0] blk.column\[2\].row\[15\].yc/lin[1] blk.column\[3\].row\[15\].yc/rin[0]
+ blk.column\[3\].row\[15\].yc/rin[1] blk.column\[1\].row\[15\].yc/hempty blk.column\[2\].row\[15\].yc/reset
+ blk.column\[2\].row\[15\].yc/reseto blk.column\[2\].row\[15\].yc/rin[0] blk.column\[2\].row\[15\].yc/rin[1]
+ blk.column\[1\].row\[15\].yc/lin[0] blk.column\[1\].row\[15\].yc/lin[1] blk.column\[2\].row\[15\].yc/uempty
+ blk.column\[2\].row\[15\].yc/uin[0] blk.column\[2\].row\[15\].yc/uin[1] blk.column\[2\].row\[14\].yc/din[0]
+ blk.column\[2\].row\[14\].yc/din[1] blk.column\[2\].row\[14\].yc/dempty blk.column\[2\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_453_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_287_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_336_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_541_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_403_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_425_ _391_/A wbs_dat_o[0] _314_/A _382_/A VGND VGND VPWR VPWR _425_/X sky130_fd_sc_hd__o22a_4
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_387_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_356_ _356_/A VGND VGND VPWR VPWR _356_/Y sky130_fd_sc_hd__inv_2
XFILLER_536_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_457_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_271_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_523_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_539_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_538_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_505_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_369_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_448_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_384_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[3\].row\[0\].yc la_data_in[99] blk.column\[3\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[3\].row\[1\].yc/confclk blk.column\[3\].row\[0\].yc/dempty blk.column\[3\].row\[0\].yc/din[0]
+ blk.column\[3\].row\[0\].yc/din[1] blk.column\[3\].row\[1\].yc/uin[0] blk.column\[3\].row\[1\].yc/uin[1]
+ blk.column\[3\].row\[0\].yc/hempty blk.column\[2\].row\[0\].yc/lempty blk.column\[3\].row\[0\].yc/lempty
+ blk.column\[3\].row\[0\].yc/lin[0] blk.column\[3\].row\[0\].yc/lin[1] blk.column\[4\].row\[0\].yc/rin[0]
+ blk.column\[4\].row\[0\].yc/rin[1] blk.column\[2\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[3\].row\[1\].yc/reset blk.column\[3\].row\[0\].yc/rin[0] blk.column\[3\].row\[0\].yc/rin[1]
+ blk.column\[2\].row\[0\].yc/lin[0] blk.column\[2\].row\[0\].yc/lin[1] _567_/LO la_data_in[70]
+ la_data_in[71] la_data_out[6] la_data_out[7] blk.column\[3\].row\[0\].yc/vempty
+ blk.column\[3\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_439_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_310_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_367_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_408_ _405_/X wbs_dat_o[13] _323_/A _403_/X VGND VGND VPWR VPWR _408_/X sky130_fd_sc_hd__o22a_4
XFILLER_358_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_509_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_339_ _338_/X VGND VGND VPWR VPWR _339_/X sky130_fd_sc_hd__buf_2
XFILLER_15_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_488_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_271_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_261_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_437_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_690_ VGND VGND VPWR VPWR _690_/HI la_data_out[74] sky130_fd_sc_hd__conb_1
XPHY_6957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_507_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_531_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_351_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_475_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_515_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_491_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_486_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_368_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_507_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_482_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_442_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_483_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[9\].yc blk.column\[9\].row\[9\].yc/cbitin blk.column\[9\].row\[9\].yc/cbitout
+ blk.column\[9\].row\[9\].yc/confclk blk.column\[9\].row\[9\].yc/confclko blk.column\[9\].row\[9\].yc/dempty
+ blk.column\[9\].row\[9\].yc/din[0] blk.column\[9\].row\[9\].yc/din[1] blk.column\[9\].row\[9\].yc/dout[0]
+ blk.column\[9\].row\[9\].yc/dout[1] blk.column\[9\].row\[9\].yc/hempty blk.column\[8\].row\[9\].yc/lempty
+ blk.column\[9\].row\[9\].yc/lempty blk.column\[9\].row\[9\].yc/lin[0] blk.column\[9\].row\[9\].yc/lin[1]
+ blk.column\[9\].row\[9\].yc/lout[0] blk.column\[9\].row\[9\].yc/lout[1] blk.column\[8\].row\[9\].yc/hempty
+ blk.column\[9\].row\[9\].yc/reset blk.column\[9\].row\[9\].yc/reseto blk.column\[9\].row\[9\].yc/rin[0]
+ blk.column\[9\].row\[9\].yc/rin[1] blk.column\[8\].row\[9\].yc/lin[0] blk.column\[8\].row\[9\].yc/lin[1]
+ blk.column\[9\].row\[9\].yc/uempty blk.column\[9\].row\[9\].yc/uin[0] blk.column\[9\].row\[9\].yc/uin[1]
+ blk.column\[9\].row\[8\].yc/din[0] blk.column\[9\].row\[8\].yc/din[1] blk.column\[9\].row\[8\].yc/dempty
+ blk.column\[9\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_253_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[10\].yc blk.column\[4\].row\[9\].yc/cbitout blk.column\[4\].row\[11\].yc/cbitin
+ blk.column\[4\].row\[9\].yc/confclko blk.column\[4\].row\[11\].yc/confclk blk.column\[4\].row\[10\].yc/dempty
+ blk.column\[4\].row\[10\].yc/din[0] blk.column\[4\].row\[10\].yc/din[1] blk.column\[4\].row\[11\].yc/uin[0]
+ blk.column\[4\].row\[11\].yc/uin[1] blk.column\[4\].row\[10\].yc/hempty blk.column\[3\].row\[10\].yc/lempty
+ blk.column\[4\].row\[10\].yc/lempty blk.column\[4\].row\[10\].yc/lin[0] blk.column\[4\].row\[10\].yc/lin[1]
+ blk.column\[5\].row\[10\].yc/rin[0] blk.column\[5\].row\[10\].yc/rin[1] blk.column\[3\].row\[10\].yc/hempty
+ blk.column\[4\].row\[9\].yc/reseto blk.column\[4\].row\[11\].yc/reset blk.column\[4\].row\[10\].yc/rin[0]
+ blk.column\[4\].row\[10\].yc/rin[1] blk.column\[3\].row\[10\].yc/lin[0] blk.column\[3\].row\[10\].yc/lin[1]
+ blk.column\[4\].row\[9\].yc/vempty2 blk.column\[4\].row\[9\].yc/dout[0] blk.column\[4\].row\[9\].yc/dout[1]
+ blk.column\[4\].row\[9\].yc/din[0] blk.column\[4\].row\[9\].yc/din[1] blk.column\[4\].row\[9\].yc/dempty
+ blk.column\[4\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_520_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_312_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_367_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_398_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_742_ VGND VGND VPWR VPWR _742_/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XPHY_7477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_2097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_524_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_673_ VGND VGND VPWR VPWR _673_/HI la_data_out[57] sky130_fd_sc_hd__conb_1
XFILLER_483_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_250_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_496_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_503_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_533_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[1\].yc blk.column\[13\].row\[1\].yc/cbitin blk.column\[13\].row\[2\].yc/cbitin
+ blk.column\[13\].row\[1\].yc/confclk blk.column\[13\].row\[2\].yc/confclk blk.column\[13\].row\[1\].yc/dempty
+ blk.column\[13\].row\[1\].yc/din[0] blk.column\[13\].row\[1\].yc/din[1] blk.column\[13\].row\[2\].yc/uin[0]
+ blk.column\[13\].row\[2\].yc/uin[1] blk.column\[13\].row\[1\].yc/hempty blk.column\[12\].row\[1\].yc/lempty
+ blk.column\[13\].row\[1\].yc/lempty blk.column\[13\].row\[1\].yc/lin[0] blk.column\[13\].row\[1\].yc/lin[1]
+ blk.column\[14\].row\[1\].yc/rin[0] blk.column\[14\].row\[1\].yc/rin[1] blk.column\[12\].row\[1\].yc/hempty
+ blk.column\[13\].row\[1\].yc/reset blk.column\[13\].row\[2\].yc/reset blk.column\[13\].row\[1\].yc/rin[0]
+ blk.column\[13\].row\[1\].yc/rin[1] blk.column\[12\].row\[1\].yc/lin[0] blk.column\[12\].row\[1\].yc/lin[1]
+ blk.column\[13\].row\[1\].yc/uempty blk.column\[13\].row\[1\].yc/uin[0] blk.column\[13\].row\[1\].yc/uin[1]
+ blk.column\[13\].row\[0\].yc/din[0] blk.column\[13\].row\[0\].yc/din[1] blk.column\[13\].row\[0\].yc/dempty
+ blk.column\[13\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_525_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_217_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_519_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[2\].yc blk.column\[4\].row\[2\].yc/cbitin blk.column\[4\].row\[3\].yc/cbitin
+ blk.column\[4\].row\[2\].yc/confclk blk.column\[4\].row\[3\].yc/confclk blk.column\[4\].row\[2\].yc/dempty
+ blk.column\[4\].row\[2\].yc/din[0] blk.column\[4\].row\[2\].yc/din[1] blk.column\[4\].row\[3\].yc/uin[0]
+ blk.column\[4\].row\[3\].yc/uin[1] blk.column\[4\].row\[2\].yc/hempty blk.column\[3\].row\[2\].yc/lempty
+ blk.column\[4\].row\[2\].yc/lempty blk.column\[4\].row\[2\].yc/lin[0] blk.column\[4\].row\[2\].yc/lin[1]
+ blk.column\[5\].row\[2\].yc/rin[0] blk.column\[5\].row\[2\].yc/rin[1] blk.column\[3\].row\[2\].yc/hempty
+ blk.column\[4\].row\[2\].yc/reset blk.column\[4\].row\[3\].yc/reset blk.column\[4\].row\[2\].yc/rin[0]
+ blk.column\[4\].row\[2\].yc/rin[1] blk.column\[3\].row\[2\].yc/lin[0] blk.column\[3\].row\[2\].yc/lin[1]
+ blk.column\[4\].row\[2\].yc/uempty blk.column\[4\].row\[2\].yc/uin[0] blk.column\[4\].row\[2\].yc/uin[1]
+ blk.column\[4\].row\[1\].yc/din[0] blk.column\[4\].row\[1\].yc/din[1] blk.column\[4\].row\[1\].yc/dempty
+ blk.column\[4\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_538_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_309_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[12\].yc blk.column\[11\].row\[12\].yc/cbitin blk.column\[11\].row\[13\].yc/cbitin
+ blk.column\[11\].row\[12\].yc/confclk blk.column\[11\].row\[13\].yc/confclk blk.column\[11\].row\[12\].yc/dempty
+ blk.column\[11\].row\[12\].yc/din[0] blk.column\[11\].row\[12\].yc/din[1] blk.column\[11\].row\[13\].yc/uin[0]
+ blk.column\[11\].row\[13\].yc/uin[1] blk.column\[11\].row\[12\].yc/hempty blk.column\[10\].row\[12\].yc/lempty
+ blk.column\[11\].row\[12\].yc/lempty blk.column\[11\].row\[12\].yc/lin[0] blk.column\[11\].row\[12\].yc/lin[1]
+ blk.column\[12\].row\[12\].yc/rin[0] blk.column\[12\].row\[12\].yc/rin[1] blk.column\[10\].row\[12\].yc/hempty
+ blk.column\[11\].row\[12\].yc/reset blk.column\[11\].row\[13\].yc/reset blk.column\[11\].row\[12\].yc/rin[0]
+ blk.column\[11\].row\[12\].yc/rin[1] blk.column\[10\].row\[12\].yc/lin[0] blk.column\[10\].row\[12\].yc/lin[1]
+ blk.column\[11\].row\[12\].yc/uempty blk.column\[11\].row\[12\].yc/uin[0] blk.column\[11\].row\[12\].yc/uin[1]
+ blk.column\[11\].row\[11\].yc/din[0] blk.column\[11\].row\[11\].yc/din[1] blk.column\[11\].row\[11\].yc/dempty
+ blk.column\[11\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_87_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_254_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_489_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_725_ VGND VGND VPWR VPWR _725_/HI la_data_out[109] sky130_fd_sc_hd__conb_1
XPHY_6562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_263_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_656_ VGND VGND VPWR VPWR _656_/HI io_out[30] sky130_fd_sc_hd__conb_1
XFILLER_480_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_587_ VGND VGND VPWR VPWR _587_/HI _587_/LO sky130_fd_sc_hd__conb_1
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_433_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_509_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_214_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_368_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_301_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_516_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_478_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_514_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_510_ VGND VGND VPWR VPWR _510_/HI _510_/LO sky130_fd_sc_hd__conb_1
XPHY_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_441_ VGND VGND VPWR VPWR _441_/HI _441_/LO sky130_fd_sc_hd__conb_1
XFILLER_497_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_402_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_372_ _778_/Q VGND VGND VPWR VPWR _372_/Y sky130_fd_sc_hd__inv_2
XPHY_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_493_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[13\].yc blk.column\[8\].row\[13\].yc/cbitin blk.column\[8\].row\[14\].yc/cbitin
+ blk.column\[8\].row\[13\].yc/confclk blk.column\[8\].row\[14\].yc/confclk blk.column\[8\].row\[13\].yc/dempty
+ blk.column\[8\].row\[13\].yc/din[0] blk.column\[8\].row\[13\].yc/din[1] blk.column\[8\].row\[14\].yc/uin[0]
+ blk.column\[8\].row\[14\].yc/uin[1] blk.column\[8\].row\[13\].yc/hempty blk.column\[7\].row\[13\].yc/lempty
+ blk.column\[8\].row\[13\].yc/lempty blk.column\[8\].row\[13\].yc/lin[0] blk.column\[8\].row\[13\].yc/lin[1]
+ blk.column\[9\].row\[13\].yc/rin[0] blk.column\[9\].row\[13\].yc/rin[1] blk.column\[7\].row\[13\].yc/hempty
+ blk.column\[8\].row\[13\].yc/reset blk.column\[8\].row\[14\].yc/reset blk.column\[8\].row\[13\].yc/rin[0]
+ blk.column\[8\].row\[13\].yc/rin[1] blk.column\[7\].row\[13\].yc/lin[0] blk.column\[7\].row\[13\].yc/lin[1]
+ blk.column\[8\].row\[13\].yc/uempty blk.column\[8\].row\[13\].yc/uin[0] blk.column\[8\].row\[13\].yc/uin[1]
+ blk.column\[8\].row\[12\].yc/din[0] blk.column\[8\].row\[12\].yc/din[1] blk.column\[8\].row\[12\].yc/dempty
+ blk.column\[8\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_13_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_708_ VGND VGND VPWR VPWR _708_/HI la_data_out[92] sky130_fd_sc_hd__conb_1
XFILLER_221_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_639_ VGND VGND VPWR VPWR _639_/HI io_out[13] sky130_fd_sc_hd__conb_1
XFILLER_526_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_377_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_511_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_505_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_503_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_527_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_287_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_382_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_407_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_424_ _419_/X wbs_dat_o[1] _312_/A _382_/A VGND VGND VPWR VPWR _745_/D sky130_fd_sc_hd__o22a_4
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _354_/Y _352_/X wbs_dat_i[17] _352_/X VGND VGND VPWR VPWR _355_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_518_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_515_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_472_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_541_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_419_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_407_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xblk.column\[14\].row\[3\].yc blk.column\[14\].row\[3\].yc/cbitin blk.column\[14\].row\[4\].yc/cbitin
+ blk.column\[14\].row\[3\].yc/confclk blk.column\[14\].row\[4\].yc/confclk blk.column\[14\].row\[3\].yc/dempty
+ blk.column\[14\].row\[3\].yc/din[0] blk.column\[14\].row\[3\].yc/din[1] blk.column\[14\].row\[4\].yc/uin[0]
+ blk.column\[14\].row\[4\].yc/uin[1] blk.column\[14\].row\[3\].yc/hempty blk.column\[13\].row\[3\].yc/lempty
+ blk.column\[14\].row\[3\].yc/lempty blk.column\[14\].row\[3\].yc/lin[0] blk.column\[14\].row\[3\].yc/lin[1]
+ blk.column\[15\].row\[3\].yc/rin[0] blk.column\[15\].row\[3\].yc/rin[1] blk.column\[13\].row\[3\].yc/hempty
+ blk.column\[14\].row\[3\].yc/reset blk.column\[14\].row\[4\].yc/reset blk.column\[14\].row\[3\].yc/rin[0]
+ blk.column\[14\].row\[3\].yc/rin[1] blk.column\[13\].row\[3\].yc/lin[0] blk.column\[13\].row\[3\].yc/lin[1]
+ blk.column\[14\].row\[3\].yc/uempty blk.column\[14\].row\[3\].yc/uin[0] blk.column\[14\].row\[3\].yc/uin[1]
+ blk.column\[14\].row\[2\].yc/din[0] blk.column\[14\].row\[2\].yc/din[1] blk.column\[14\].row\[2\].yc/dempty
+ blk.column\[14\].row\[4\].yc/uempty VPWR VGND ycell
XPHY_8508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[15\].yc blk.column\[15\].row\[15\].yc/cbitin la_data_out[47]
+ blk.column\[15\].row\[15\].yc/confclk blk.column\[15\].row\[15\].yc/confclko _456_/HI
+ _539_/LO _540_/LO blk.column\[15\].row\[15\].yc/dout[0] blk.column\[15\].row\[15\].yc/dout[1]
+ blk.column\[15\].row\[15\].yc/hempty blk.column\[14\].row\[15\].yc/lempty _457_/HI
+ _541_/LO _542_/LO blk.column\[15\].row\[15\].yc/lout[0] blk.column\[15\].row\[15\].yc/lout[1]
+ blk.column\[14\].row\[15\].yc/hempty blk.column\[15\].row\[15\].yc/reset blk.column\[15\].row\[15\].yc/reseto
+ blk.column\[15\].row\[15\].yc/rin[0] blk.column\[15\].row\[15\].yc/rin[1] blk.column\[14\].row\[15\].yc/lin[0]
+ blk.column\[14\].row\[15\].yc/lin[1] blk.column\[15\].row\[15\].yc/uempty blk.column\[15\].row\[15\].yc/uin[0]
+ blk.column\[15\].row\[15\].yc/uin[1] blk.column\[15\].row\[14\].yc/din[0] blk.column\[15\].row\[14\].yc/din[1]
+ blk.column\[15\].row\[14\].yc/dempty blk.column\[15\].row\[15\].yc/vempty2 VPWR
+ VGND ycell
XFILLER_112_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_509_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[4\].yc blk.column\[5\].row\[4\].yc/cbitin blk.column\[5\].row\[5\].yc/cbitin
+ blk.column\[5\].row\[4\].yc/confclk blk.column\[5\].row\[5\].yc/confclk blk.column\[5\].row\[4\].yc/dempty
+ blk.column\[5\].row\[4\].yc/din[0] blk.column\[5\].row\[4\].yc/din[1] blk.column\[5\].row\[5\].yc/uin[0]
+ blk.column\[5\].row\[5\].yc/uin[1] blk.column\[5\].row\[4\].yc/hempty blk.column\[4\].row\[4\].yc/lempty
+ blk.column\[5\].row\[4\].yc/lempty blk.column\[5\].row\[4\].yc/lin[0] blk.column\[5\].row\[4\].yc/lin[1]
+ blk.column\[6\].row\[4\].yc/rin[0] blk.column\[6\].row\[4\].yc/rin[1] blk.column\[4\].row\[4\].yc/hempty
+ blk.column\[5\].row\[4\].yc/reset blk.column\[5\].row\[5\].yc/reset blk.column\[5\].row\[4\].yc/rin[0]
+ blk.column\[5\].row\[4\].yc/rin[1] blk.column\[4\].row\[4\].yc/lin[0] blk.column\[4\].row\[4\].yc/lin[1]
+ blk.column\[5\].row\[4\].yc/uempty blk.column\[5\].row\[4\].yc/uin[0] blk.column\[5\].row\[4\].yc/uin[1]
+ blk.column\[5\].row\[3\].yc/din[0] blk.column\[5\].row\[3\].yc/din[1] blk.column\[5\].row\[3\].yc/dempty
+ blk.column\[5\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_215_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_527_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_317_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_486_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_454_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_489_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_520_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_407_ _405_/X wbs_dat_o[14] _321_/A _403_/X VGND VGND VPWR VPWR _758_/D sky130_fd_sc_hd__o22a_4
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_499_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_338_ _295_/Y wbs_we_i wbs_sel_i[2] VGND VGND VPWR VPWR _338_/X sky130_fd_sc_hd__and3_4
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_319_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_258_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_512_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_445_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_506_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_517_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_450_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_408_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_531_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_488_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_525_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_271_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_300_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_539_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_476_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_741_ VGND VGND VPWR VPWR _741_/HI la_data_out[125] sky130_fd_sc_hd__conb_1
XPHY_6733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_409_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_672_ VGND VGND VPWR VPWR _672_/HI la_data_out[56] sky130_fd_sc_hd__conb_1
XFILLER_21_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_379_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[14\].yc blk.column\[3\].row\[14\].yc/cbitin blk.column\[3\].row\[15\].yc/cbitin
+ blk.column\[3\].row\[14\].yc/confclk blk.column\[3\].row\[15\].yc/confclk blk.column\[3\].row\[14\].yc/dempty
+ blk.column\[3\].row\[14\].yc/din[0] blk.column\[3\].row\[14\].yc/din[1] blk.column\[3\].row\[15\].yc/uin[0]
+ blk.column\[3\].row\[15\].yc/uin[1] blk.column\[3\].row\[14\].yc/hempty blk.column\[2\].row\[14\].yc/lempty
+ blk.column\[3\].row\[14\].yc/lempty blk.column\[3\].row\[14\].yc/lin[0] blk.column\[3\].row\[14\].yc/lin[1]
+ blk.column\[4\].row\[14\].yc/rin[0] blk.column\[4\].row\[14\].yc/rin[1] blk.column\[2\].row\[14\].yc/hempty
+ blk.column\[3\].row\[14\].yc/reset blk.column\[3\].row\[15\].yc/reset blk.column\[3\].row\[14\].yc/rin[0]
+ blk.column\[3\].row\[14\].yc/rin[1] blk.column\[2\].row\[14\].yc/lin[0] blk.column\[2\].row\[14\].yc/lin[1]
+ blk.column\[3\].row\[14\].yc/uempty blk.column\[3\].row\[14\].yc/uin[0] blk.column\[3\].row\[14\].yc/uin[1]
+ blk.column\[3\].row\[13\].yc/din[0] blk.column\[3\].row\[13\].yc/din[1] blk.column\[3\].row\[13\].yc/dempty
+ blk.column\[3\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_199_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_520_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_496_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_439_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_511_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_505_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_474_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_531_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[5\].yc blk.column\[15\].row\[5\].yc/cbitin blk.column\[15\].row\[6\].yc/cbitin
+ blk.column\[15\].row\[5\].yc/confclk blk.column\[15\].row\[6\].yc/confclk blk.column\[15\].row\[5\].yc/dempty
+ blk.column\[15\].row\[5\].yc/din[0] blk.column\[15\].row\[5\].yc/din[1] blk.column\[15\].row\[6\].yc/uin[0]
+ blk.column\[15\].row\[6\].yc/uin[1] blk.column\[15\].row\[5\].yc/hempty blk.column\[14\].row\[5\].yc/lempty
+ _462_/HI _551_/LO _552_/LO blk.column\[15\].row\[5\].yc/lout[0] blk.column\[15\].row\[5\].yc/lout[1]
+ blk.column\[14\].row\[5\].yc/hempty blk.column\[15\].row\[5\].yc/reset blk.column\[15\].row\[6\].yc/reset
+ blk.column\[15\].row\[5\].yc/rin[0] blk.column\[15\].row\[5\].yc/rin[1] blk.column\[14\].row\[5\].yc/lin[0]
+ blk.column\[14\].row\[5\].yc/lin[1] blk.column\[15\].row\[5\].yc/uempty blk.column\[15\].row\[5\].yc/uin[0]
+ blk.column\[15\].row\[5\].yc/uin[1] blk.column\[15\].row\[4\].yc/din[0] blk.column\[15\].row\[4\].yc/din[1]
+ blk.column\[15\].row\[4\].yc/dempty blk.column\[15\].row\[6\].yc/uempty VPWR VGND
+ ycell
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_494_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_484_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[6\].yc blk.column\[6\].row\[6\].yc/cbitin blk.column\[6\].row\[7\].yc/cbitin
+ blk.column\[6\].row\[6\].yc/confclk blk.column\[6\].row\[7\].yc/confclk blk.column\[6\].row\[6\].yc/dempty
+ blk.column\[6\].row\[6\].yc/din[0] blk.column\[6\].row\[6\].yc/din[1] blk.column\[6\].row\[7\].yc/uin[0]
+ blk.column\[6\].row\[7\].yc/uin[1] blk.column\[6\].row\[6\].yc/hempty blk.column\[5\].row\[6\].yc/lempty
+ blk.column\[6\].row\[6\].yc/lempty blk.column\[6\].row\[6\].yc/lin[0] blk.column\[6\].row\[6\].yc/lin[1]
+ blk.column\[7\].row\[6\].yc/rin[0] blk.column\[7\].row\[6\].yc/rin[1] blk.column\[5\].row\[6\].yc/hempty
+ blk.column\[6\].row\[6\].yc/reset blk.column\[6\].row\[7\].yc/reset blk.column\[6\].row\[6\].yc/rin[0]
+ blk.column\[6\].row\[6\].yc/rin[1] blk.column\[5\].row\[6\].yc/lin[0] blk.column\[5\].row\[6\].yc/lin[1]
+ blk.column\[6\].row\[6\].yc/uempty blk.column\[6\].row\[6\].yc/uin[0] blk.column\[6\].row\[6\].yc/uin[1]
+ blk.column\[6\].row\[5\].yc/din[0] blk.column\[6\].row\[5\].yc/din[1] blk.column\[6\].row\[5\].yc/dempty
+ blk.column\[6\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_480_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_225_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_724_ VGND VGND VPWR VPWR _724_/HI la_data_out[108] sky130_fd_sc_hd__conb_1
XFILLER_79_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_655_ VGND VGND VPWR VPWR _655_/HI io_out[29] sky130_fd_sc_hd__conb_1
XPHY_5862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_242_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_586_ VGND VGND VPWR VPWR _586_/HI _586_/LO sky130_fd_sc_hd__conb_1
XFILLER_405_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_357_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_479_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_301_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_401_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_292_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_438_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_440_ VGND VGND VPWR VPWR _440_/HI _440_/LO sky130_fd_sc_hd__conb_1
XPHY_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_359_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_371_ _370_/Y _366_/X wbs_dat_i[27] _366_/X VGND VGND VPWR VPWR _779_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_402_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_475_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_352_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_707_ VGND VGND VPWR VPWR _707_/HI la_data_out[91] sky130_fd_sc_hd__conb_1
XPHY_6382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_638_ VGND VGND VPWR VPWR _638_/HI io_out[12] sky130_fd_sc_hd__conb_1
XFILLER_523_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_569_ VGND VGND VPWR VPWR _569_/HI _569_/LO sky130_fd_sc_hd__conb_1
XFILLER_539_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_435_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_286_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_416_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_481_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_479_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_503_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_527_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_513_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_386_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_527_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_527_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_402_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_423_ _419_/X wbs_dat_o[2] _802_/Q _417_/X VGND VGND VPWR VPWR _423_/X sky130_fd_sc_hd__o22a_4
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_354_ _354_/A VGND VGND VPWR VPWR _354_/Y sky130_fd_sc_hd__inv_2
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_393_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_533_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_10871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_506_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_504_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[8\].yc blk.column\[7\].row\[8\].yc/cbitin blk.column\[7\].row\[9\].yc/cbitin
+ blk.column\[7\].row\[8\].yc/confclk blk.column\[7\].row\[9\].yc/confclk blk.column\[7\].row\[8\].yc/dempty
+ blk.column\[7\].row\[8\].yc/din[0] blk.column\[7\].row\[8\].yc/din[1] blk.column\[7\].row\[9\].yc/uin[0]
+ blk.column\[7\].row\[9\].yc/uin[1] blk.column\[7\].row\[8\].yc/hempty blk.column\[6\].row\[8\].yc/lempty
+ blk.column\[7\].row\[8\].yc/lempty blk.column\[7\].row\[8\].yc/lin[0] blk.column\[7\].row\[8\].yc/lin[1]
+ blk.column\[8\].row\[8\].yc/rin[0] blk.column\[8\].row\[8\].yc/rin[1] blk.column\[6\].row\[8\].yc/hempty
+ blk.column\[7\].row\[8\].yc/reset blk.column\[7\].row\[9\].yc/reset blk.column\[7\].row\[8\].yc/rin[0]
+ blk.column\[7\].row\[8\].yc/rin[1] blk.column\[6\].row\[8\].yc/lin[0] blk.column\[6\].row\[8\].yc/lin[1]
+ blk.column\[7\].row\[8\].yc/uempty blk.column\[7\].row\[8\].yc/uin[0] blk.column\[7\].row\[8\].yc/uin[1]
+ blk.column\[7\].row\[7\].yc/din[0] blk.column\[7\].row\[7\].yc/din[1] blk.column\[7\].row\[7\].yc/dempty
+ blk.column\[7\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_533_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_524_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_483_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_227_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_418_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_448_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_507_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_395_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_278_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_406_ _405_/X wbs_dat_o[15] _316_/A _403_/X VGND VGND VPWR VPWR _406_/X sky130_fd_sc_hd__o22a_4
XFILLER_15_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_375_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_337_ _337_/A VGND VGND VPWR VPWR _337_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_390_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[11\].yc blk.column\[12\].row\[11\].yc/cbitin blk.column\[12\].row\[12\].yc/cbitin
+ blk.column\[12\].row\[11\].yc/confclk blk.column\[12\].row\[12\].yc/confclk blk.column\[12\].row\[11\].yc/dempty
+ blk.column\[12\].row\[11\].yc/din[0] blk.column\[12\].row\[11\].yc/din[1] blk.column\[12\].row\[12\].yc/uin[0]
+ blk.column\[12\].row\[12\].yc/uin[1] blk.column\[12\].row\[11\].yc/hempty blk.column\[11\].row\[11\].yc/lempty
+ blk.column\[12\].row\[11\].yc/lempty blk.column\[12\].row\[11\].yc/lin[0] blk.column\[12\].row\[11\].yc/lin[1]
+ blk.column\[13\].row\[11\].yc/rin[0] blk.column\[13\].row\[11\].yc/rin[1] blk.column\[11\].row\[11\].yc/hempty
+ blk.column\[12\].row\[11\].yc/reset blk.column\[12\].row\[12\].yc/reset blk.column\[12\].row\[11\].yc/rin[0]
+ blk.column\[12\].row\[11\].yc/rin[1] blk.column\[11\].row\[11\].yc/lin[0] blk.column\[11\].row\[11\].yc/lin[1]
+ blk.column\[12\].row\[11\].yc/uempty blk.column\[12\].row\[11\].yc/uin[0] blk.column\[12\].row\[11\].yc/uin[1]
+ blk.column\[12\].row\[10\].yc/din[0] blk.column\[12\].row\[10\].yc/din[1] blk.column\[12\].row\[10\].yc/dempty
+ blk.column\[12\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_508_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_528_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_401_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_498_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_307_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_413_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_517_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_514_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_309_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_239_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_372_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[0\].yc la_data_in[107] blk.column\[11\].row\[1\].yc/cbitin
+ la_data_in[112] blk.column\[11\].row\[1\].yc/confclk blk.column\[11\].row\[0\].yc/dempty
+ blk.column\[11\].row\[0\].yc/din[0] blk.column\[11\].row\[0\].yc/din[1] blk.column\[11\].row\[1\].yc/uin[0]
+ blk.column\[11\].row\[1\].yc/uin[1] blk.column\[11\].row\[0\].yc/hempty blk.column\[10\].row\[0\].yc/lempty
+ blk.column\[11\].row\[0\].yc/lempty blk.column\[11\].row\[0\].yc/lin[0] blk.column\[11\].row\[0\].yc/lin[1]
+ blk.column\[12\].row\[0\].yc/rin[0] blk.column\[12\].row\[0\].yc/rin[1] blk.column\[10\].row\[0\].yc/hempty
+ la_data_in[113] blk.column\[11\].row\[1\].yc/reset blk.column\[11\].row\[0\].yc/rin[0]
+ blk.column\[11\].row\[0\].yc/rin[1] blk.column\[10\].row\[0\].yc/lin[0] blk.column\[10\].row\[0\].yc/lin[1]
+ _514_/LO la_data_in[86] la_data_in[87] la_data_out[22] la_data_out[23] blk.column\[11\].row\[0\].yc/vempty
+ blk.column\[11\].row\[1\].yc/uempty VPWR VGND ycell
XPHY_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_390_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[2\].row\[1\].yc blk.column\[2\].row\[1\].yc/cbitin blk.column\[2\].row\[2\].yc/cbitin
+ blk.column\[2\].row\[1\].yc/confclk blk.column\[2\].row\[2\].yc/confclk blk.column\[2\].row\[1\].yc/dempty
+ blk.column\[2\].row\[1\].yc/din[0] blk.column\[2\].row\[1\].yc/din[1] blk.column\[2\].row\[2\].yc/uin[0]
+ blk.column\[2\].row\[2\].yc/uin[1] blk.column\[2\].row\[1\].yc/hempty blk.column\[1\].row\[1\].yc/lempty
+ blk.column\[2\].row\[1\].yc/lempty blk.column\[2\].row\[1\].yc/lin[0] blk.column\[2\].row\[1\].yc/lin[1]
+ blk.column\[3\].row\[1\].yc/rin[0] blk.column\[3\].row\[1\].yc/rin[1] blk.column\[1\].row\[1\].yc/hempty
+ blk.column\[2\].row\[1\].yc/reset blk.column\[2\].row\[2\].yc/reset blk.column\[2\].row\[1\].yc/rin[0]
+ blk.column\[2\].row\[1\].yc/rin[1] blk.column\[1\].row\[1\].yc/lin[0] blk.column\[1\].row\[1\].yc/lin[1]
+ blk.column\[2\].row\[1\].yc/uempty blk.column\[2\].row\[1\].yc/uin[0] blk.column\[2\].row\[1\].yc/uin[1]
+ blk.column\[2\].row\[0\].yc/din[0] blk.column\[2\].row\[0\].yc/din[1] blk.column\[2\].row\[0\].yc/dempty
+ blk.column\[2\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_542_3125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_409_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_427_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_395_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[9\].row\[12\].yc blk.column\[9\].row\[12\].yc/cbitin blk.column\[9\].row\[13\].yc/cbitin
+ blk.column\[9\].row\[12\].yc/confclk blk.column\[9\].row\[13\].yc/confclk blk.column\[9\].row\[12\].yc/dempty
+ blk.column\[9\].row\[12\].yc/din[0] blk.column\[9\].row\[12\].yc/din[1] blk.column\[9\].row\[13\].yc/uin[0]
+ blk.column\[9\].row\[13\].yc/uin[1] blk.column\[9\].row\[12\].yc/hempty blk.column\[8\].row\[12\].yc/lempty
+ blk.column\[9\].row\[12\].yc/lempty blk.column\[9\].row\[12\].yc/lin[0] blk.column\[9\].row\[12\].yc/lin[1]
+ blk.column\[9\].row\[12\].yc/lout[0] blk.column\[9\].row\[12\].yc/lout[1] blk.column\[8\].row\[12\].yc/hempty
+ blk.column\[9\].row\[12\].yc/reset blk.column\[9\].row\[13\].yc/reset blk.column\[9\].row\[12\].yc/rin[0]
+ blk.column\[9\].row\[12\].yc/rin[1] blk.column\[8\].row\[12\].yc/lin[0] blk.column\[8\].row\[12\].yc/lin[1]
+ blk.column\[9\].row\[12\].yc/uempty blk.column\[9\].row\[12\].yc/uin[0] blk.column\[9\].row\[12\].yc/uin[1]
+ blk.column\[9\].row\[11\].yc/din[0] blk.column\[9\].row\[11\].yc/din[1] blk.column\[9\].row\[11\].yc/dempty
+ blk.column\[9\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_238_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_436_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_477_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_492_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_334_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_244_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_270_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_443_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_420_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_541_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_510_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2033 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_244_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_740_ VGND VGND VPWR VPWR _740_/HI la_data_out[124] sky130_fd_sc_hd__conb_1
XPHY_7457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_309_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_671_ VGND VGND VPWR VPWR _671_/HI la_data_out[55] sky130_fd_sc_hd__conb_1
XPHY_6767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_523_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_478_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_490_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_439_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_433_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_316_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_345_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_474_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_470_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_542_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_503_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_506_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[10\].yc blk.column\[0\].row\[9\].yc/cbitout blk.column\[0\].row\[11\].yc/cbitin
+ blk.column\[0\].row\[9\].yc/confclko blk.column\[0\].row\[11\].yc/confclk blk.column\[0\].row\[10\].yc/dempty
+ blk.column\[0\].row\[10\].yc/din[0] blk.column\[0\].row\[10\].yc/din[1] blk.column\[0\].row\[11\].yc/uin[0]
+ blk.column\[0\].row\[11\].yc/uin[1] blk.column\[0\].row\[10\].yc/hempty blk.column\[0\].row\[10\].yc/hempty2
+ blk.column\[0\].row\[10\].yc/lempty blk.column\[0\].row\[10\].yc/lin[0] blk.column\[0\].row\[10\].yc/lin[1]
+ blk.column\[1\].row\[10\].yc/rin[0] blk.column\[1\].row\[10\].yc/rin[1] _429_/HI
+ blk.column\[0\].row\[9\].yc/reseto blk.column\[0\].row\[11\].yc/reset _479_/LO _480_/LO
+ blk.column\[0\].row\[10\].yc/rout[0] blk.column\[0\].row\[10\].yc/rout[1] blk.column\[0\].row\[9\].yc/vempty2
+ blk.column\[0\].row\[9\].yc/dout[0] blk.column\[0\].row\[9\].yc/dout[1] blk.column\[0\].row\[9\].yc/din[0]
+ blk.column\[0\].row\[9\].yc/din[1] blk.column\[0\].row\[9\].yc/dempty blk.column\[0\].row\[11\].yc/uempty
+ VPWR VGND ycell
XFILLER_484_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_406_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_228_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_508_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_341_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_519_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_532_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_473_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_723_ VGND VGND VPWR VPWR _723_/HI la_data_out[107] sky130_fd_sc_hd__conb_1
XFILLER_208_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_654_ VGND VGND VPWR VPWR _654_/HI io_out[28] sky130_fd_sc_hd__conb_1
XPHY_6586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_585_ VGND VGND VPWR VPWR _585_/HI _585_/LO sky130_fd_sc_hd__conb_1
XFILLER_261_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_537_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_484_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_481_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_507_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_479_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_440_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_520_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_309_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_522_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[12\].row\[2\].yc blk.column\[12\].row\[2\].yc/cbitin blk.column\[12\].row\[3\].yc/cbitin
+ blk.column\[12\].row\[2\].yc/confclk blk.column\[12\].row\[3\].yc/confclk blk.column\[12\].row\[2\].yc/dempty
+ blk.column\[12\].row\[2\].yc/din[0] blk.column\[12\].row\[2\].yc/din[1] blk.column\[12\].row\[3\].yc/uin[0]
+ blk.column\[12\].row\[3\].yc/uin[1] blk.column\[12\].row\[2\].yc/hempty blk.column\[11\].row\[2\].yc/lempty
+ blk.column\[12\].row\[2\].yc/lempty blk.column\[12\].row\[2\].yc/lin[0] blk.column\[12\].row\[2\].yc/lin[1]
+ blk.column\[13\].row\[2\].yc/rin[0] blk.column\[13\].row\[2\].yc/rin[1] blk.column\[11\].row\[2\].yc/hempty
+ blk.column\[12\].row\[2\].yc/reset blk.column\[12\].row\[3\].yc/reset blk.column\[12\].row\[2\].yc/rin[0]
+ blk.column\[12\].row\[2\].yc/rin[1] blk.column\[11\].row\[2\].yc/lin[0] blk.column\[11\].row\[2\].yc/lin[1]
+ blk.column\[12\].row\[2\].yc/uempty blk.column\[12\].row\[2\].yc/uin[0] blk.column\[12\].row\[2\].yc/uin[1]
+ blk.column\[12\].row\[1\].yc/din[0] blk.column\[12\].row\[1\].yc/din[1] blk.column\[12\].row\[1\].yc/dempty
+ blk.column\[12\].row\[3\].yc/uempty VPWR VGND ycell
XPHY_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_325_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_399_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_370_ _779_/Q VGND VGND VPWR VPWR _370_/Y sky130_fd_sc_hd__inv_2
XFILLER_359_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[3\].yc blk.column\[3\].row\[3\].yc/cbitin blk.column\[3\].row\[4\].yc/cbitin
+ blk.column\[3\].row\[3\].yc/confclk blk.column\[3\].row\[4\].yc/confclk blk.column\[3\].row\[3\].yc/dempty
+ blk.column\[3\].row\[3\].yc/din[0] blk.column\[3\].row\[3\].yc/din[1] blk.column\[3\].row\[4\].yc/uin[0]
+ blk.column\[3\].row\[4\].yc/uin[1] blk.column\[3\].row\[3\].yc/hempty blk.column\[2\].row\[3\].yc/lempty
+ blk.column\[3\].row\[3\].yc/lempty blk.column\[3\].row\[3\].yc/lin[0] blk.column\[3\].row\[3\].yc/lin[1]
+ blk.column\[4\].row\[3\].yc/rin[0] blk.column\[4\].row\[3\].yc/rin[1] blk.column\[2\].row\[3\].yc/hempty
+ blk.column\[3\].row\[3\].yc/reset blk.column\[3\].row\[4\].yc/reset blk.column\[3\].row\[3\].yc/rin[0]
+ blk.column\[3\].row\[3\].yc/rin[1] blk.column\[2\].row\[3\].yc/lin[0] blk.column\[2\].row\[3\].yc/lin[1]
+ blk.column\[3\].row\[3\].yc/uempty blk.column\[3\].row\[3\].yc/uin[0] blk.column\[3\].row\[3\].yc/uin[1]
+ blk.column\[3\].row\[2\].yc/din[0] blk.column\[3\].row\[2\].yc/din[1] blk.column\[3\].row\[2\].yc/dempty
+ blk.column\[3\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_512_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_706_ VGND VGND VPWR VPWR _706_/HI la_data_out[90] sky130_fd_sc_hd__conb_1
XFILLER_504_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_324_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_637_ VGND VGND VPWR VPWR _637_/HI io_out[11] sky130_fd_sc_hd__conb_1
XFILLER_480_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_568_ VGND VGND VPWR VPWR _568_/HI _568_/LO sky130_fd_sc_hd__conb_1
XPHY_4981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_499_ VGND VGND VPWR VPWR _499_/HI _499_/LO sky130_fd_sc_hd__conb_1
XFILLER_13_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_393_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_522_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_492_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_516_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_331_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_422_ _419_/X wbs_dat_o[3] _307_/A _417_/X VGND VGND VPWR VPWR _747_/D sky130_fd_sc_hd__o22a_4
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_353_ _351_/Y _352_/X wbs_dat_i[18] _352_/X VGND VGND VPWR VPWR _786_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_319_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_393_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_457_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[13\].yc blk.column\[4\].row\[13\].yc/cbitin blk.column\[4\].row\[14\].yc/cbitin
+ blk.column\[4\].row\[13\].yc/confclk blk.column\[4\].row\[14\].yc/confclk blk.column\[4\].row\[13\].yc/dempty
+ blk.column\[4\].row\[13\].yc/din[0] blk.column\[4\].row\[13\].yc/din[1] blk.column\[4\].row\[14\].yc/uin[0]
+ blk.column\[4\].row\[14\].yc/uin[1] blk.column\[4\].row\[13\].yc/hempty blk.column\[3\].row\[13\].yc/lempty
+ blk.column\[4\].row\[13\].yc/lempty blk.column\[4\].row\[13\].yc/lin[0] blk.column\[4\].row\[13\].yc/lin[1]
+ blk.column\[5\].row\[13\].yc/rin[0] blk.column\[5\].row\[13\].yc/rin[1] blk.column\[3\].row\[13\].yc/hempty
+ blk.column\[4\].row\[13\].yc/reset blk.column\[4\].row\[14\].yc/reset blk.column\[4\].row\[13\].yc/rin[0]
+ blk.column\[4\].row\[13\].yc/rin[1] blk.column\[3\].row\[13\].yc/lin[0] blk.column\[3\].row\[13\].yc/lin[1]
+ blk.column\[4\].row\[13\].yc/uempty blk.column\[4\].row\[13\].yc/uin[0] blk.column\[4\].row\[13\].yc/uin[1]
+ blk.column\[4\].row\[12\].yc/din[0] blk.column\[4\].row\[12\].yc/din[1] blk.column\[4\].row\[12\].yc/dempty
+ blk.column\[4\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_18_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_498_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_518_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_448_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_513_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_386_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_505_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ _419_/A VGND VGND VPWR VPWR _405_/X sky130_fd_sc_hd__buf_2
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_336_ _335_/Y _331_/X wbs_dat_i[8] _319_/A VGND VGND VPWR VPWR _336_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_471_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_358_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_316_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_432_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_512_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_498_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_523_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_418_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_535_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[4\].yc blk.column\[13\].row\[4\].yc/cbitin blk.column\[13\].row\[5\].yc/cbitin
+ blk.column\[13\].row\[4\].yc/confclk blk.column\[13\].row\[5\].yc/confclk blk.column\[13\].row\[4\].yc/dempty
+ blk.column\[13\].row\[4\].yc/din[0] blk.column\[13\].row\[4\].yc/din[1] blk.column\[13\].row\[5\].yc/uin[0]
+ blk.column\[13\].row\[5\].yc/uin[1] blk.column\[13\].row\[4\].yc/hempty blk.column\[12\].row\[4\].yc/lempty
+ blk.column\[13\].row\[4\].yc/lempty blk.column\[13\].row\[4\].yc/lin[0] blk.column\[13\].row\[4\].yc/lin[1]
+ blk.column\[14\].row\[4\].yc/rin[0] blk.column\[14\].row\[4\].yc/rin[1] blk.column\[12\].row\[4\].yc/hempty
+ blk.column\[13\].row\[4\].yc/reset blk.column\[13\].row\[5\].yc/reset blk.column\[13\].row\[4\].yc/rin[0]
+ blk.column\[13\].row\[4\].yc/rin[1] blk.column\[12\].row\[4\].yc/lin[0] blk.column\[12\].row\[4\].yc/lin[1]
+ blk.column\[13\].row\[4\].yc/uempty blk.column\[13\].row\[4\].yc/uin[0] blk.column\[13\].row\[4\].yc/uin[1]
+ blk.column\[13\].row\[3\].yc/din[0] blk.column\[13\].row\[3\].yc/din[1] blk.column\[13\].row\[3\].yc/dempty
+ blk.column\[13\].row\[5\].yc/uempty VPWR VGND ycell
XPHY_6905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_383_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[5\].yc blk.column\[4\].row\[5\].yc/cbitin blk.column\[4\].row\[6\].yc/cbitin
+ blk.column\[4\].row\[5\].yc/confclk blk.column\[4\].row\[6\].yc/confclk blk.column\[4\].row\[5\].yc/dempty
+ blk.column\[4\].row\[5\].yc/din[0] blk.column\[4\].row\[5\].yc/din[1] blk.column\[4\].row\[6\].yc/uin[0]
+ blk.column\[4\].row\[6\].yc/uin[1] blk.column\[4\].row\[5\].yc/hempty blk.column\[3\].row\[5\].yc/lempty
+ blk.column\[4\].row\[5\].yc/lempty blk.column\[4\].row\[5\].yc/lin[0] blk.column\[4\].row\[5\].yc/lin[1]
+ blk.column\[5\].row\[5\].yc/rin[0] blk.column\[5\].row\[5\].yc/rin[1] blk.column\[3\].row\[5\].yc/hempty
+ blk.column\[4\].row\[5\].yc/reset blk.column\[4\].row\[6\].yc/reset blk.column\[4\].row\[5\].yc/rin[0]
+ blk.column\[4\].row\[5\].yc/rin[1] blk.column\[3\].row\[5\].yc/lin[0] blk.column\[3\].row\[5\].yc/lin[1]
+ blk.column\[4\].row\[5\].yc/uempty blk.column\[4\].row\[5\].yc/uin[0] blk.column\[4\].row\[5\].yc/uin[1]
+ blk.column\[4\].row\[4\].yc/din[0] blk.column\[4\].row\[4\].yc/din[1] blk.column\[4\].row\[4\].yc/dempty
+ blk.column\[4\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_494_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xblk.column\[11\].row\[15\].yc blk.column\[11\].row\[15\].yc/cbitin la_data_out[43]
+ blk.column\[11\].row\[15\].yc/confclk blk.column\[11\].row\[15\].yc/confclko _446_/HI
+ _515_/LO _516_/LO blk.column\[11\].row\[15\].yc/dout[0] blk.column\[11\].row\[15\].yc/dout[1]
+ blk.column\[11\].row\[15\].yc/hempty blk.column\[10\].row\[15\].yc/lempty blk.column\[11\].row\[15\].yc/lempty
+ blk.column\[11\].row\[15\].yc/lin[0] blk.column\[11\].row\[15\].yc/lin[1] blk.column\[12\].row\[15\].yc/rin[0]
+ blk.column\[12\].row\[15\].yc/rin[1] blk.column\[10\].row\[15\].yc/hempty blk.column\[11\].row\[15\].yc/reset
+ blk.column\[11\].row\[15\].yc/reseto blk.column\[11\].row\[15\].yc/rin[0] blk.column\[11\].row\[15\].yc/rin[1]
+ blk.column\[10\].row\[15\].yc/lin[0] blk.column\[10\].row\[15\].yc/lin[1] blk.column\[11\].row\[15\].yc/uempty
+ blk.column\[11\].row\[15\].yc/uin[0] blk.column\[11\].row\[15\].yc/uin[1] blk.column\[11\].row\[14\].yc/din[0]
+ blk.column\[11\].row\[14\].yc/din[1] blk.column\[11\].row\[14\].yc/dempty blk.column\[11\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XPHY_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_515_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_514_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_499_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_435_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_319_ _319_/A VGND VGND VPWR VPWR _319_/X sky130_fd_sc_hd__buf_2
XFILLER_497_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_493_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_217_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_518_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_408_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_350_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_525_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_394_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_429_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_517_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_268_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_670_ VGND VGND VPWR VPWR _670_/HI la_data_out[54] sky130_fd_sc_hd__conb_1
XPHY_6757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_309_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_377_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_478_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_339_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_374_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_474_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_799_ wb_clk_i _320_/X VGND VGND VPWR VPWR _316_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_1_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_542_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_403_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_342_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_249_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_293_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_514_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_380_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_538_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_299_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_722_ VGND VGND VPWR VPWR _722_/HI la_data_out[106] sky130_fd_sc_hd__conb_1
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_653_ VGND VGND VPWR VPWR _653_/HI io_out[27] sky130_fd_sc_hd__conb_1
XPHY_6576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_584_ VGND VGND VPWR VPWR _584_/HI _584_/LO sky130_fd_sc_hd__conb_1
XPHY_5886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_358_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_508_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_534_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_516_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_433_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[10\].yc blk.column\[13\].row\[9\].yc/cbitout blk.column\[13\].row\[11\].yc/cbitin
+ blk.column\[13\].row\[9\].yc/confclko blk.column\[13\].row\[11\].yc/confclk blk.column\[13\].row\[10\].yc/dempty
+ blk.column\[13\].row\[10\].yc/din[0] blk.column\[13\].row\[10\].yc/din[1] blk.column\[13\].row\[11\].yc/uin[0]
+ blk.column\[13\].row\[11\].yc/uin[1] blk.column\[13\].row\[10\].yc/hempty blk.column\[12\].row\[10\].yc/lempty
+ blk.column\[13\].row\[10\].yc/lempty blk.column\[13\].row\[10\].yc/lin[0] blk.column\[13\].row\[10\].yc/lin[1]
+ blk.column\[14\].row\[10\].yc/rin[0] blk.column\[14\].row\[10\].yc/rin[1] blk.column\[12\].row\[10\].yc/hempty
+ blk.column\[13\].row\[9\].yc/reseto blk.column\[13\].row\[11\].yc/reset blk.column\[13\].row\[10\].yc/rin[0]
+ blk.column\[13\].row\[10\].yc/rin[1] blk.column\[12\].row\[10\].yc/lin[0] blk.column\[12\].row\[10\].yc/lin[1]
+ blk.column\[13\].row\[9\].yc/vempty2 blk.column\[13\].row\[9\].yc/dout[0] blk.column\[13\].row\[9\].yc/dout[1]
+ blk.column\[13\].row\[9\].yc/din[0] blk.column\[13\].row\[9\].yc/din[1] blk.column\[13\].row\[9\].yc/dempty
+ blk.column\[13\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_258_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_271_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[6\].yc blk.column\[14\].row\[6\].yc/cbitin blk.column\[14\].row\[7\].yc/cbitin
+ blk.column\[14\].row\[6\].yc/confclk blk.column\[14\].row\[7\].yc/confclk blk.column\[14\].row\[6\].yc/dempty
+ blk.column\[14\].row\[6\].yc/din[0] blk.column\[14\].row\[6\].yc/din[1] blk.column\[14\].row\[7\].yc/uin[0]
+ blk.column\[14\].row\[7\].yc/uin[1] blk.column\[14\].row\[6\].yc/hempty blk.column\[13\].row\[6\].yc/lempty
+ blk.column\[14\].row\[6\].yc/lempty blk.column\[14\].row\[6\].yc/lin[0] blk.column\[14\].row\[6\].yc/lin[1]
+ blk.column\[15\].row\[6\].yc/rin[0] blk.column\[15\].row\[6\].yc/rin[1] blk.column\[13\].row\[6\].yc/hempty
+ blk.column\[14\].row\[6\].yc/reset blk.column\[14\].row\[7\].yc/reset blk.column\[14\].row\[6\].yc/rin[0]
+ blk.column\[14\].row\[6\].yc/rin[1] blk.column\[13\].row\[6\].yc/lin[0] blk.column\[13\].row\[6\].yc/lin[1]
+ blk.column\[14\].row\[6\].yc/uempty blk.column\[14\].row\[6\].yc/uin[0] blk.column\[14\].row\[6\].yc/uin[1]
+ blk.column\[14\].row\[5\].yc/din[0] blk.column\[14\].row\[5\].yc/din[1] blk.column\[14\].row\[5\].yc/dempty
+ blk.column\[14\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_209_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_324_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_429_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[5\].row\[7\].yc blk.column\[5\].row\[7\].yc/cbitin blk.column\[5\].row\[8\].yc/cbitin
+ blk.column\[5\].row\[7\].yc/confclk blk.column\[5\].row\[8\].yc/confclk blk.column\[5\].row\[7\].yc/dempty
+ blk.column\[5\].row\[7\].yc/din[0] blk.column\[5\].row\[7\].yc/din[1] blk.column\[5\].row\[8\].yc/uin[0]
+ blk.column\[5\].row\[8\].yc/uin[1] blk.column\[5\].row\[7\].yc/hempty blk.column\[4\].row\[7\].yc/lempty
+ blk.column\[5\].row\[7\].yc/lempty blk.column\[5\].row\[7\].yc/lin[0] blk.column\[5\].row\[7\].yc/lin[1]
+ blk.column\[6\].row\[7\].yc/rin[0] blk.column\[6\].row\[7\].yc/rin[1] blk.column\[4\].row\[7\].yc/hempty
+ blk.column\[5\].row\[7\].yc/reset blk.column\[5\].row\[8\].yc/reset blk.column\[5\].row\[7\].yc/rin[0]
+ blk.column\[5\].row\[7\].yc/rin[1] blk.column\[4\].row\[7\].yc/lin[0] blk.column\[4\].row\[7\].yc/lin[1]
+ blk.column\[5\].row\[7\].yc/uempty blk.column\[5\].row\[7\].yc/uin[0] blk.column\[5\].row\[7\].yc/uin[1]
+ blk.column\[5\].row\[6\].yc/din[0] blk.column\[5\].row\[6\].yc/din[1] blk.column\[5\].row\[6\].yc/dempty
+ blk.column\[5\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_245_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_325_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_359_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_336_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_313_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_705_ VGND VGND VPWR VPWR _705_/HI la_data_out[89] sky130_fd_sc_hd__conb_1
XFILLER_189_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_636_ VGND VGND VPWR VPWR _636_/HI io_out[10] sky130_fd_sc_hd__conb_1
XPHY_5672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_400_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_567_ VGND VGND VPWR VPWR _567_/HI _567_/LO sky130_fd_sc_hd__conb_1
XPHY_4982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_500_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_498_ VGND VGND VPWR VPWR _498_/HI _498_/LO sky130_fd_sc_hd__conb_1
XFILLER_474_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_523_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_361_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_331_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_416_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_522_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_520_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_542_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_394_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_437_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_352_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_271_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_442_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_421_ _419_/X wbs_dat_o[4] _305_/A _417_/X VGND VGND VPWR VPWR _748_/D sky130_fd_sc_hd__o22a_4
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_352_ _339_/X VGND VGND VPWR VPWR _352_/X sky130_fd_sc_hd__buf_2
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_331_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_319_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_519_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_469_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_430_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_472_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_504_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_619_ VGND VGND VPWR VPWR _619_/HI io_oeb[31] sky130_fd_sc_hd__conb_1
XFILLER_476_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[0\].yc la_data_in[96] blk.column\[0\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[0\].row\[1\].yc/confclk blk.column\[0\].row\[0\].yc/dempty blk.column\[0\].row\[0\].yc/din[0]
+ blk.column\[0\].row\[0\].yc/din[1] blk.column\[0\].row\[1\].yc/uin[0] blk.column\[0\].row\[1\].yc/uin[1]
+ blk.column\[0\].row\[0\].yc/hempty blk.column\[0\].row\[0\].yc/hempty2 blk.column\[0\].row\[0\].yc/lempty
+ blk.column\[0\].row\[0\].yc/lin[0] blk.column\[0\].row\[0\].yc/lin[1] blk.column\[1\].row\[0\].yc/rin[0]
+ blk.column\[1\].row\[0\].yc/rin[1] _428_/HI la_data_in[113] blk.column\[0\].row\[1\].yc/reset
+ _476_/LO _477_/LO blk.column\[0\].row\[0\].yc/rout[0] blk.column\[0\].row\[0\].yc/rout[1]
+ _478_/LO la_data_in[64] la_data_in[65] la_data_out[0] la_data_out[1] blk.column\[0\].row\[0\].yc/vempty
+ blk.column\[0\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_393_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_492_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_334_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_259_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_509_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_342_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_528_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_321_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_227_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_404_ _398_/X wbs_dat_o[16] _356_/A _403_/X VGND VGND VPWR VPWR _760_/D sky130_fd_sc_hd__o22a_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_335_ _335_/A VGND VGND VPWR VPWR _335_/Y sky130_fd_sc_hd__inv_2
XFILLER_375_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_291_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_319_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_307_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_384_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[8\].yc blk.column\[15\].row\[8\].yc/cbitin blk.column\[15\].row\[9\].yc/cbitin
+ blk.column\[15\].row\[8\].yc/confclk blk.column\[15\].row\[9\].yc/confclk blk.column\[15\].row\[8\].yc/dempty
+ blk.column\[15\].row\[8\].yc/din[0] blk.column\[15\].row\[8\].yc/din[1] blk.column\[15\].row\[9\].yc/uin[0]
+ blk.column\[15\].row\[9\].yc/uin[1] blk.column\[15\].row\[8\].yc/hempty blk.column\[14\].row\[8\].yc/lempty
+ _465_/HI _557_/LO _558_/LO blk.column\[15\].row\[8\].yc/lout[0] blk.column\[15\].row\[8\].yc/lout[1]
+ blk.column\[14\].row\[8\].yc/hempty blk.column\[15\].row\[8\].yc/reset blk.column\[15\].row\[9\].yc/reset
+ blk.column\[15\].row\[8\].yc/rin[0] blk.column\[15\].row\[8\].yc/rin[1] blk.column\[14\].row\[8\].yc/lin[0]
+ blk.column\[14\].row\[8\].yc/lin[1] blk.column\[15\].row\[8\].yc/uempty blk.column\[15\].row\[8\].yc/uin[0]
+ blk.column\[15\].row\[8\].yc/uin[1] blk.column\[15\].row\[7\].yc/din[0] blk.column\[15\].row\[7\].yc/din[1]
+ blk.column\[15\].row\[7\].yc/dempty blk.column\[15\].row\[9\].yc/uempty VPWR VGND
+ ycell
XFILLER_177_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_524_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_434_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xblk.column\[6\].row\[9\].yc blk.column\[6\].row\[9\].yc/cbitin blk.column\[6\].row\[9\].yc/cbitout
+ blk.column\[6\].row\[9\].yc/confclk blk.column\[6\].row\[9\].yc/confclko blk.column\[6\].row\[9\].yc/dempty
+ blk.column\[6\].row\[9\].yc/din[0] blk.column\[6\].row\[9\].yc/din[1] blk.column\[6\].row\[9\].yc/dout[0]
+ blk.column\[6\].row\[9\].yc/dout[1] blk.column\[6\].row\[9\].yc/hempty blk.column\[5\].row\[9\].yc/lempty
+ blk.column\[6\].row\[9\].yc/lempty blk.column\[6\].row\[9\].yc/lin[0] blk.column\[6\].row\[9\].yc/lin[1]
+ blk.column\[7\].row\[9\].yc/rin[0] blk.column\[7\].row\[9\].yc/rin[1] blk.column\[5\].row\[9\].yc/hempty
+ blk.column\[6\].row\[9\].yc/reset blk.column\[6\].row\[9\].yc/reseto blk.column\[6\].row\[9\].yc/rin[0]
+ blk.column\[6\].row\[9\].yc/rin[1] blk.column\[5\].row\[9\].yc/lin[0] blk.column\[5\].row\[9\].yc/lin[1]
+ blk.column\[6\].row\[9\].yc/uempty blk.column\[6\].row\[9\].yc/uin[0] blk.column\[6\].row\[9\].yc/uin[1]
+ blk.column\[6\].row\[8\].yc/din[0] blk.column\[6\].row\[8\].yc/din[1] blk.column\[6\].row\[8\].yc/dempty
+ blk.column\[6\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_520_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_383_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_320_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_344_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_507_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_318_ _317_/X VGND VGND VPWR VPWR _319_/A sky130_fd_sc_hd__buf_2
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_534_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_331_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_485_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_334_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_503_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_415_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_311_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_489_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_367_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_432_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_243_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_244_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1010 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_478_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_411_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_374_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[1\].yc blk.column\[10\].row\[1\].yc/cbitin blk.column\[10\].row\[2\].yc/cbitin
+ blk.column\[10\].row\[1\].yc/confclk blk.column\[10\].row\[2\].yc/confclk blk.column\[10\].row\[1\].yc/dempty
+ blk.column\[10\].row\[1\].yc/din[0] blk.column\[10\].row\[1\].yc/din[1] blk.column\[10\].row\[2\].yc/uin[0]
+ blk.column\[10\].row\[2\].yc/uin[1] blk.column\[10\].row\[1\].yc/hempty blk.column\[9\].row\[1\].yc/lempty
+ blk.column\[10\].row\[1\].yc/lempty blk.column\[10\].row\[1\].yc/lin[0] blk.column\[10\].row\[1\].yc/lin[1]
+ blk.column\[11\].row\[1\].yc/rin[0] blk.column\[11\].row\[1\].yc/rin[1] blk.column\[9\].row\[1\].yc/hempty
+ blk.column\[10\].row\[1\].yc/reset blk.column\[10\].row\[2\].yc/reset blk.column\[9\].row\[1\].yc/lout[0]
+ blk.column\[9\].row\[1\].yc/lout[1] blk.column\[9\].row\[1\].yc/lin[0] blk.column\[9\].row\[1\].yc/lin[1]
+ blk.column\[10\].row\[1\].yc/uempty blk.column\[10\].row\[1\].yc/uin[0] blk.column\[10\].row\[1\].yc/uin[1]
+ blk.column\[10\].row\[0\].yc/din[0] blk.column\[10\].row\[0\].yc/din[1] blk.column\[10\].row\[0\].yc/dempty
+ blk.column\[10\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_136_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_335_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_798_ wb_clk_i _798_/D VGND VGND VPWR VPWR _321_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_5_1890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[2\].yc blk.column\[1\].row\[2\].yc/cbitin blk.column\[1\].row\[3\].yc/cbitin
+ blk.column\[1\].row\[2\].yc/confclk blk.column\[1\].row\[3\].yc/confclk blk.column\[1\].row\[2\].yc/dempty
+ blk.column\[1\].row\[2\].yc/din[0] blk.column\[1\].row\[2\].yc/din[1] blk.column\[1\].row\[3\].yc/uin[0]
+ blk.column\[1\].row\[3\].yc/uin[1] blk.column\[1\].row\[2\].yc/hempty blk.column\[0\].row\[2\].yc/lempty
+ blk.column\[1\].row\[2\].yc/lempty blk.column\[1\].row\[2\].yc/lin[0] blk.column\[1\].row\[2\].yc/lin[1]
+ blk.column\[2\].row\[2\].yc/rin[0] blk.column\[2\].row\[2\].yc/rin[1] blk.column\[0\].row\[2\].yc/hempty
+ blk.column\[1\].row\[2\].yc/reset blk.column\[1\].row\[3\].yc/reset blk.column\[1\].row\[2\].yc/rin[0]
+ blk.column\[1\].row\[2\].yc/rin[1] blk.column\[0\].row\[2\].yc/lin[0] blk.column\[0\].row\[2\].yc/lin[1]
+ blk.column\[1\].row\[2\].yc/uempty blk.column\[1\].row\[2\].yc/uin[0] blk.column\[1\].row\[2\].yc/uin[1]
+ blk.column\[1\].row\[1\].yc/din[0] blk.column\[1\].row\[1\].yc/din[1] blk.column\[1\].row\[1\].yc/dempty
+ blk.column\[1\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_499_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_403_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[12\].yc blk.column\[5\].row\[12\].yc/cbitin blk.column\[5\].row\[13\].yc/cbitin
+ blk.column\[5\].row\[12\].yc/confclk blk.column\[5\].row\[13\].yc/confclk blk.column\[5\].row\[12\].yc/dempty
+ blk.column\[5\].row\[12\].yc/din[0] blk.column\[5\].row\[12\].yc/din[1] blk.column\[5\].row\[13\].yc/uin[0]
+ blk.column\[5\].row\[13\].yc/uin[1] blk.column\[5\].row\[12\].yc/hempty blk.column\[4\].row\[12\].yc/lempty
+ blk.column\[5\].row\[12\].yc/lempty blk.column\[5\].row\[12\].yc/lin[0] blk.column\[5\].row\[12\].yc/lin[1]
+ blk.column\[6\].row\[12\].yc/rin[0] blk.column\[6\].row\[12\].yc/rin[1] blk.column\[4\].row\[12\].yc/hempty
+ blk.column\[5\].row\[12\].yc/reset blk.column\[5\].row\[13\].yc/reset blk.column\[5\].row\[12\].yc/rin[0]
+ blk.column\[5\].row\[12\].yc/rin[1] blk.column\[4\].row\[12\].yc/lin[0] blk.column\[4\].row\[12\].yc/lin[1]
+ blk.column\[5\].row\[12\].yc/uempty blk.column\[5\].row\[12\].yc/uin[0] blk.column\[5\].row\[12\].yc/uin[1]
+ blk.column\[5\].row\[11\].yc/din[0] blk.column\[5\].row\[11\].yc/din[1] blk.column\[5\].row\[11\].yc/dempty
+ blk.column\[5\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_414_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_335_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_536_1893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_721_ VGND VGND VPWR VPWR _721_/HI la_data_out[105] sky130_fd_sc_hd__conb_1
XPHY_7267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_483_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_652_ VGND VGND VPWR VPWR _652_/HI io_out[26] sky130_fd_sc_hd__conb_1
XPHY_5832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_361_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_583_ VGND VGND VPWR VPWR _583_/HI _583_/LO sky130_fd_sc_hd__conb_1
XFILLER_508_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_508_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_485_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_509_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_507_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_522_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_542_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_258_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_525_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_534_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_486_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_442_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_493_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_325_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_538_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_532_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_500_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_704_ VGND VGND VPWR VPWR _704_/HI la_data_out[88] sky130_fd_sc_hd__conb_1
XPHY_6352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_635_ VGND VGND VPWR VPWR _635_/HI io_out[9] sky130_fd_sc_hd__conb_1
XFILLER_504_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_566_ VGND VGND VPWR VPWR _566_/HI _566_/LO sky130_fd_sc_hd__conb_1
XFILLER_400_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_497_ VGND VGND VPWR VPWR _497_/HI _497_/LO sky130_fd_sc_hd__conb_1
Xblk.column\[12\].row\[14\].yc blk.column\[12\].row\[14\].yc/cbitin blk.column\[12\].row\[15\].yc/cbitin
+ blk.column\[12\].row\[14\].yc/confclk blk.column\[12\].row\[15\].yc/confclk blk.column\[12\].row\[14\].yc/dempty
+ blk.column\[12\].row\[14\].yc/din[0] blk.column\[12\].row\[14\].yc/din[1] blk.column\[12\].row\[15\].yc/uin[0]
+ blk.column\[12\].row\[15\].yc/uin[1] blk.column\[12\].row\[14\].yc/hempty blk.column\[11\].row\[14\].yc/lempty
+ blk.column\[12\].row\[14\].yc/lempty blk.column\[12\].row\[14\].yc/lin[0] blk.column\[12\].row\[14\].yc/lin[1]
+ blk.column\[13\].row\[14\].yc/rin[0] blk.column\[13\].row\[14\].yc/rin[1] blk.column\[11\].row\[14\].yc/hempty
+ blk.column\[12\].row\[14\].yc/reset blk.column\[12\].row\[15\].yc/reset blk.column\[12\].row\[14\].yc/rin[0]
+ blk.column\[12\].row\[14\].yc/rin[1] blk.column\[11\].row\[14\].yc/lin[0] blk.column\[11\].row\[14\].yc/lin[1]
+ blk.column\[12\].row\[14\].yc/uempty blk.column\[12\].row\[14\].yc/uin[0] blk.column\[12\].row\[14\].yc/uin[1]
+ blk.column\[12\].row\[13\].yc/din[0] blk.column\[12\].row\[13\].yc/din[1] blk.column\[12\].row\[13\].yc/dempty
+ blk.column\[12\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_537_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_527_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_396_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_312_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_494_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_442_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_420_ _419_/X wbs_dat_o[5] _805_/Q _417_/X VGND VGND VPWR VPWR _420_/X sky130_fd_sc_hd__o22a_4
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_351_ _786_/Q VGND VGND VPWR VPWR _351_/Y sky130_fd_sc_hd__inv_2
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_497_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_358_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[3\].yc blk.column\[11\].row\[3\].yc/cbitin blk.column\[11\].row\[4\].yc/cbitin
+ blk.column\[11\].row\[3\].yc/confclk blk.column\[11\].row\[4\].yc/confclk blk.column\[11\].row\[3\].yc/dempty
+ blk.column\[11\].row\[3\].yc/din[0] blk.column\[11\].row\[3\].yc/din[1] blk.column\[11\].row\[4\].yc/uin[0]
+ blk.column\[11\].row\[4\].yc/uin[1] blk.column\[11\].row\[3\].yc/hempty blk.column\[10\].row\[3\].yc/lempty
+ blk.column\[11\].row\[3\].yc/lempty blk.column\[11\].row\[3\].yc/lin[0] blk.column\[11\].row\[3\].yc/lin[1]
+ blk.column\[12\].row\[3\].yc/rin[0] blk.column\[12\].row\[3\].yc/rin[1] blk.column\[10\].row\[3\].yc/hempty
+ blk.column\[11\].row\[3\].yc/reset blk.column\[11\].row\[4\].yc/reset blk.column\[11\].row\[3\].yc/rin[0]
+ blk.column\[11\].row\[3\].yc/rin[1] blk.column\[10\].row\[3\].yc/lin[0] blk.column\[10\].row\[3\].yc/lin[1]
+ blk.column\[11\].row\[3\].yc/uempty blk.column\[11\].row\[3\].yc/uin[0] blk.column\[11\].row\[3\].yc/uin[1]
+ blk.column\[11\].row\[2\].yc/din[0] blk.column\[11\].row\[2\].yc/din[1] blk.column\[11\].row\[2\].yc/dempty
+ blk.column\[11\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_518_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_311_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_330_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[4\].yc blk.column\[2\].row\[4\].yc/cbitin blk.column\[2\].row\[5\].yc/cbitin
+ blk.column\[2\].row\[4\].yc/confclk blk.column\[2\].row\[5\].yc/confclk blk.column\[2\].row\[4\].yc/dempty
+ blk.column\[2\].row\[4\].yc/din[0] blk.column\[2\].row\[4\].yc/din[1] blk.column\[2\].row\[5\].yc/uin[0]
+ blk.column\[2\].row\[5\].yc/uin[1] blk.column\[2\].row\[4\].yc/hempty blk.column\[1\].row\[4\].yc/lempty
+ blk.column\[2\].row\[4\].yc/lempty blk.column\[2\].row\[4\].yc/lin[0] blk.column\[2\].row\[4\].yc/lin[1]
+ blk.column\[3\].row\[4\].yc/rin[0] blk.column\[3\].row\[4\].yc/rin[1] blk.column\[1\].row\[4\].yc/hempty
+ blk.column\[2\].row\[4\].yc/reset blk.column\[2\].row\[5\].yc/reset blk.column\[2\].row\[4\].yc/rin[0]
+ blk.column\[2\].row\[4\].yc/rin[1] blk.column\[1\].row\[4\].yc/lin[0] blk.column\[1\].row\[4\].yc/lin[1]
+ blk.column\[2\].row\[4\].yc/uempty blk.column\[2\].row\[4\].yc/uin[0] blk.column\[2\].row\[4\].yc/uin[1]
+ blk.column\[2\].row\[3\].yc/din[0] blk.column\[2\].row\[3\].yc/din[1] blk.column\[2\].row\[3\].yc/dempty
+ blk.column\[2\].row\[5\].yc/uempty VPWR VGND ycell
XPHY_11564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_326_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_413_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_618_ VGND VGND VPWR VPWR _618_/HI io_oeb[30] sky130_fd_sc_hd__conb_1
XFILLER_504_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_308_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_388_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_549_ VGND VGND VPWR VPWR _549_/HI _549_/LO sky130_fd_sc_hd__conb_1
XFILLER_144_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[15\].yc blk.column\[9\].row\[15\].yc/cbitin la_data_out[41]
+ blk.column\[9\].row\[15\].yc/confclk blk.column\[9\].row\[15\].yc/confclko _475_/HI
+ _586_/LO _587_/LO blk.column\[9\].row\[15\].yc/dout[0] blk.column\[9\].row\[15\].yc/dout[1]
+ blk.column\[9\].row\[15\].yc/hempty blk.column\[8\].row\[15\].yc/lempty blk.column\[9\].row\[15\].yc/lempty
+ blk.column\[9\].row\[15\].yc/lin[0] blk.column\[9\].row\[15\].yc/lin[1] blk.column\[9\].row\[15\].yc/lout[0]
+ blk.column\[9\].row\[15\].yc/lout[1] blk.column\[8\].row\[15\].yc/hempty blk.column\[9\].row\[15\].yc/reset
+ blk.column\[9\].row\[15\].yc/reseto blk.column\[9\].row\[15\].yc/rin[0] blk.column\[9\].row\[15\].yc/rin[1]
+ blk.column\[8\].row\[15\].yc/lin[0] blk.column\[8\].row\[15\].yc/lin[1] blk.column\[9\].row\[15\].yc/uempty
+ blk.column\[9\].row\[15\].yc/uin[0] blk.column\[9\].row\[15\].yc/uin[1] blk.column\[9\].row\[14\].yc/din[0]
+ blk.column\[9\].row\[14\].yc/din[1] blk.column\[9\].row\[14\].yc/dempty blk.column\[9\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_378_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_257_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_419_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_487_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_503_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_369_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_412_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_298_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_377_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_448_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_439_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_413_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_403_ wb_rst_i VGND VGND VPWR VPWR _403_/X sky130_fd_sc_hd__buf_2
XFILLER_50_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_358_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_521_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_334_ _333_/Y _331_/X wbs_dat_i[9] _331_/X VGND VGND VPWR VPWR _334_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_19_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_278_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_375_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_482_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_517_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[13\].yc blk.column\[0\].row\[13\].yc/cbitin blk.column\[0\].row\[14\].yc/cbitin
+ blk.column\[0\].row\[13\].yc/confclk blk.column\[0\].row\[14\].yc/confclk blk.column\[0\].row\[13\].yc/dempty
+ blk.column\[0\].row\[13\].yc/din[0] blk.column\[0\].row\[13\].yc/din[1] blk.column\[0\].row\[14\].yc/uin[0]
+ blk.column\[0\].row\[14\].yc/uin[1] blk.column\[0\].row\[13\].yc/hempty blk.column\[0\].row\[13\].yc/hempty2
+ blk.column\[0\].row\[13\].yc/lempty blk.column\[0\].row\[13\].yc/lin[0] blk.column\[0\].row\[13\].yc/lin[1]
+ blk.column\[1\].row\[13\].yc/rin[0] blk.column\[1\].row\[13\].yc/rin[1] _432_/HI
+ blk.column\[0\].row\[13\].yc/reset blk.column\[0\].row\[14\].yc/reset _485_/LO _486_/LO
+ blk.column\[0\].row\[13\].yc/rout[0] blk.column\[0\].row\[13\].yc/rout[1] blk.column\[0\].row\[13\].yc/uempty
+ blk.column\[0\].row\[13\].yc/uin[0] blk.column\[0\].row\[13\].yc/uin[1] blk.column\[0\].row\[12\].yc/din[0]
+ blk.column\[0\].row\[12\].yc/din[1] blk.column\[0\].row\[12\].yc/dempty blk.column\[0\].row\[14\].yc/uempty
+ VPWR VGND ycell
XFILLER_322_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_520_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_450_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_530_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_372_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_513_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_391_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_483_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_317_ _295_/Y wbs_we_i wbs_sel_i[1] VGND VGND VPWR VPWR _317_/X sky130_fd_sc_hd__and3_4
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_455_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_418_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_473_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_408_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_449_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_508_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[5\].yc blk.column\[12\].row\[5\].yc/cbitin blk.column\[12\].row\[6\].yc/cbitin
+ blk.column\[12\].row\[5\].yc/confclk blk.column\[12\].row\[6\].yc/confclk blk.column\[12\].row\[5\].yc/dempty
+ blk.column\[12\].row\[5\].yc/din[0] blk.column\[12\].row\[5\].yc/din[1] blk.column\[12\].row\[6\].yc/uin[0]
+ blk.column\[12\].row\[6\].yc/uin[1] blk.column\[12\].row\[5\].yc/hempty blk.column\[11\].row\[5\].yc/lempty
+ blk.column\[12\].row\[5\].yc/lempty blk.column\[12\].row\[5\].yc/lin[0] blk.column\[12\].row\[5\].yc/lin[1]
+ blk.column\[13\].row\[5\].yc/rin[0] blk.column\[13\].row\[5\].yc/rin[1] blk.column\[11\].row\[5\].yc/hempty
+ blk.column\[12\].row\[5\].yc/reset blk.column\[12\].row\[6\].yc/reset blk.column\[12\].row\[5\].yc/rin[0]
+ blk.column\[12\].row\[5\].yc/rin[1] blk.column\[11\].row\[5\].yc/lin[0] blk.column\[11\].row\[5\].yc/lin[1]
+ blk.column\[12\].row\[5\].yc/uempty blk.column\[12\].row\[5\].yc/uin[0] blk.column\[12\].row\[5\].yc/uin[1]
+ blk.column\[12\].row\[4\].yc/din[0] blk.column\[12\].row\[4\].yc/din[1] blk.column\[12\].row\[4\].yc/dempty
+ blk.column\[12\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_528_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_389_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_385_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_486_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_355_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_404_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[6\].yc blk.column\[3\].row\[6\].yc/cbitin blk.column\[3\].row\[7\].yc/cbitin
+ blk.column\[3\].row\[6\].yc/confclk blk.column\[3\].row\[7\].yc/confclk blk.column\[3\].row\[6\].yc/dempty
+ blk.column\[3\].row\[6\].yc/din[0] blk.column\[3\].row\[6\].yc/din[1] blk.column\[3\].row\[7\].yc/uin[0]
+ blk.column\[3\].row\[7\].yc/uin[1] blk.column\[3\].row\[6\].yc/hempty blk.column\[2\].row\[6\].yc/lempty
+ blk.column\[3\].row\[6\].yc/lempty blk.column\[3\].row\[6\].yc/lin[0] blk.column\[3\].row\[6\].yc/lin[1]
+ blk.column\[4\].row\[6\].yc/rin[0] blk.column\[4\].row\[6\].yc/rin[1] blk.column\[2\].row\[6\].yc/hempty
+ blk.column\[3\].row\[6\].yc/reset blk.column\[3\].row\[7\].yc/reset blk.column\[3\].row\[6\].yc/rin[0]
+ blk.column\[3\].row\[6\].yc/rin[1] blk.column\[2\].row\[6\].yc/lin[0] blk.column\[2\].row\[6\].yc/lin[1]
+ blk.column\[3\].row\[6\].yc/uempty blk.column\[3\].row\[6\].yc/uin[0] blk.column\[3\].row\[6\].yc/uin[1]
+ blk.column\[3\].row\[5\].yc/din[0] blk.column\[3\].row\[5\].yc/din[1] blk.column\[3\].row\[5\].yc/dempty
+ blk.column\[3\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_499_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_371_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_371_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_542_2202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_362_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_797_ wb_clk_i _797_/D VGND VGND VPWR VPWR _323_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_542_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_423_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_524_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_336_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_534_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_514_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_257_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_521_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_421_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_274_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[0\].yc la_data_in[104] blk.column\[8\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[8\].row\[1\].yc/confclk blk.column\[8\].row\[0\].yc/dempty blk.column\[8\].row\[0\].yc/din[0]
+ blk.column\[8\].row\[0\].yc/din[1] blk.column\[8\].row\[1\].yc/uin[0] blk.column\[8\].row\[1\].yc/uin[1]
+ blk.column\[8\].row\[0\].yc/hempty blk.column\[7\].row\[0\].yc/lempty blk.column\[8\].row\[0\].yc/lempty
+ blk.column\[8\].row\[0\].yc/lin[0] blk.column\[8\].row\[0\].yc/lin[1] blk.column\[9\].row\[0\].yc/rin[0]
+ blk.column\[9\].row\[0\].yc/rin[1] blk.column\[7\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[8\].row\[1\].yc/reset blk.column\[8\].row\[0\].yc/rin[0] blk.column\[8\].row\[0\].yc/rin[1]
+ blk.column\[7\].row\[0\].yc/lin[0] blk.column\[7\].row\[0\].yc/lin[1] _582_/LO la_data_in[80]
+ la_data_in[81] la_data_out[16] la_data_out[17] blk.column\[8\].row\[0\].yc/vempty
+ blk.column\[8\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_497_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_720_ VGND VGND VPWR VPWR _720_/HI la_data_out[104] sky130_fd_sc_hd__conb_1
XFILLER_102_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_480_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_651_ VGND VGND VPWR VPWR _651_/HI io_out[25] sky130_fd_sc_hd__conb_1
XPHY_6556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_582_ VGND VGND VPWR VPWR _582_/HI _582_/LO sky130_fd_sc_hd__conb_1
XFILLER_496_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_354_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_357_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_385_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_462_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_522_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_494_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_449_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_265_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_364_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_253_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_276_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_703_ VGND VGND VPWR VPWR _703_/HI la_data_out[87] sky130_fd_sc_hd__conb_1
XPHY_6353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_634_ VGND VGND VPWR VPWR _634_/HI io_out[8] sky130_fd_sc_hd__conb_1
XPHY_6386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_565_ VGND VGND VPWR VPWR _565_/HI _565_/LO sky130_fd_sc_hd__conb_1
XPHY_5696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_400_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_496_ VGND VGND VPWR VPWR _496_/HI _496_/LO sky130_fd_sc_hd__conb_1
XFILLER_301_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_522_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_411_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_498_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_535_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[7\].yc blk.column\[13\].row\[7\].yc/cbitin blk.column\[13\].row\[8\].yc/cbitin
+ blk.column\[13\].row\[7\].yc/confclk blk.column\[13\].row\[8\].yc/confclk blk.column\[13\].row\[7\].yc/dempty
+ blk.column\[13\].row\[7\].yc/din[0] blk.column\[13\].row\[7\].yc/din[1] blk.column\[13\].row\[8\].yc/uin[0]
+ blk.column\[13\].row\[8\].yc/uin[1] blk.column\[13\].row\[7\].yc/hempty blk.column\[12\].row\[7\].yc/lempty
+ blk.column\[13\].row\[7\].yc/lempty blk.column\[13\].row\[7\].yc/lin[0] blk.column\[13\].row\[7\].yc/lin[1]
+ blk.column\[14\].row\[7\].yc/rin[0] blk.column\[14\].row\[7\].yc/rin[1] blk.column\[12\].row\[7\].yc/hempty
+ blk.column\[13\].row\[7\].yc/reset blk.column\[13\].row\[8\].yc/reset blk.column\[13\].row\[7\].yc/rin[0]
+ blk.column\[13\].row\[7\].yc/rin[1] blk.column\[12\].row\[7\].yc/lin[0] blk.column\[12\].row\[7\].yc/lin[1]
+ blk.column\[13\].row\[7\].yc/uempty blk.column\[13\].row\[7\].yc/uin[0] blk.column\[13\].row\[7\].yc/uin[1]
+ blk.column\[13\].row\[6\].yc/din[0] blk.column\[13\].row\[6\].yc/din[1] blk.column\[13\].row\[6\].yc/dempty
+ blk.column\[13\].row\[8\].yc/uempty VPWR VGND ycell
XPHY_10308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ _349_/Y _345_/X wbs_dat_i[19] _345_/X VGND VGND VPWR VPWR _787_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[4\].row\[8\].yc blk.column\[4\].row\[8\].yc/cbitin blk.column\[4\].row\[9\].yc/cbitin
+ blk.column\[4\].row\[8\].yc/confclk blk.column\[4\].row\[9\].yc/confclk blk.column\[4\].row\[8\].yc/dempty
+ blk.column\[4\].row\[8\].yc/din[0] blk.column\[4\].row\[8\].yc/din[1] blk.column\[4\].row\[9\].yc/uin[0]
+ blk.column\[4\].row\[9\].yc/uin[1] blk.column\[4\].row\[8\].yc/hempty blk.column\[3\].row\[8\].yc/lempty
+ blk.column\[4\].row\[8\].yc/lempty blk.column\[4\].row\[8\].yc/lin[0] blk.column\[4\].row\[8\].yc/lin[1]
+ blk.column\[5\].row\[8\].yc/rin[0] blk.column\[5\].row\[8\].yc/rin[1] blk.column\[3\].row\[8\].yc/hempty
+ blk.column\[4\].row\[8\].yc/reset blk.column\[4\].row\[9\].yc/reset blk.column\[4\].row\[8\].yc/rin[0]
+ blk.column\[4\].row\[8\].yc/rin[1] blk.column\[3\].row\[8\].yc/lin[0] blk.column\[3\].row\[8\].yc/lin[1]
+ blk.column\[4\].row\[8\].yc/uempty blk.column\[4\].row\[8\].yc/uin[0] blk.column\[4\].row\[8\].yc/uin[1]
+ blk.column\[4\].row\[7\].yc/din[0] blk.column\[4\].row\[7\].yc/din[1] blk.column\[4\].row\[7\].yc/dempty
+ blk.column\[4\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_505_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_478_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_536_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_497_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_529_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_347_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_370_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_512_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_527_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_413_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_617_ VGND VGND VPWR VPWR _617_/HI io_oeb[29] sky130_fd_sc_hd__conb_1
XPHY_5482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_548_ VGND VGND VPWR VPWR _548_/HI _548_/LO sky130_fd_sc_hd__conb_1
XFILLER_232_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_479_ VGND VGND VPWR VPWR _479_/HI _479_/LO sky130_fd_sc_hd__conb_1
XFILLER_179_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_346_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_523_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_485_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_522_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_322_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_448_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_492_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_527_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[2\].yc blk.column\[9\].row\[2\].yc/cbitin blk.column\[9\].row\[3\].yc/cbitin
+ blk.column\[9\].row\[2\].yc/confclk blk.column\[9\].row\[3\].yc/confclk blk.column\[9\].row\[2\].yc/dempty
+ blk.column\[9\].row\[2\].yc/din[0] blk.column\[9\].row\[2\].yc/din[1] blk.column\[9\].row\[3\].yc/uin[0]
+ blk.column\[9\].row\[3\].yc/uin[1] blk.column\[9\].row\[2\].yc/hempty blk.column\[8\].row\[2\].yc/lempty
+ blk.column\[9\].row\[2\].yc/lempty blk.column\[9\].row\[2\].yc/lin[0] blk.column\[9\].row\[2\].yc/lin[1]
+ blk.column\[9\].row\[2\].yc/lout[0] blk.column\[9\].row\[2\].yc/lout[1] blk.column\[8\].row\[2\].yc/hempty
+ blk.column\[9\].row\[2\].yc/reset blk.column\[9\].row\[3\].yc/reset blk.column\[9\].row\[2\].yc/rin[0]
+ blk.column\[9\].row\[2\].yc/rin[1] blk.column\[8\].row\[2\].yc/lin[0] blk.column\[8\].row\[2\].yc/lin[1]
+ blk.column\[9\].row\[2\].yc/uempty blk.column\[9\].row\[2\].yc/uin[0] blk.column\[9\].row\[2\].yc/uin[1]
+ blk.column\[9\].row\[1\].yc/din[0] blk.column\[9\].row\[1\].yc/din[1] blk.column\[9\].row\[1\].yc/dempty
+ blk.column\[9\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_195_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_429_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[11\].yc blk.column\[6\].row\[11\].yc/cbitin blk.column\[6\].row\[12\].yc/cbitin
+ blk.column\[6\].row\[11\].yc/confclk blk.column\[6\].row\[12\].yc/confclk blk.column\[6\].row\[11\].yc/dempty
+ blk.column\[6\].row\[11\].yc/din[0] blk.column\[6\].row\[11\].yc/din[1] blk.column\[6\].row\[12\].yc/uin[0]
+ blk.column\[6\].row\[12\].yc/uin[1] blk.column\[6\].row\[11\].yc/hempty blk.column\[5\].row\[11\].yc/lempty
+ blk.column\[6\].row\[11\].yc/lempty blk.column\[6\].row\[11\].yc/lin[0] blk.column\[6\].row\[11\].yc/lin[1]
+ blk.column\[7\].row\[11\].yc/rin[0] blk.column\[7\].row\[11\].yc/rin[1] blk.column\[5\].row\[11\].yc/hempty
+ blk.column\[6\].row\[11\].yc/reset blk.column\[6\].row\[12\].yc/reset blk.column\[6\].row\[11\].yc/rin[0]
+ blk.column\[6\].row\[11\].yc/rin[1] blk.column\[5\].row\[11\].yc/lin[0] blk.column\[5\].row\[11\].yc/lin[1]
+ blk.column\[6\].row\[11\].yc/uempty blk.column\[6\].row\[11\].yc/uin[0] blk.column\[6\].row\[11\].yc/uin[1]
+ blk.column\[6\].row\[10\].yc/din[0] blk.column\[6\].row\[10\].yc/din[1] blk.column\[6\].row\[10\].yc/dempty
+ blk.column\[6\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_494_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_447_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_402_ _398_/X wbs_dat_o[17] _354_/A _396_/X VGND VGND VPWR VPWR _761_/D sky130_fd_sc_hd__o22a_4
XFILLER_14_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_434_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_509_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_333_ _333_/A VGND VGND VPWR VPWR _333_/Y sky130_fd_sc_hd__inv_2
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_358_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_375_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_471_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_390_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_331_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_11384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_252_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_517_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_530_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_528_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_459_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_498_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_320_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_516_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_429_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_409_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_369_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_316_ _316_/A VGND VGND VPWR VPWR _316_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_514_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_502_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[13\].yc blk.column\[13\].row\[13\].yc/cbitin blk.column\[13\].row\[14\].yc/cbitin
+ blk.column\[13\].row\[13\].yc/confclk blk.column\[13\].row\[14\].yc/confclk blk.column\[13\].row\[13\].yc/dempty
+ blk.column\[13\].row\[13\].yc/din[0] blk.column\[13\].row\[13\].yc/din[1] blk.column\[13\].row\[14\].yc/uin[0]
+ blk.column\[13\].row\[14\].yc/uin[1] blk.column\[13\].row\[13\].yc/hempty blk.column\[12\].row\[13\].yc/lempty
+ blk.column\[13\].row\[13\].yc/lempty blk.column\[13\].row\[13\].yc/lin[0] blk.column\[13\].row\[13\].yc/lin[1]
+ blk.column\[14\].row\[13\].yc/rin[0] blk.column\[14\].row\[13\].yc/rin[1] blk.column\[12\].row\[13\].yc/hempty
+ blk.column\[13\].row\[13\].yc/reset blk.column\[13\].row\[14\].yc/reset blk.column\[13\].row\[13\].yc/rin[0]
+ blk.column\[13\].row\[13\].yc/rin[1] blk.column\[12\].row\[13\].yc/lin[0] blk.column\[12\].row\[13\].yc/lin[1]
+ blk.column\[13\].row\[13\].yc/uempty blk.column\[13\].row\[13\].yc/uin[0] blk.column\[13\].row\[13\].yc/uin[1]
+ blk.column\[13\].row\[12\].yc/din[0] blk.column\[13\].row\[12\].yc/din[1] blk.column\[13\].row\[12\].yc/dempty
+ blk.column\[13\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_33_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_240_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_509_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_354_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[9\].yc blk.column\[14\].row\[9\].yc/cbitin blk.column\[14\].row\[9\].yc/cbitout
+ blk.column\[14\].row\[9\].yc/confclk blk.column\[14\].row\[9\].yc/confclko blk.column\[14\].row\[9\].yc/dempty
+ blk.column\[14\].row\[9\].yc/din[0] blk.column\[14\].row\[9\].yc/din[1] blk.column\[14\].row\[9\].yc/dout[0]
+ blk.column\[14\].row\[9\].yc/dout[1] blk.column\[14\].row\[9\].yc/hempty blk.column\[13\].row\[9\].yc/lempty
+ blk.column\[14\].row\[9\].yc/lempty blk.column\[14\].row\[9\].yc/lin[0] blk.column\[14\].row\[9\].yc/lin[1]
+ blk.column\[15\].row\[9\].yc/rin[0] blk.column\[15\].row\[9\].yc/rin[1] blk.column\[13\].row\[9\].yc/hempty
+ blk.column\[14\].row\[9\].yc/reset blk.column\[14\].row\[9\].yc/reseto blk.column\[14\].row\[9\].yc/rin[0]
+ blk.column\[14\].row\[9\].yc/rin[1] blk.column\[13\].row\[9\].yc/lin[0] blk.column\[13\].row\[9\].yc/lin[1]
+ blk.column\[14\].row\[9\].yc/uempty blk.column\[14\].row\[9\].yc/uin[0] blk.column\[14\].row\[9\].yc/uin[1]
+ blk.column\[14\].row\[8\].yc/din[0] blk.column\[14\].row\[8\].yc/din[1] blk.column\[14\].row\[8\].yc/dempty
+ blk.column\[14\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_468_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_502_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_478_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_459_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_385_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_419_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_419_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_507_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_796_ wb_clk_i _327_/X VGND VGND VPWR VPWR _326_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_5_1870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_503_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_381_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_396_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_329_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_336_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_490_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_531_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_456_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_438_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_530_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_650_ VGND VGND VPWR VPWR _650_/HI io_out[24] sky130_fd_sc_hd__conb_1
XPHY_6557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_581_ VGND VGND VPWR VPWR _581_/HI _581_/LO sky130_fd_sc_hd__conb_1
XPHY_5867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_496_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_514_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_366_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_318_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_253_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_341_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_531_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_779_ wb_clk_i _779_/D VGND VGND VPWR VPWR _779_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_79_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[3\].yc blk.column\[0\].row\[3\].yc/cbitin blk.column\[0\].row\[4\].yc/cbitin
+ blk.column\[0\].row\[3\].yc/confclk blk.column\[0\].row\[4\].yc/confclk blk.column\[0\].row\[4\].yc/vempty
+ blk.column\[0\].row\[3\].yc/din[0] blk.column\[0\].row\[3\].yc/din[1] blk.column\[0\].row\[4\].yc/uin[0]
+ blk.column\[0\].row\[4\].yc/uin[1] blk.column\[0\].row\[3\].yc/hempty blk.column\[0\].row\[3\].yc/hempty2
+ blk.column\[0\].row\[3\].yc/lempty blk.column\[0\].row\[3\].yc/lin[0] blk.column\[0\].row\[3\].yc/lin[1]
+ blk.column\[1\].row\[3\].yc/rin[0] blk.column\[1\].row\[3\].yc/rin[1] _438_/HI blk.column\[0\].row\[3\].yc/reset
+ blk.column\[0\].row\[4\].yc/reset _497_/LO _498_/LO blk.column\[0\].row\[3\].yc/rout[0]
+ blk.column\[0\].row\[3\].yc/rout[1] blk.column\[0\].row\[3\].yc/uempty blk.column\[0\].row\[3\].yc/uin[0]
+ blk.column\[0\].row\[3\].yc/uin[1] blk.column\[0\].row\[2\].yc/din[0] blk.column\[0\].row\[2\].yc/din[1]
+ blk.column\[0\].row\[2\].yc/dempty blk.column\[0\].row\[4\].yc/uempty VPWR VGND
+ ycell
XFILLER_520_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_525_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_522_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_364_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_221_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_517_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_495_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[12\].yc blk.column\[1\].row\[12\].yc/cbitin blk.column\[1\].row\[13\].yc/cbitin
+ blk.column\[1\].row\[12\].yc/confclk blk.column\[1\].row\[13\].yc/confclk blk.column\[1\].row\[12\].yc/dempty
+ blk.column\[1\].row\[12\].yc/din[0] blk.column\[1\].row\[12\].yc/din[1] blk.column\[1\].row\[13\].yc/uin[0]
+ blk.column\[1\].row\[13\].yc/uin[1] blk.column\[1\].row\[12\].yc/hempty blk.column\[0\].row\[12\].yc/lempty
+ blk.column\[1\].row\[12\].yc/lempty blk.column\[1\].row\[12\].yc/lin[0] blk.column\[1\].row\[12\].yc/lin[1]
+ blk.column\[2\].row\[12\].yc/rin[0] blk.column\[2\].row\[12\].yc/rin[1] blk.column\[0\].row\[12\].yc/hempty
+ blk.column\[1\].row\[12\].yc/reset blk.column\[1\].row\[13\].yc/reset blk.column\[1\].row\[12\].yc/rin[0]
+ blk.column\[1\].row\[12\].yc/rin[1] blk.column\[0\].row\[12\].yc/lin[0] blk.column\[0\].row\[12\].yc/lin[1]
+ blk.column\[1\].row\[12\].yc/uempty blk.column\[1\].row\[12\].yc/uin[0] blk.column\[1\].row\[12\].yc/uin[1]
+ blk.column\[1\].row\[11\].yc/din[0] blk.column\[1\].row\[11\].yc/din[1] blk.column\[1\].row\[11\].yc/dempty
+ blk.column\[1\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_81_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_489_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_437_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_702_ VGND VGND VPWR VPWR _702_/HI la_data_out[86] sky130_fd_sc_hd__conb_1
XPHY_7077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_633_ VGND VGND VPWR VPWR _633_/HI io_out[7] sky130_fd_sc_hd__conb_1
XPHY_5642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_564_ VGND VGND VPWR VPWR _564_/HI _564_/LO sky130_fd_sc_hd__conb_1
XPHY_4963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_460_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_495_ VGND VGND VPWR VPWR _495_/HI _495_/LO sky130_fd_sc_hd__conb_1
XFILLER_377_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_346_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_507_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_541_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_517_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_527_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_442_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_538_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_198_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_495_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_212_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_504_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_512_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_308_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_440_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_616_ VGND VGND VPWR VPWR _616_/HI io_oeb[28] sky130_fd_sc_hd__conb_1
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_398_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_547_ VGND VGND VPWR VPWR _547_/HI _547_/LO sky130_fd_sc_hd__conb_1
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_232_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_294_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_478_ VGND VGND VPWR VPWR _478_/HI _478_/LO sky130_fd_sc_hd__conb_1
XFILLER_439_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_255_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_536_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_448_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_465_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_528_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_352_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_273_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_403_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_401_ _398_/X wbs_dat_o[18] _786_/Q _396_/X VGND VGND VPWR VPWR _762_/D sky130_fd_sc_hd__o22a_4
XFILLER_15_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_540_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_332_ _330_/Y _331_/X wbs_dat_i[10] _331_/X VGND VGND VPWR VPWR _332_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_517_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_358_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[4\].yc blk.column\[10\].row\[4\].yc/cbitin blk.column\[10\].row\[5\].yc/cbitin
+ blk.column\[10\].row\[4\].yc/confclk blk.column\[10\].row\[5\].yc/confclk blk.column\[10\].row\[4\].yc/dempty
+ blk.column\[10\].row\[4\].yc/din[0] blk.column\[10\].row\[4\].yc/din[1] blk.column\[10\].row\[5\].yc/uin[0]
+ blk.column\[10\].row\[5\].yc/uin[1] blk.column\[10\].row\[4\].yc/hempty blk.column\[9\].row\[4\].yc/lempty
+ blk.column\[10\].row\[4\].yc/lempty blk.column\[10\].row\[4\].yc/lin[0] blk.column\[10\].row\[4\].yc/lin[1]
+ blk.column\[11\].row\[4\].yc/rin[0] blk.column\[11\].row\[4\].yc/rin[1] blk.column\[9\].row\[4\].yc/hempty
+ blk.column\[10\].row\[4\].yc/reset blk.column\[10\].row\[5\].yc/reset blk.column\[9\].row\[4\].yc/lout[0]
+ blk.column\[9\].row\[4\].yc/lout[1] blk.column\[9\].row\[4\].yc/lin[0] blk.column\[9\].row\[4\].yc/lin[1]
+ blk.column\[10\].row\[4\].yc/uempty blk.column\[10\].row\[4\].yc/uin[0] blk.column\[10\].row\[4\].yc/uin[1]
+ blk.column\[10\].row\[3\].yc/din[0] blk.column\[10\].row\[3\].yc/din[1] blk.column\[10\].row\[3\].yc/dempty
+ blk.column\[10\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_178_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_534_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_497_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_365_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[5\].yc blk.column\[1\].row\[5\].yc/cbitin blk.column\[1\].row\[6\].yc/cbitin
+ blk.column\[1\].row\[5\].yc/confclk blk.column\[1\].row\[6\].yc/confclk blk.column\[1\].row\[5\].yc/dempty
+ blk.column\[1\].row\[5\].yc/din[0] blk.column\[1\].row\[5\].yc/din[1] blk.column\[1\].row\[6\].yc/uin[0]
+ blk.column\[1\].row\[6\].yc/uin[1] blk.column\[1\].row\[5\].yc/hempty blk.column\[0\].row\[5\].yc/lempty
+ blk.column\[1\].row\[5\].yc/lempty blk.column\[1\].row\[5\].yc/lin[0] blk.column\[1\].row\[5\].yc/lin[1]
+ blk.column\[2\].row\[5\].yc/rin[0] blk.column\[2\].row\[5\].yc/rin[1] blk.column\[0\].row\[5\].yc/hempty
+ blk.column\[1\].row\[5\].yc/reset blk.column\[1\].row\[6\].yc/reset blk.column\[1\].row\[5\].yc/rin[0]
+ blk.column\[1\].row\[5\].yc/rin[1] blk.column\[0\].row\[5\].yc/lin[0] blk.column\[0\].row\[5\].yc/lin[1]
+ blk.column\[1\].row\[5\].yc/uempty blk.column\[1\].row\[5\].yc/uin[0] blk.column\[1\].row\[5\].yc/uin[1]
+ blk.column\[1\].row\[4\].yc/din[0] blk.column\[1\].row\[4\].yc/din[1] blk.column\[1\].row\[4\].yc/dempty
+ blk.column\[1\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_482_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[15\].yc blk.column\[5\].row\[15\].yc/cbitin la_data_out[37]
+ blk.column\[5\].row\[15\].yc/confclk blk.column\[5\].row\[15\].yc/confclko _471_/HI
+ _574_/LO _575_/LO blk.column\[5\].row\[15\].yc/dout[0] blk.column\[5\].row\[15\].yc/dout[1]
+ blk.column\[5\].row\[15\].yc/hempty blk.column\[4\].row\[15\].yc/lempty blk.column\[5\].row\[15\].yc/lempty
+ blk.column\[5\].row\[15\].yc/lin[0] blk.column\[5\].row\[15\].yc/lin[1] blk.column\[6\].row\[15\].yc/rin[0]
+ blk.column\[6\].row\[15\].yc/rin[1] blk.column\[4\].row\[15\].yc/hempty blk.column\[5\].row\[15\].yc/reset
+ blk.column\[5\].row\[15\].yc/reseto blk.column\[5\].row\[15\].yc/rin[0] blk.column\[5\].row\[15\].yc/rin[1]
+ blk.column\[4\].row\[15\].yc/lin[0] blk.column\[4\].row\[15\].yc/lin[1] blk.column\[5\].row\[15\].yc/uempty
+ blk.column\[5\].row\[15\].yc/uin[0] blk.column\[5\].row\[15\].yc/uin[1] blk.column\[5\].row\[14\].yc/din[0]
+ blk.column\[5\].row\[14\].yc/din[1] blk.column\[5\].row\[14\].yc/dempty blk.column\[5\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_101_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_429_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_481_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_498_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_355_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_499_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_325_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_535_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_274_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_429_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_362_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_542_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_315_ _314_/Y _310_/X wbs_dat_i[0] _298_/A VGND VGND VPWR VPWR _800_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_455_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_385_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_11160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_385_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1046 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_313_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_795_ wb_clk_i _795_/D VGND VGND VPWR VPWR _795_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_542_2226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_483_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_520_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_536_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_536_2019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_493_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_487_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_460_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_213_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_367_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_419_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_274_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_255_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_489_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_580_ VGND VGND VPWR VPWR _580_/HI _580_/LO sky130_fd_sc_hd__conb_1
XFILLER_483_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_341_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xblk.column\[11\].row\[6\].yc blk.column\[11\].row\[6\].yc/cbitin blk.column\[11\].row\[7\].yc/cbitin
+ blk.column\[11\].row\[6\].yc/confclk blk.column\[11\].row\[7\].yc/confclk blk.column\[11\].row\[6\].yc/dempty
+ blk.column\[11\].row\[6\].yc/din[0] blk.column\[11\].row\[6\].yc/din[1] blk.column\[11\].row\[7\].yc/uin[0]
+ blk.column\[11\].row\[7\].yc/uin[1] blk.column\[11\].row\[6\].yc/hempty blk.column\[10\].row\[6\].yc/lempty
+ blk.column\[11\].row\[6\].yc/lempty blk.column\[11\].row\[6\].yc/lin[0] blk.column\[11\].row\[6\].yc/lin[1]
+ blk.column\[12\].row\[6\].yc/rin[0] blk.column\[12\].row\[6\].yc/rin[1] blk.column\[10\].row\[6\].yc/hempty
+ blk.column\[11\].row\[6\].yc/reset blk.column\[11\].row\[7\].yc/reset blk.column\[11\].row\[6\].yc/rin[0]
+ blk.column\[11\].row\[6\].yc/rin[1] blk.column\[10\].row\[6\].yc/lin[0] blk.column\[10\].row\[6\].yc/lin[1]
+ blk.column\[11\].row\[6\].yc/uempty blk.column\[11\].row\[6\].yc/uin[0] blk.column\[11\].row\[6\].yc/uin[1]
+ blk.column\[11\].row\[5\].yc/din[0] blk.column\[11\].row\[5\].yc/din[1] blk.column\[11\].row\[5\].yc/dempty
+ blk.column\[11\].row\[7\].yc/uempty VPWR VGND ycell
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_437_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_385_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[7\].yc blk.column\[2\].row\[7\].yc/cbitin blk.column\[2\].row\[8\].yc/cbitin
+ blk.column\[2\].row\[7\].yc/confclk blk.column\[2\].row\[8\].yc/confclk blk.column\[2\].row\[7\].yc/dempty
+ blk.column\[2\].row\[7\].yc/din[0] blk.column\[2\].row\[7\].yc/din[1] blk.column\[2\].row\[8\].yc/uin[0]
+ blk.column\[2\].row\[8\].yc/uin[1] blk.column\[2\].row\[7\].yc/hempty blk.column\[1\].row\[7\].yc/lempty
+ blk.column\[2\].row\[7\].yc/lempty blk.column\[2\].row\[7\].yc/lin[0] blk.column\[2\].row\[7\].yc/lin[1]
+ blk.column\[3\].row\[7\].yc/rin[0] blk.column\[3\].row\[7\].yc/rin[1] blk.column\[1\].row\[7\].yc/hempty
+ blk.column\[2\].row\[7\].yc/reset blk.column\[2\].row\[8\].yc/reset blk.column\[2\].row\[7\].yc/rin[0]
+ blk.column\[2\].row\[7\].yc/rin[1] blk.column\[1\].row\[7\].yc/lin[0] blk.column\[1\].row\[7\].yc/lin[1]
+ blk.column\[2\].row\[7\].yc/uempty blk.column\[2\].row\[7\].yc/uin[0] blk.column\[2\].row\[7\].yc/uin[1]
+ blk.column\[2\].row\[6\].yc/din[0] blk.column\[2\].row\[6\].yc/din[1] blk.column\[2\].row\[6\].yc/dempty
+ blk.column\[2\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_10_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[10\].yc blk.column\[7\].row\[9\].yc/cbitout blk.column\[7\].row\[11\].yc/cbitin
+ blk.column\[7\].row\[9\].yc/confclko blk.column\[7\].row\[11\].yc/confclk blk.column\[7\].row\[10\].yc/dempty
+ blk.column\[7\].row\[10\].yc/din[0] blk.column\[7\].row\[10\].yc/din[1] blk.column\[7\].row\[11\].yc/uin[0]
+ blk.column\[7\].row\[11\].yc/uin[1] blk.column\[7\].row\[10\].yc/hempty blk.column\[6\].row\[10\].yc/lempty
+ blk.column\[7\].row\[10\].yc/lempty blk.column\[7\].row\[10\].yc/lin[0] blk.column\[7\].row\[10\].yc/lin[1]
+ blk.column\[8\].row\[10\].yc/rin[0] blk.column\[8\].row\[10\].yc/rin[1] blk.column\[6\].row\[10\].yc/hempty
+ blk.column\[7\].row\[9\].yc/reseto blk.column\[7\].row\[11\].yc/reset blk.column\[7\].row\[10\].yc/rin[0]
+ blk.column\[7\].row\[10\].yc/rin[1] blk.column\[6\].row\[10\].yc/lin[0] blk.column\[6\].row\[10\].yc/lin[1]
+ blk.column\[7\].row\[9\].yc/vempty2 blk.column\[7\].row\[9\].yc/dout[0] blk.column\[7\].row\[9\].yc/dout[1]
+ blk.column\[7\].row\[9\].yc/din[0] blk.column\[7\].row\[9\].yc/din[1] blk.column\[7\].row\[9\].yc/dempty
+ blk.column\[7\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_23_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_239_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_254_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_778_ wb_clk_i _778_/D VGND VGND VPWR VPWR _778_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_520_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_499_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_449_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_367_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_371_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_323_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[1\].yc blk.column\[7\].row\[1\].yc/cbitin blk.column\[7\].row\[2\].yc/cbitin
+ blk.column\[7\].row\[1\].yc/confclk blk.column\[7\].row\[2\].yc/confclk blk.column\[7\].row\[1\].yc/dempty
+ blk.column\[7\].row\[1\].yc/din[0] blk.column\[7\].row\[1\].yc/din[1] blk.column\[7\].row\[2\].yc/uin[0]
+ blk.column\[7\].row\[2\].yc/uin[1] blk.column\[7\].row\[1\].yc/hempty blk.column\[6\].row\[1\].yc/lempty
+ blk.column\[7\].row\[1\].yc/lempty blk.column\[7\].row\[1\].yc/lin[0] blk.column\[7\].row\[1\].yc/lin[1]
+ blk.column\[8\].row\[1\].yc/rin[0] blk.column\[8\].row\[1\].yc/rin[1] blk.column\[6\].row\[1\].yc/hempty
+ blk.column\[7\].row\[1\].yc/reset blk.column\[7\].row\[2\].yc/reset blk.column\[7\].row\[1\].yc/rin[0]
+ blk.column\[7\].row\[1\].yc/rin[1] blk.column\[6\].row\[1\].yc/lin[0] blk.column\[6\].row\[1\].yc/lin[1]
+ blk.column\[7\].row\[1\].yc/uempty blk.column\[7\].row\[1\].yc/uin[0] blk.column\[7\].row\[1\].yc/uin[1]
+ blk.column\[7\].row\[0\].yc/din[0] blk.column\[7\].row\[0\].yc/din[1] blk.column\[7\].row\[0\].yc/dempty
+ blk.column\[7\].row\[2\].yc/uempty VPWR VGND ycell
XPHY_7034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_701_ VGND VGND VPWR VPWR _701_/HI la_data_out[85] sky130_fd_sc_hd__conb_1
XPHY_7067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_236_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_632_ VGND VGND VPWR VPWR _632_/HI io_out[6] sky130_fd_sc_hd__conb_1
XPHY_6366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_563_ VGND VGND VPWR VPWR _563_/HI _563_/LO sky130_fd_sc_hd__conb_1
XPHY_5676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_494_ VGND VGND VPWR VPWR _494_/HI _494_/LO sky130_fd_sc_hd__conb_1
XFILLER_521_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_400_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_515_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_507_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_504_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_515_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_428_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_264_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_522_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_520_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_305_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_312_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_243_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[12\].yc blk.column\[14\].row\[12\].yc/cbitin blk.column\[14\].row\[13\].yc/cbitin
+ blk.column\[14\].row\[12\].yc/confclk blk.column\[14\].row\[13\].yc/confclk blk.column\[14\].row\[12\].yc/dempty
+ blk.column\[14\].row\[12\].yc/din[0] blk.column\[14\].row\[12\].yc/din[1] blk.column\[14\].row\[13\].yc/uin[0]
+ blk.column\[14\].row\[13\].yc/uin[1] blk.column\[14\].row\[12\].yc/hempty blk.column\[13\].row\[12\].yc/lempty
+ blk.column\[14\].row\[12\].yc/lempty blk.column\[14\].row\[12\].yc/lin[0] blk.column\[14\].row\[12\].yc/lin[1]
+ blk.column\[15\].row\[12\].yc/rin[0] blk.column\[15\].row\[12\].yc/rin[1] blk.column\[13\].row\[12\].yc/hempty
+ blk.column\[14\].row\[12\].yc/reset blk.column\[14\].row\[13\].yc/reset blk.column\[14\].row\[12\].yc/rin[0]
+ blk.column\[14\].row\[12\].yc/rin[1] blk.column\[13\].row\[12\].yc/lin[0] blk.column\[13\].row\[12\].yc/lin[1]
+ blk.column\[14\].row\[12\].yc/uempty blk.column\[14\].row\[12\].yc/uin[0] blk.column\[14\].row\[12\].yc/uin[1]
+ blk.column\[14\].row\[11\].yc/din[0] blk.column\[14\].row\[11\].yc/din[1] blk.column\[14\].row\[11\].yc/dempty
+ blk.column\[14\].row\[13\].yc/uempty VPWR VGND ycell
XPHY_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_497_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_485_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_287_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_10833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_10844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_308_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_615_ VGND VGND VPWR VPWR _615_/HI io_oeb[27] sky130_fd_sc_hd__conb_1
XPHY_6196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_5484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_546_ VGND VGND VPWR VPWR _546_/HI _546_/LO sky130_fd_sc_hd__conb_1
XFILLER_109_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_539_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_477_ VGND VGND VPWR VPWR _477_/HI _477_/LO sky130_fd_sc_hd__conb_1
XFILLER_536_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_521_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_335_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_250_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_353_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[8\].yc blk.column\[12\].row\[8\].yc/cbitin blk.column\[12\].row\[9\].yc/cbitin
+ blk.column\[12\].row\[8\].yc/confclk blk.column\[12\].row\[9\].yc/confclk blk.column\[12\].row\[8\].yc/dempty
+ blk.column\[12\].row\[8\].yc/din[0] blk.column\[12\].row\[8\].yc/din[1] blk.column\[12\].row\[9\].yc/uin[0]
+ blk.column\[12\].row\[9\].yc/uin[1] blk.column\[12\].row\[8\].yc/hempty blk.column\[11\].row\[8\].yc/lempty
+ blk.column\[12\].row\[8\].yc/lempty blk.column\[12\].row\[8\].yc/lin[0] blk.column\[12\].row\[8\].yc/lin[1]
+ blk.column\[13\].row\[8\].yc/rin[0] blk.column\[13\].row\[8\].yc/rin[1] blk.column\[11\].row\[8\].yc/hempty
+ blk.column\[12\].row\[8\].yc/reset blk.column\[12\].row\[9\].yc/reset blk.column\[12\].row\[8\].yc/rin[0]
+ blk.column\[12\].row\[8\].yc/rin[1] blk.column\[11\].row\[8\].yc/lin[0] blk.column\[11\].row\[8\].yc/lin[1]
+ blk.column\[12\].row\[8\].yc/uempty blk.column\[12\].row\[8\].yc/uin[0] blk.column\[12\].row\[8\].yc/uin[1]
+ blk.column\[12\].row\[7\].yc/din[0] blk.column\[12\].row\[7\].yc/din[1] blk.column\[12\].row\[7\].yc/dempty
+ blk.column\[12\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_505_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_407_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_400_ _398_/X wbs_dat_o[19] _349_/A _396_/X VGND VGND VPWR VPWR _400_/X sky130_fd_sc_hd__o22a_4
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_403_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_475_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ _319_/A VGND VGND VPWR VPWR _331_/X sky130_fd_sc_hd__buf_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_401_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_397_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_521_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xblk.column\[3\].row\[9\].yc blk.column\[3\].row\[9\].yc/cbitin blk.column\[3\].row\[9\].yc/cbitout
+ blk.column\[3\].row\[9\].yc/confclk blk.column\[3\].row\[9\].yc/confclko blk.column\[3\].row\[9\].yc/dempty
+ blk.column\[3\].row\[9\].yc/din[0] blk.column\[3\].row\[9\].yc/din[1] blk.column\[3\].row\[9\].yc/dout[0]
+ blk.column\[3\].row\[9\].yc/dout[1] blk.column\[3\].row\[9\].yc/hempty blk.column\[2\].row\[9\].yc/lempty
+ blk.column\[3\].row\[9\].yc/lempty blk.column\[3\].row\[9\].yc/lin[0] blk.column\[3\].row\[9\].yc/lin[1]
+ blk.column\[4\].row\[9\].yc/rin[0] blk.column\[4\].row\[9\].yc/rin[1] blk.column\[2\].row\[9\].yc/hempty
+ blk.column\[3\].row\[9\].yc/reset blk.column\[3\].row\[9\].yc/reseto blk.column\[3\].row\[9\].yc/rin[0]
+ blk.column\[3\].row\[9\].yc/rin[1] blk.column\[2\].row\[9\].yc/lin[0] blk.column\[2\].row\[9\].yc/lin[1]
+ blk.column\[3\].row\[9\].yc/uempty blk.column\[3\].row\[9\].yc/uin[0] blk.column\[3\].row\[9\].yc/uin[1]
+ blk.column\[3\].row\[8\].yc/din[0] blk.column\[3\].row\[8\].yc/din[1] blk.column\[3\].row\[8\].yc/dempty
+ blk.column\[3\].row\[9\].yc/vempty2 VPWR VGND ycell
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_532_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_383_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_482_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_482_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_529_ VGND VGND VPWR VPWR _529_/HI _529_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_536_2927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_337_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_508_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_506_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_270_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_522_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[3\].yc blk.column\[8\].row\[3\].yc/cbitin blk.column\[8\].row\[4\].yc/cbitin
+ blk.column\[8\].row\[3\].yc/confclk blk.column\[8\].row\[4\].yc/confclk blk.column\[8\].row\[3\].yc/dempty
+ blk.column\[8\].row\[3\].yc/din[0] blk.column\[8\].row\[3\].yc/din[1] blk.column\[8\].row\[4\].yc/uin[0]
+ blk.column\[8\].row\[4\].yc/uin[1] blk.column\[8\].row\[3\].yc/hempty blk.column\[7\].row\[3\].yc/lempty
+ blk.column\[8\].row\[3\].yc/lempty blk.column\[8\].row\[3\].yc/lin[0] blk.column\[8\].row\[3\].yc/lin[1]
+ blk.column\[9\].row\[3\].yc/rin[0] blk.column\[9\].row\[3\].yc/rin[1] blk.column\[7\].row\[3\].yc/hempty
+ blk.column\[8\].row\[3\].yc/reset blk.column\[8\].row\[4\].yc/reset blk.column\[8\].row\[3\].yc/rin[0]
+ blk.column\[8\].row\[3\].yc/rin[1] blk.column\[7\].row\[3\].yc/lin[0] blk.column\[7\].row\[3\].yc/lin[1]
+ blk.column\[8\].row\[3\].yc/uempty blk.column\[8\].row\[3\].yc/uin[0] blk.column\[8\].row\[3\].yc/uin[1]
+ blk.column\[8\].row\[2\].yc/din[0] blk.column\[8\].row\[2\].yc/din[1] blk.column\[8\].row\[2\].yc/dempty
+ blk.column\[8\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_10_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_429_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_362_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_272_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_497_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ _314_/A VGND VGND VPWR VPWR _314_/Y sky130_fd_sc_hd__inv_2
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_436_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[11\].yc blk.column\[2\].row\[11\].yc/cbitin blk.column\[2\].row\[12\].yc/cbitin
+ blk.column\[2\].row\[11\].yc/confclk blk.column\[2\].row\[12\].yc/confclk blk.column\[2\].row\[11\].yc/dempty
+ blk.column\[2\].row\[11\].yc/din[0] blk.column\[2\].row\[11\].yc/din[1] blk.column\[2\].row\[12\].yc/uin[0]
+ blk.column\[2\].row\[12\].yc/uin[1] blk.column\[2\].row\[11\].yc/hempty blk.column\[1\].row\[11\].yc/lempty
+ blk.column\[2\].row\[11\].yc/lempty blk.column\[2\].row\[11\].yc/lin[0] blk.column\[2\].row\[11\].yc/lin[1]
+ blk.column\[3\].row\[11\].yc/rin[0] blk.column\[3\].row\[11\].yc/rin[1] blk.column\[1\].row\[11\].yc/hempty
+ blk.column\[2\].row\[11\].yc/reset blk.column\[2\].row\[12\].yc/reset blk.column\[2\].row\[11\].yc/rin[0]
+ blk.column\[2\].row\[11\].yc/rin[1] blk.column\[1\].row\[11\].yc/lin[0] blk.column\[1\].row\[11\].yc/lin[1]
+ blk.column\[2\].row\[11\].yc/uempty blk.column\[2\].row\[11\].yc/uin[0] blk.column\[2\].row\[11\].yc/uin[1]
+ blk.column\[2\].row\[10\].yc/din[0] blk.column\[2\].row\[10\].yc/din[1] blk.column\[2\].row\[10\].yc/dempty
+ blk.column\[2\].row\[12\].yc/uempty VPWR VGND ycell
XPHY_1784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_256_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_324_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_541_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_487_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_528_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_419_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_435_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_327_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_451_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_451_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_794_ wb_clk_i _332_/X VGND VGND VPWR VPWR _330_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_21_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_258_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_514_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_488_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_432_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_540_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_358_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_231_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_472_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_235_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_777_ wb_clk_i _777_/D VGND VGND VPWR VPWR _375_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_526_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_501_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_518_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_522_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_289_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[5\].yc blk.column\[9\].row\[5\].yc/cbitin blk.column\[9\].row\[6\].yc/cbitin
+ blk.column\[9\].row\[5\].yc/confclk blk.column\[9\].row\[6\].yc/confclk blk.column\[9\].row\[5\].yc/dempty
+ blk.column\[9\].row\[5\].yc/din[0] blk.column\[9\].row\[5\].yc/din[1] blk.column\[9\].row\[6\].yc/uin[0]
+ blk.column\[9\].row\[6\].yc/uin[1] blk.column\[9\].row\[5\].yc/hempty blk.column\[8\].row\[5\].yc/lempty
+ blk.column\[9\].row\[5\].yc/lempty blk.column\[9\].row\[5\].yc/lin[0] blk.column\[9\].row\[5\].yc/lin[1]
+ blk.column\[9\].row\[5\].yc/lout[0] blk.column\[9\].row\[5\].yc/lout[1] blk.column\[8\].row\[5\].yc/hempty
+ blk.column\[9\].row\[5\].yc/reset blk.column\[9\].row\[6\].yc/reset blk.column\[9\].row\[5\].yc/rin[0]
+ blk.column\[9\].row\[5\].yc/rin[1] blk.column\[8\].row\[5\].yc/lin[0] blk.column\[8\].row\[5\].yc/lin[1]
+ blk.column\[9\].row\[5\].yc/uempty blk.column\[9\].row\[5\].yc/uin[0] blk.column\[9\].row\[5\].yc/uin[1]
+ blk.column\[9\].row\[4\].yc/din[0] blk.column\[9\].row\[4\].yc/din[1] blk.column\[9\].row\[4\].yc/dempty
+ blk.column\[9\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_206_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_516_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_432_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[6\].row\[14\].yc blk.column\[6\].row\[14\].yc/cbitin blk.column\[6\].row\[15\].yc/cbitin
+ blk.column\[6\].row\[14\].yc/confclk blk.column\[6\].row\[15\].yc/confclk blk.column\[6\].row\[14\].yc/dempty
+ blk.column\[6\].row\[14\].yc/din[0] blk.column\[6\].row\[14\].yc/din[1] blk.column\[6\].row\[15\].yc/uin[0]
+ blk.column\[6\].row\[15\].yc/uin[1] blk.column\[6\].row\[14\].yc/hempty blk.column\[5\].row\[14\].yc/lempty
+ blk.column\[6\].row\[14\].yc/lempty blk.column\[6\].row\[14\].yc/lin[0] blk.column\[6\].row\[14\].yc/lin[1]
+ blk.column\[7\].row\[14\].yc/rin[0] blk.column\[7\].row\[14\].yc/rin[1] blk.column\[5\].row\[14\].yc/hempty
+ blk.column\[6\].row\[14\].yc/reset blk.column\[6\].row\[15\].yc/reset blk.column\[6\].row\[14\].yc/rin[0]
+ blk.column\[6\].row\[14\].yc/rin[1] blk.column\[5\].row\[14\].yc/lin[0] blk.column\[5\].row\[14\].yc/lin[1]
+ blk.column\[6\].row\[14\].yc/uempty blk.column\[6\].row\[14\].yc/uin[0] blk.column\[6\].row\[14\].yc/uin[1]
+ blk.column\[6\].row\[13\].yc/din[0] blk.column\[6\].row\[13\].yc/din[1] blk.column\[6\].row\[13\].yc/dempty
+ blk.column\[6\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_7_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_700_ VGND VGND VPWR VPWR _700_/HI la_data_out[84] sky130_fd_sc_hd__conb_1
XPHY_7057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_631_ VGND VGND VPWR VPWR _631_/HI io_out[5] sky130_fd_sc_hd__conb_1
XPHY_6367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_562_ VGND VGND VPWR VPWR _562_/HI _562_/LO sky130_fd_sc_hd__conb_1
XPHY_5666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_352_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_493_ VGND VGND VPWR VPWR _493_/HI _493_/LO sky130_fd_sc_hd__conb_1
XFILLER_496_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_401_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_537_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_522_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_520_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_522_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_531_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_533_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_393_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_614_ VGND VGND VPWR VPWR _614_/HI io_oeb[26] sky130_fd_sc_hd__conb_1
XPHY_5452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_308_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_5463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_545_ VGND VGND VPWR VPWR _545_/HI _545_/LO sky130_fd_sc_hd__conb_1
XFILLER_504_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_476_ VGND VGND VPWR VPWR _476_/HI _476_/LO sky130_fd_sc_hd__conb_1
XFILLER_517_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_319_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_259_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_247_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_360_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_521_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_403_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_330_ _330_/A VGND VGND VPWR VPWR _330_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_540_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_319_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_288_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_254_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_438_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_384_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_399_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_252_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_528_ VGND VGND VPWR VPWR _528_/HI _528_/LO sky130_fd_sc_hd__conb_1
XFILLER_220_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_459_ VGND VGND VPWR VPWR _459_/HI _459_/LO sky130_fd_sc_hd__conb_1
XFILLER_536_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_302_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_337_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_500_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_522_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_277_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_408_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_251_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_435_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_344_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_403_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ _312_/Y _310_/X wbs_dat_i[1] _310_/X VGND VGND VPWR VPWR _313_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_475_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_348_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_295_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_436_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_505_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[6\].yc blk.column\[0\].row\[6\].yc/cbitin blk.column\[0\].row\[7\].yc/cbitin
+ blk.column\[0\].row\[6\].yc/confclk blk.column\[0\].row\[7\].yc/confclk blk.column\[0\].row\[6\].yc/dempty
+ blk.column\[0\].row\[6\].yc/din[0] blk.column\[0\].row\[6\].yc/din[1] blk.column\[0\].row\[7\].yc/uin[0]
+ blk.column\[0\].row\[7\].yc/uin[1] blk.column\[0\].row\[6\].yc/hempty blk.column\[0\].row\[6\].yc/hempty2
+ blk.column\[0\].row\[6\].yc/lempty blk.column\[0\].row\[6\].yc/lin[0] blk.column\[0\].row\[6\].yc/lin[1]
+ blk.column\[1\].row\[6\].yc/rin[0] blk.column\[1\].row\[6\].yc/rin[1] _441_/HI blk.column\[0\].row\[6\].yc/reset
+ blk.column\[0\].row\[7\].yc/reset _503_/LO _504_/LO blk.column\[0\].row\[6\].yc/rout[0]
+ blk.column\[0\].row\[6\].yc/rout[1] blk.column\[0\].row\[6\].yc/uempty blk.column\[0\].row\[6\].yc/uin[0]
+ blk.column\[0\].row\[6\].yc/uin[1] blk.column\[0\].row\[5\].yc/din[0] blk.column\[0\].row\[5\].yc/din[1]
+ blk.column\[0\].row\[5\].yc/dempty blk.column\[0\].row\[7\].yc/uempty VPWR VGND
+ ycell
XPHY_5090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_419_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_228_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_476_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_432_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_269_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_486_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_269_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_385_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_528_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[15\].yc blk.column\[1\].row\[15\].yc/cbitin la_data_out[33]
+ blk.column\[1\].row\[15\].yc/confclk blk.column\[1\].row\[15\].yc/confclko _467_/HI
+ _562_/LO _563_/LO blk.column\[1\].row\[15\].yc/dout[0] blk.column\[1\].row\[15\].yc/dout[1]
+ blk.column\[1\].row\[15\].yc/hempty blk.column\[0\].row\[15\].yc/lempty blk.column\[1\].row\[15\].yc/lempty
+ blk.column\[1\].row\[15\].yc/lin[0] blk.column\[1\].row\[15\].yc/lin[1] blk.column\[2\].row\[15\].yc/rin[0]
+ blk.column\[2\].row\[15\].yc/rin[1] blk.column\[0\].row\[15\].yc/hempty blk.column\[1\].row\[15\].yc/reset
+ blk.column\[1\].row\[15\].yc/reseto blk.column\[1\].row\[15\].yc/rin[0] blk.column\[1\].row\[15\].yc/rin[1]
+ blk.column\[0\].row\[15\].yc/lin[0] blk.column\[0\].row\[15\].yc/lin[1] blk.column\[1\].row\[15\].yc/uempty
+ blk.column\[1\].row\[15\].yc/uin[0] blk.column\[1\].row\[15\].yc/uin[1] blk.column\[1\].row\[14\].yc/din[0]
+ blk.column\[1\].row\[14\].yc/din[1] blk.column\[1\].row\[14\].yc/dempty blk.column\[1\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_10_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_542_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_270_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_435_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_327_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_281_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_793_ wb_clk_i _334_/X VGND VGND VPWR VPWR _333_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_112_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_451_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[15\].row\[11\].yc blk.column\[15\].row\[11\].yc/cbitin blk.column\[15\].row\[12\].yc/cbitin
+ blk.column\[15\].row\[11\].yc/confclk blk.column\[15\].row\[12\].yc/confclk blk.column\[15\].row\[11\].yc/dempty
+ blk.column\[15\].row\[11\].yc/din[0] blk.column\[15\].row\[11\].yc/din[1] blk.column\[15\].row\[12\].yc/uin[0]
+ blk.column\[15\].row\[12\].yc/uin[1] blk.column\[15\].row\[11\].yc/hempty blk.column\[14\].row\[11\].yc/lempty
+ _452_/HI _531_/LO _532_/LO blk.column\[15\].row\[11\].yc/lout[0] blk.column\[15\].row\[11\].yc/lout[1]
+ blk.column\[14\].row\[11\].yc/hempty blk.column\[15\].row\[11\].yc/reset blk.column\[15\].row\[12\].yc/reset
+ blk.column\[15\].row\[11\].yc/rin[0] blk.column\[15\].row\[11\].yc/rin[1] blk.column\[14\].row\[11\].yc/lin[0]
+ blk.column\[14\].row\[11\].yc/lin[1] blk.column\[15\].row\[11\].yc/uempty blk.column\[15\].row\[11\].yc/uin[0]
+ blk.column\[15\].row\[11\].yc/uin[1] blk.column\[15\].row\[10\].yc/din[0] blk.column\[15\].row\[10\].yc/din[1]
+ blk.column\[15\].row\[10\].yc/dempty blk.column\[15\].row\[12\].yc/uempty VPWR VGND
+ ycell
XFILLER_408_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_520_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[0\].yc la_data_in[101] blk.column\[5\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[5\].row\[1\].yc/confclk blk.column\[5\].row\[0\].yc/dempty blk.column\[5\].row\[0\].yc/din[0]
+ blk.column\[5\].row\[0\].yc/din[1] blk.column\[5\].row\[1\].yc/uin[0] blk.column\[5\].row\[1\].yc/uin[1]
+ blk.column\[5\].row\[0\].yc/hempty blk.column\[4\].row\[0\].yc/lempty blk.column\[5\].row\[0\].yc/lempty
+ blk.column\[5\].row\[0\].yc/lin[0] blk.column\[5\].row\[0\].yc/lin[1] blk.column\[6\].row\[0\].yc/rin[0]
+ blk.column\[6\].row\[0\].yc/rin[1] blk.column\[4\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[5\].row\[1\].yc/reset blk.column\[5\].row\[0\].yc/rin[0] blk.column\[5\].row\[0\].yc/rin[1]
+ blk.column\[4\].row\[0\].yc/lin[0] blk.column\[4\].row\[0\].yc/lin[1] _573_/LO la_data_in[74]
+ la_data_in[75] la_data_out[10] la_data_out[11] blk.column\[5\].row\[0\].yc/vempty
+ blk.column\[5\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_179_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_501_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_476_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_512_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_361_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_225_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_367_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_536_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_315_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_246_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_472_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_358_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_476_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_535_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_531_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_8485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_470_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_776_ wb_clk_i _378_/X VGND VGND VPWR VPWR _776_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2047 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_496_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_297_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_364_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_502_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_505_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_504_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_630_ VGND VGND VPWR VPWR _630_/HI io_out[4] sky130_fd_sc_hd__conb_1
XPHY_6346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_561_ VGND VGND VPWR VPWR _561_/HI _561_/LO sky130_fd_sc_hd__conb_1
XFILLER_508_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_492_ VGND VGND VPWR VPWR _492_/HI _492_/LO sky130_fd_sc_hd__conb_1
XFILLER_2_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_345_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[7\].yc blk.column\[10\].row\[7\].yc/cbitin blk.column\[10\].row\[8\].yc/cbitin
+ blk.column\[10\].row\[7\].yc/confclk blk.column\[10\].row\[8\].yc/confclk blk.column\[10\].row\[7\].yc/dempty
+ blk.column\[10\].row\[7\].yc/din[0] blk.column\[10\].row\[7\].yc/din[1] blk.column\[10\].row\[8\].yc/uin[0]
+ blk.column\[10\].row\[8\].yc/uin[1] blk.column\[10\].row\[7\].yc/hempty blk.column\[9\].row\[7\].yc/lempty
+ blk.column\[10\].row\[7\].yc/lempty blk.column\[10\].row\[7\].yc/lin[0] blk.column\[10\].row\[7\].yc/lin[1]
+ blk.column\[11\].row\[7\].yc/rin[0] blk.column\[11\].row\[7\].yc/rin[1] blk.column\[9\].row\[7\].yc/hempty
+ blk.column\[10\].row\[7\].yc/reset blk.column\[10\].row\[8\].yc/reset blk.column\[9\].row\[7\].yc/lout[0]
+ blk.column\[9\].row\[7\].yc/lout[1] blk.column\[9\].row\[7\].yc/lin[0] blk.column\[9\].row\[7\].yc/lin[1]
+ blk.column\[10\].row\[7\].yc/uempty blk.column\[10\].row\[7\].yc/uin[0] blk.column\[10\].row\[7\].yc/uin[1]
+ blk.column\[10\].row\[6\].yc/din[0] blk.column\[10\].row\[6\].yc/din[1] blk.column\[10\].row\[6\].yc/dempty
+ blk.column\[10\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_537_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_300_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_218_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[8\].yc blk.column\[1\].row\[8\].yc/cbitin blk.column\[1\].row\[9\].yc/cbitin
+ blk.column\[1\].row\[8\].yc/confclk blk.column\[1\].row\[9\].yc/confclk blk.column\[1\].row\[8\].yc/dempty
+ blk.column\[1\].row\[8\].yc/din[0] blk.column\[1\].row\[8\].yc/din[1] blk.column\[1\].row\[9\].yc/uin[0]
+ blk.column\[1\].row\[9\].yc/uin[1] blk.column\[1\].row\[8\].yc/hempty blk.column\[0\].row\[8\].yc/lempty
+ blk.column\[1\].row\[8\].yc/lempty blk.column\[1\].row\[8\].yc/lin[0] blk.column\[1\].row\[8\].yc/lin[1]
+ blk.column\[2\].row\[8\].yc/rin[0] blk.column\[2\].row\[8\].yc/rin[1] blk.column\[0\].row\[8\].yc/hempty
+ blk.column\[1\].row\[8\].yc/reset blk.column\[1\].row\[9\].yc/reset blk.column\[1\].row\[8\].yc/rin[0]
+ blk.column\[1\].row\[8\].yc/rin[1] blk.column\[0\].row\[8\].yc/lin[0] blk.column\[0\].row\[8\].yc/lin[1]
+ blk.column\[1\].row\[8\].yc/uempty blk.column\[1\].row\[8\].yc/uin[0] blk.column\[1\].row\[8\].yc/uin[1]
+ blk.column\[1\].row\[7\].yc/din[0] blk.column\[1\].row\[7\].yc/din[1] blk.column\[1\].row\[7\].yc/dempty
+ blk.column\[1\].row\[9\].yc/uempty VPWR VGND ycell
XPHY_8271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_759_ wb_clk_i _406_/X VGND VGND VPWR VPWR wbs_dat_o[15] sky130_fd_sc_hd__dfxtp_4
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_520_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[10\].yc blk.column\[3\].row\[9\].yc/cbitout blk.column\[3\].row\[11\].yc/cbitin
+ blk.column\[3\].row\[9\].yc/confclko blk.column\[3\].row\[11\].yc/confclk blk.column\[3\].row\[10\].yc/dempty
+ blk.column\[3\].row\[10\].yc/din[0] blk.column\[3\].row\[10\].yc/din[1] blk.column\[3\].row\[11\].yc/uin[0]
+ blk.column\[3\].row\[11\].yc/uin[1] blk.column\[3\].row\[10\].yc/hempty blk.column\[2\].row\[10\].yc/lempty
+ blk.column\[3\].row\[10\].yc/lempty blk.column\[3\].row\[10\].yc/lin[0] blk.column\[3\].row\[10\].yc/lin[1]
+ blk.column\[4\].row\[10\].yc/rin[0] blk.column\[4\].row\[10\].yc/rin[1] blk.column\[2\].row\[10\].yc/hempty
+ blk.column\[3\].row\[9\].yc/reseto blk.column\[3\].row\[11\].yc/reset blk.column\[3\].row\[10\].yc/rin[0]
+ blk.column\[3\].row\[10\].yc/rin[1] blk.column\[2\].row\[10\].yc/lin[0] blk.column\[2\].row\[10\].yc/lin[1]
+ blk.column\[3\].row\[9\].yc/vempty2 blk.column\[3\].row\[9\].yc/dout[0] blk.column\[3\].row\[9\].yc/dout[1]
+ blk.column\[3\].row\[9\].yc/din[0] blk.column\[3\].row\[9\].yc/din[1] blk.column\[3\].row\[9\].yc/dempty
+ blk.column\[3\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_195_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_367_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_434_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_277_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_519_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[1\].yc blk.column\[15\].row\[1\].yc/cbitin blk.column\[15\].row\[2\].yc/cbitin
+ blk.column\[15\].row\[1\].yc/confclk blk.column\[15\].row\[2\].yc/confclk blk.column\[15\].row\[1\].yc/dempty
+ blk.column\[15\].row\[1\].yc/din[0] blk.column\[15\].row\[1\].yc/din[1] blk.column\[15\].row\[2\].yc/uin[0]
+ blk.column\[15\].row\[2\].yc/uin[1] blk.column\[15\].row\[1\].yc/hempty blk.column\[14\].row\[1\].yc/lempty
+ _458_/HI _543_/LO _544_/LO blk.column\[15\].row\[1\].yc/lout[0] blk.column\[15\].row\[1\].yc/lout[1]
+ blk.column\[14\].row\[1\].yc/hempty blk.column\[15\].row\[1\].yc/reset blk.column\[15\].row\[2\].yc/reset
+ blk.column\[15\].row\[1\].yc/rin[0] blk.column\[15\].row\[1\].yc/rin[1] blk.column\[14\].row\[1\].yc/lin[0]
+ blk.column\[14\].row\[1\].yc/lin[1] blk.column\[15\].row\[1\].yc/uempty blk.column\[15\].row\[1\].yc/uin[0]
+ blk.column\[15\].row\[1\].yc/uin[1] blk.column\[15\].row\[0\].yc/din[0] blk.column\[15\].row\[0\].yc/din[1]
+ blk.column\[15\].row\[0\].yc/dempty blk.column\[15\].row\[2\].yc/uempty VPWR VGND
+ ycell
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[2\].yc blk.column\[6\].row\[2\].yc/cbitin blk.column\[6\].row\[3\].yc/cbitin
+ blk.column\[6\].row\[2\].yc/confclk blk.column\[6\].row\[3\].yc/confclk blk.column\[6\].row\[2\].yc/dempty
+ blk.column\[6\].row\[2\].yc/din[0] blk.column\[6\].row\[2\].yc/din[1] blk.column\[6\].row\[3\].yc/uin[0]
+ blk.column\[6\].row\[3\].yc/uin[1] blk.column\[6\].row\[2\].yc/hempty blk.column\[5\].row\[2\].yc/lempty
+ blk.column\[6\].row\[2\].yc/lempty blk.column\[6\].row\[2\].yc/lin[0] blk.column\[6\].row\[2\].yc/lin[1]
+ blk.column\[7\].row\[2\].yc/rin[0] blk.column\[7\].row\[2\].yc/rin[1] blk.column\[5\].row\[2\].yc/hempty
+ blk.column\[6\].row\[2\].yc/reset blk.column\[6\].row\[3\].yc/reset blk.column\[6\].row\[2\].yc/rin[0]
+ blk.column\[6\].row\[2\].yc/rin[1] blk.column\[5\].row\[2\].yc/lin[0] blk.column\[5\].row\[2\].yc/lin[1]
+ blk.column\[6\].row\[2\].yc/uempty blk.column\[6\].row\[2\].yc/uin[0] blk.column\[6\].row\[2\].yc/uin[1]
+ blk.column\[6\].row\[1\].yc/din[0] blk.column\[6\].row\[1\].yc/din[1] blk.column\[6\].row\[1\].yc/dempty
+ blk.column\[6\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_183_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_613_ VGND VGND VPWR VPWR _613_/HI io_oeb[25] sky130_fd_sc_hd__conb_1
XPHY_6176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_418_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_544_ VGND VGND VPWR VPWR _544_/HI _544_/LO sky130_fd_sc_hd__conb_1
XFILLER_521_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_378_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_475_ VGND VGND VPWR VPWR _475_/HI _475_/LO sky130_fd_sc_hd__conb_1
XPHY_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_478_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_298_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_521_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_534_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_416_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_522_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_508_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_439_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_521_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_430_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_475_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_319_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_377_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[12\].yc blk.column\[10\].row\[12\].yc/cbitin blk.column\[10\].row\[13\].yc/cbitin
+ blk.column\[10\].row\[12\].yc/confclk blk.column\[10\].row\[13\].yc/confclk blk.column\[10\].row\[12\].yc/dempty
+ blk.column\[10\].row\[12\].yc/din[0] blk.column\[10\].row\[12\].yc/din[1] blk.column\[10\].row\[13\].yc/uin[0]
+ blk.column\[10\].row\[13\].yc/uin[1] blk.column\[10\].row\[12\].yc/hempty blk.column\[9\].row\[12\].yc/lempty
+ blk.column\[10\].row\[12\].yc/lempty blk.column\[10\].row\[12\].yc/lin[0] blk.column\[10\].row\[12\].yc/lin[1]
+ blk.column\[11\].row\[12\].yc/rin[0] blk.column\[11\].row\[12\].yc/rin[1] blk.column\[9\].row\[12\].yc/hempty
+ blk.column\[10\].row\[12\].yc/reset blk.column\[10\].row\[13\].yc/reset blk.column\[9\].row\[12\].yc/lout[0]
+ blk.column\[9\].row\[12\].yc/lout[1] blk.column\[9\].row\[12\].yc/lin[0] blk.column\[9\].row\[12\].yc/lin[1]
+ blk.column\[10\].row\[12\].yc/uempty blk.column\[10\].row\[12\].yc/uin[0] blk.column\[10\].row\[12\].yc/uin[1]
+ blk.column\[10\].row\[11\].yc/din[0] blk.column\[10\].row\[11\].yc/din[1] blk.column\[10\].row\[11\].yc/dempty
+ blk.column\[10\].row\[13\].yc/uempty VPWR VGND ycell
XPHY_11300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_527_ VGND VGND VPWR VPWR _527_/HI _527_/LO sky130_fd_sc_hd__conb_1
XPHY_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_458_ VGND VGND VPWR VPWR _458_/HI _458_/LO sky130_fd_sc_hd__conb_1
XFILLER_70_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_517_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_389_ _382_/A VGND VGND VPWR VPWR _389_/X sky130_fd_sc_hd__buf_2
XFILLER_374_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_524_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_431_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[9\].yc blk.column\[11\].row\[9\].yc/cbitin blk.column\[11\].row\[9\].yc/cbitout
+ blk.column\[11\].row\[9\].yc/confclk blk.column\[11\].row\[9\].yc/confclko blk.column\[11\].row\[9\].yc/dempty
+ blk.column\[11\].row\[9\].yc/din[0] blk.column\[11\].row\[9\].yc/din[1] blk.column\[11\].row\[9\].yc/dout[0]
+ blk.column\[11\].row\[9\].yc/dout[1] blk.column\[11\].row\[9\].yc/hempty blk.column\[10\].row\[9\].yc/lempty
+ blk.column\[11\].row\[9\].yc/lempty blk.column\[11\].row\[9\].yc/lin[0] blk.column\[11\].row\[9\].yc/lin[1]
+ blk.column\[12\].row\[9\].yc/rin[0] blk.column\[12\].row\[9\].yc/rin[1] blk.column\[10\].row\[9\].yc/hempty
+ blk.column\[11\].row\[9\].yc/reset blk.column\[11\].row\[9\].yc/reseto blk.column\[11\].row\[9\].yc/rin[0]
+ blk.column\[11\].row\[9\].yc/rin[1] blk.column\[10\].row\[9\].yc/lin[0] blk.column\[10\].row\[9\].yc/lin[1]
+ blk.column\[11\].row\[9\].yc/uempty blk.column\[11\].row\[9\].yc/uin[0] blk.column\[11\].row\[9\].yc/uin[1]
+ blk.column\[11\].row\[8\].yc/din[0] blk.column\[11\].row\[8\].yc/din[1] blk.column\[11\].row\[8\].yc/dempty
+ blk.column\[11\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_58_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_399_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _312_/A VGND VGND VPWR VPWR _312_/Y sky130_fd_sc_hd__inv_2
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_295_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_291_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_533_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_488_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[13\].yc blk.column\[7\].row\[13\].yc/cbitin blk.column\[7\].row\[14\].yc/cbitin
+ blk.column\[7\].row\[13\].yc/confclk blk.column\[7\].row\[14\].yc/confclk blk.column\[7\].row\[13\].yc/dempty
+ blk.column\[7\].row\[13\].yc/din[0] blk.column\[7\].row\[13\].yc/din[1] blk.column\[7\].row\[14\].yc/uin[0]
+ blk.column\[7\].row\[14\].yc/uin[1] blk.column\[7\].row\[13\].yc/hempty blk.column\[6\].row\[13\].yc/lempty
+ blk.column\[7\].row\[13\].yc/lempty blk.column\[7\].row\[13\].yc/lin[0] blk.column\[7\].row\[13\].yc/lin[1]
+ blk.column\[8\].row\[13\].yc/rin[0] blk.column\[8\].row\[13\].yc/rin[1] blk.column\[6\].row\[13\].yc/hempty
+ blk.column\[7\].row\[13\].yc/reset blk.column\[7\].row\[14\].yc/reset blk.column\[7\].row\[13\].yc/rin[0]
+ blk.column\[7\].row\[13\].yc/rin[1] blk.column\[6\].row\[13\].yc/lin[0] blk.column\[6\].row\[13\].yc/lin[1]
+ blk.column\[7\].row\[13\].yc/uempty blk.column\[7\].row\[13\].yc/uin[0] blk.column\[7\].row\[13\].yc/uin[1]
+ blk.column\[7\].row\[12\].yc/din[0] blk.column\[7\].row\[12\].yc/din[1] blk.column\[7\].row\[12\].yc/dempty
+ blk.column\[7\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_152_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_473_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_541_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_394_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_359_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_307_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_502_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_498_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_269_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_539_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_499_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_270_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[4\].yc blk.column\[7\].row\[4\].yc/cbitin blk.column\[7\].row\[5\].yc/cbitin
+ blk.column\[7\].row\[4\].yc/confclk blk.column\[7\].row\[5\].yc/confclk blk.column\[7\].row\[4\].yc/dempty
+ blk.column\[7\].row\[4\].yc/din[0] blk.column\[7\].row\[4\].yc/din[1] blk.column\[7\].row\[5\].yc/uin[0]
+ blk.column\[7\].row\[5\].yc/uin[1] blk.column\[7\].row\[4\].yc/hempty blk.column\[6\].row\[4\].yc/lempty
+ blk.column\[7\].row\[4\].yc/lempty blk.column\[7\].row\[4\].yc/lin[0] blk.column\[7\].row\[4\].yc/lin[1]
+ blk.column\[8\].row\[4\].yc/rin[0] blk.column\[8\].row\[4\].yc/rin[1] blk.column\[6\].row\[4\].yc/hempty
+ blk.column\[7\].row\[4\].yc/reset blk.column\[7\].row\[5\].yc/reset blk.column\[7\].row\[4\].yc/rin[0]
+ blk.column\[7\].row\[4\].yc/rin[1] blk.column\[6\].row\[4\].yc/lin[0] blk.column\[6\].row\[4\].yc/lin[1]
+ blk.column\[7\].row\[4\].yc/uempty blk.column\[7\].row\[4\].yc/uin[0] blk.column\[7\].row\[4\].yc/uin[1]
+ blk.column\[7\].row\[3\].yc/din[0] blk.column\[7\].row\[3\].yc/din[1] blk.column\[7\].row\[3\].yc/dempty
+ blk.column\[7\].row\[5\].yc/uempty VPWR VGND ycell
XPHY_9357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_251_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_331_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_792_ wb_clk_i _336_/X VGND VGND VPWR VPWR _335_/A sky130_fd_sc_hd__dfxtp_4
XPHY_7977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_327_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_375_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_507_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_414_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_535_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_523_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_221_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_397_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_501_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_278_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_540_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_303_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[15\].yc blk.column\[14\].row\[15\].yc/cbitin la_data_out[46]
+ blk.column\[14\].row\[15\].yc/confclk blk.column\[14\].row\[15\].yc/confclko _449_/HI
+ _524_/LO _525_/LO blk.column\[14\].row\[15\].yc/dout[0] blk.column\[14\].row\[15\].yc/dout[1]
+ blk.column\[14\].row\[15\].yc/hempty blk.column\[13\].row\[15\].yc/lempty blk.column\[14\].row\[15\].yc/lempty
+ blk.column\[14\].row\[15\].yc/lin[0] blk.column\[14\].row\[15\].yc/lin[1] blk.column\[15\].row\[15\].yc/rin[0]
+ blk.column\[15\].row\[15\].yc/rin[1] blk.column\[13\].row\[15\].yc/hempty blk.column\[14\].row\[15\].yc/reset
+ blk.column\[14\].row\[15\].yc/reseto blk.column\[14\].row\[15\].yc/rin[0] blk.column\[14\].row\[15\].yc/rin[1]
+ blk.column\[13\].row\[15\].yc/lin[0] blk.column\[13\].row\[15\].yc/lin[1] blk.column\[14\].row\[15\].yc/uempty
+ blk.column\[14\].row\[15\].yc/uin[0] blk.column\[14\].row\[15\].yc/uin[1] blk.column\[14\].row\[14\].yc/din[0]
+ blk.column\[14\].row\[14\].yc/din[1] blk.column\[14\].row\[14\].yc/dempty blk.column\[14\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XPHY_5816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_385_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_396_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_421_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_530_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_2383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_470_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_775_ wb_clk_i _775_/D VGND VGND VPWR VPWR wbs_dat_o[31] sky130_fd_sc_hd__dfxtp_4
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_542_2059 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_539_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_297_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_317_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_367_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_317_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_308_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_276_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_508_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_418_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_480_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_560_ VGND VGND VPWR VPWR _560_/HI _560_/LO sky130_fd_sc_hd__conb_1
XPHY_4901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_491_ VGND VGND VPWR VPWR _491_/HI _491_/LO sky130_fd_sc_hd__conb_1
XPHY_4956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_537_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_231_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_758_ wb_clk_i _758_/D VGND VGND VPWR VPWR wbs_dat_o[14] sky130_fd_sc_hd__dfxtp_4
XFILLER_480_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_689_ VGND VGND VPWR VPWR _689_/HI la_data_out[73] sky130_fd_sc_hd__conb_1
XFILLER_34_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_396_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_241_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[6\].yc blk.column\[8\].row\[6\].yc/cbitin blk.column\[8\].row\[7\].yc/cbitin
+ blk.column\[8\].row\[6\].yc/confclk blk.column\[8\].row\[7\].yc/confclk blk.column\[8\].row\[6\].yc/dempty
+ blk.column\[8\].row\[6\].yc/din[0] blk.column\[8\].row\[6\].yc/din[1] blk.column\[8\].row\[7\].yc/uin[0]
+ blk.column\[8\].row\[7\].yc/uin[1] blk.column\[8\].row\[6\].yc/hempty blk.column\[7\].row\[6\].yc/lempty
+ blk.column\[8\].row\[6\].yc/lempty blk.column\[8\].row\[6\].yc/lin[0] blk.column\[8\].row\[6\].yc/lin[1]
+ blk.column\[9\].row\[6\].yc/rin[0] blk.column\[9\].row\[6\].yc/rin[1] blk.column\[7\].row\[6\].yc/hempty
+ blk.column\[8\].row\[6\].yc/reset blk.column\[8\].row\[7\].yc/reset blk.column\[8\].row\[6\].yc/rin[0]
+ blk.column\[8\].row\[6\].yc/rin[1] blk.column\[7\].row\[6\].yc/lin[0] blk.column\[7\].row\[6\].yc/lin[1]
+ blk.column\[8\].row\[6\].yc/uempty blk.column\[8\].row\[6\].yc/uin[0] blk.column\[8\].row\[6\].yc/uin[1]
+ blk.column\[8\].row\[5\].yc/din[0] blk.column\[8\].row\[5\].yc/din[1] blk.column\[8\].row\[5\].yc/dempty
+ blk.column\[8\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_519_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_500_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_493_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_288_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_612_ VGND VGND VPWR VPWR _612_/HI io_oeb[24] sky130_fd_sc_hd__conb_1
XPHY_6177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_543_ VGND VGND VPWR VPWR _543_/HI _543_/LO sky130_fd_sc_hd__conb_1
XFILLER_57_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_378_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_474_ VGND VGND VPWR VPWR _474_/HI _474_/LO sky130_fd_sc_hd__conb_1
XFILLER_504_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_536_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[14\].yc blk.column\[2\].row\[14\].yc/cbitin blk.column\[2\].row\[15\].yc/cbitin
+ blk.column\[2\].row\[14\].yc/confclk blk.column\[2\].row\[15\].yc/confclk blk.column\[2\].row\[14\].yc/dempty
+ blk.column\[2\].row\[14\].yc/din[0] blk.column\[2\].row\[14\].yc/din[1] blk.column\[2\].row\[15\].yc/uin[0]
+ blk.column\[2\].row\[15\].yc/uin[1] blk.column\[2\].row\[14\].yc/hempty blk.column\[1\].row\[14\].yc/lempty
+ blk.column\[2\].row\[14\].yc/lempty blk.column\[2\].row\[14\].yc/lin[0] blk.column\[2\].row\[14\].yc/lin[1]
+ blk.column\[3\].row\[14\].yc/rin[0] blk.column\[3\].row\[14\].yc/rin[1] blk.column\[1\].row\[14\].yc/hempty
+ blk.column\[2\].row\[14\].yc/reset blk.column\[2\].row\[15\].yc/reset blk.column\[2\].row\[14\].yc/rin[0]
+ blk.column\[2\].row\[14\].yc/rin[1] blk.column\[1\].row\[14\].yc/lin[0] blk.column\[1\].row\[14\].yc/lin[1]
+ blk.column\[2\].row\[14\].yc/uempty blk.column\[2\].row\[14\].yc/uin[0] blk.column\[2\].row\[14\].yc/uin[1]
+ blk.column\[2\].row\[13\].yc/din[0] blk.column\[2\].row\[13\].yc/din[1] blk.column\[2\].row\[13\].yc/dempty
+ blk.column\[2\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_298_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_515_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_353_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_352_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_246_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_261_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_525_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_440_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_475_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_516_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_526_ VGND VGND VPWR VPWR _526_/HI _526_/LO sky130_fd_sc_hd__conb_1
XPHY_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_457_ VGND VGND VPWR VPWR _457_/HI _457_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_376_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_388_ _384_/X wbs_dat_o[27] _779_/Q _382_/X VGND VGND VPWR VPWR _388_/X sky130_fd_sc_hd__o22a_4
XFILLER_509_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_505_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_424_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_2924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_491_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _309_/Y _310_/X wbs_dat_i[2] _310_/X VGND VGND VPWR VPWR _311_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_475_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_493_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_418_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_334_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_473_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_292_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_482_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_509_ VGND VGND VPWR VPWR _509_/HI _509_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_511_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_348_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_528_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_361_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_408_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[8\].yc blk.column\[9\].row\[8\].yc/cbitin blk.column\[9\].row\[9\].yc/cbitin
+ blk.column\[9\].row\[8\].yc/confclk blk.column\[9\].row\[9\].yc/confclk blk.column\[9\].row\[8\].yc/dempty
+ blk.column\[9\].row\[8\].yc/din[0] blk.column\[9\].row\[8\].yc/din[1] blk.column\[9\].row\[9\].yc/uin[0]
+ blk.column\[9\].row\[9\].yc/uin[1] blk.column\[9\].row\[8\].yc/hempty blk.column\[8\].row\[8\].yc/lempty
+ blk.column\[9\].row\[8\].yc/lempty blk.column\[9\].row\[8\].yc/lin[0] blk.column\[9\].row\[8\].yc/lin[1]
+ blk.column\[9\].row\[8\].yc/lout[0] blk.column\[9\].row\[8\].yc/lout[1] blk.column\[8\].row\[8\].yc/hempty
+ blk.column\[9\].row\[8\].yc/reset blk.column\[9\].row\[9\].yc/reset blk.column\[9\].row\[8\].yc/rin[0]
+ blk.column\[9\].row\[8\].yc/rin[1] blk.column\[8\].row\[8\].yc/lin[0] blk.column\[8\].row\[8\].yc/lin[1]
+ blk.column\[9\].row\[8\].yc/uempty blk.column\[9\].row\[8\].yc/uin[0] blk.column\[9\].row\[8\].yc/uin[1]
+ blk.column\[9\].row\[7\].yc/din[0] blk.column\[9\].row\[7\].yc/din[1] blk.column\[9\].row\[7\].yc/dempty
+ blk.column\[9\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_541_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_478_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_269_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_527_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_285_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_511_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_791_ wb_clk_i _791_/D VGND VGND VPWR VPWR _337_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_507_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_327_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_520_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_373_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_279_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_531_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_458_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_542_2753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_280_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_274_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_525_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_334_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_493_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_389_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_281_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_341_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_222_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_774_ wb_clk_i _385_/X VGND VGND VPWR VPWR wbs_dat_o[30] sky130_fd_sc_hd__dfxtp_4
XFILLER_542_2016 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[13\].row\[0\].yc la_data_in[109] blk.column\[13\].row\[1\].yc/cbitin
+ la_data_in[112] blk.column\[13\].row\[1\].yc/confclk blk.column\[13\].row\[0\].yc/dempty
+ blk.column\[13\].row\[0\].yc/din[0] blk.column\[13\].row\[0\].yc/din[1] blk.column\[13\].row\[1\].yc/uin[0]
+ blk.column\[13\].row\[1\].yc/uin[1] blk.column\[13\].row\[0\].yc/hempty blk.column\[12\].row\[0\].yc/lempty
+ blk.column\[13\].row\[0\].yc/lempty blk.column\[13\].row\[0\].yc/lin[0] blk.column\[13\].row\[0\].yc/lin[1]
+ blk.column\[14\].row\[0\].yc/rin[0] blk.column\[14\].row\[0\].yc/rin[1] blk.column\[12\].row\[0\].yc/hempty
+ la_data_in[113] blk.column\[13\].row\[1\].yc/reset blk.column\[13\].row\[0\].yc/rin[0]
+ blk.column\[13\].row\[0\].yc/rin[1] blk.column\[12\].row\[0\].yc/lin[0] blk.column\[12\].row\[0\].yc/lin[1]
+ _520_/LO la_data_in[90] la_data_in[91] la_data_out[26] la_data_out[27] blk.column\[13\].row\[0\].yc/vempty
+ blk.column\[13\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_181_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_542_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_451_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_391_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[1\].yc blk.column\[4\].row\[1\].yc/cbitin blk.column\[4\].row\[2\].yc/cbitin
+ blk.column\[4\].row\[1\].yc/confclk blk.column\[4\].row\[2\].yc/confclk blk.column\[4\].row\[1\].yc/dempty
+ blk.column\[4\].row\[1\].yc/din[0] blk.column\[4\].row\[1\].yc/din[1] blk.column\[4\].row\[2\].yc/uin[0]
+ blk.column\[4\].row\[2\].yc/uin[1] blk.column\[4\].row\[1\].yc/hempty blk.column\[3\].row\[1\].yc/lempty
+ blk.column\[4\].row\[1\].yc/lempty blk.column\[4\].row\[1\].yc/lin[0] blk.column\[4\].row\[1\].yc/lin[1]
+ blk.column\[5\].row\[1\].yc/rin[0] blk.column\[5\].row\[1\].yc/rin[1] blk.column\[3\].row\[1\].yc/hempty
+ blk.column\[4\].row\[1\].yc/reset blk.column\[4\].row\[2\].yc/reset blk.column\[4\].row\[1\].yc/rin[0]
+ blk.column\[4\].row\[1\].yc/rin[1] blk.column\[3\].row\[1\].yc/lin[0] blk.column\[3\].row\[1\].yc/lin[1]
+ blk.column\[4\].row\[1\].yc/uempty blk.column\[4\].row\[1\].yc/uin[0] blk.column\[4\].row\[1\].yc/uin[1]
+ blk.column\[4\].row\[0\].yc/din[0] blk.column\[4\].row\[0\].yc/din[1] blk.column\[4\].row\[0\].yc/dempty
+ blk.column\[4\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_209_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xblk.column\[11\].row\[11\].yc blk.column\[11\].row\[11\].yc/cbitin blk.column\[11\].row\[12\].yc/cbitin
+ blk.column\[11\].row\[11\].yc/confclk blk.column\[11\].row\[12\].yc/confclk blk.column\[11\].row\[11\].yc/dempty
+ blk.column\[11\].row\[11\].yc/din[0] blk.column\[11\].row\[11\].yc/din[1] blk.column\[11\].row\[12\].yc/uin[0]
+ blk.column\[11\].row\[12\].yc/uin[1] blk.column\[11\].row\[11\].yc/hempty blk.column\[10\].row\[11\].yc/lempty
+ blk.column\[11\].row\[11\].yc/lempty blk.column\[11\].row\[11\].yc/lin[0] blk.column\[11\].row\[11\].yc/lin[1]
+ blk.column\[12\].row\[11\].yc/rin[0] blk.column\[12\].row\[11\].yc/rin[1] blk.column\[10\].row\[11\].yc/hempty
+ blk.column\[11\].row\[11\].yc/reset blk.column\[11\].row\[12\].yc/reset blk.column\[11\].row\[11\].yc/rin[0]
+ blk.column\[11\].row\[11\].yc/rin[1] blk.column\[10\].row\[11\].yc/lin[0] blk.column\[10\].row\[11\].yc/lin[1]
+ blk.column\[11\].row\[11\].yc/uempty blk.column\[11\].row\[11\].yc/uin[0] blk.column\[11\].row\[11\].yc/uin[1]
+ blk.column\[11\].row\[10\].yc/din[0] blk.column\[11\].row\[10\].yc/din[1] blk.column\[11\].row\[10\].yc/dempty
+ blk.column\[11\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_522_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_512_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_529_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_499_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_509_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_536_2365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_317_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_514_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_517_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_489_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_490_ VGND VGND VPWR VPWR _490_/HI _490_/LO sky130_fd_sc_hd__conb_1
XPHY_4957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_276_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_2238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_342_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_526_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_235_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_757_ wb_clk_i _408_/X VGND VGND VPWR VPWR wbs_dat_o[13] sky130_fd_sc_hd__dfxtp_4
XFILLER_507_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_305_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_688_ VGND VGND VPWR VPWR _688_/HI la_data_out[72] sky130_fd_sc_hd__conb_1
XFILLER_21_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[12\].yc blk.column\[8\].row\[12\].yc/cbitin blk.column\[8\].row\[13\].yc/cbitin
+ blk.column\[8\].row\[12\].yc/confclk blk.column\[8\].row\[13\].yc/confclk blk.column\[8\].row\[12\].yc/dempty
+ blk.column\[8\].row\[12\].yc/din[0] blk.column\[8\].row\[12\].yc/din[1] blk.column\[8\].row\[13\].yc/uin[0]
+ blk.column\[8\].row\[13\].yc/uin[1] blk.column\[8\].row\[12\].yc/hempty blk.column\[7\].row\[12\].yc/lempty
+ blk.column\[8\].row\[12\].yc/lempty blk.column\[8\].row\[12\].yc/lin[0] blk.column\[8\].row\[12\].yc/lin[1]
+ blk.column\[9\].row\[12\].yc/rin[0] blk.column\[9\].row\[12\].yc/rin[1] blk.column\[7\].row\[12\].yc/hempty
+ blk.column\[8\].row\[12\].yc/reset blk.column\[8\].row\[13\].yc/reset blk.column\[8\].row\[12\].yc/rin[0]
+ blk.column\[8\].row\[12\].yc/rin[1] blk.column\[7\].row\[12\].yc/lin[0] blk.column\[7\].row\[12\].yc/lin[1]
+ blk.column\[8\].row\[12\].yc/uempty blk.column\[8\].row\[12\].yc/uin[0] blk.column\[8\].row\[12\].yc/uin[1]
+ blk.column\[8\].row\[11\].yc/din[0] blk.column\[8\].row\[11\].yc/din[1] blk.column\[8\].row\[11\].yc/dempty
+ blk.column\[8\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_236_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_509_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_532_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_410_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_287_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_611_ VGND VGND VPWR VPWR _611_/HI io_oeb[23] sky130_fd_sc_hd__conb_1
XPHY_6156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_291_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_328_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_542_ VGND VGND VPWR VPWR _542_/HI _542_/LO sky130_fd_sc_hd__conb_1
XPHY_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_473_ VGND VGND VPWR VPWR _473_/HI _473_/LO sky130_fd_sc_hd__conb_1
XFILLER_378_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_496_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_497_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_416_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[9\].yc blk.column\[0\].row\[9\].yc/cbitin blk.column\[0\].row\[9\].yc/cbitout
+ blk.column\[0\].row\[9\].yc/confclk blk.column\[0\].row\[9\].yc/confclko blk.column\[0\].row\[9\].yc/dempty
+ blk.column\[0\].row\[9\].yc/din[0] blk.column\[0\].row\[9\].yc/din[1] blk.column\[0\].row\[9\].yc/dout[0]
+ blk.column\[0\].row\[9\].yc/dout[1] blk.column\[0\].row\[9\].yc/hempty blk.column\[0\].row\[9\].yc/hempty2
+ blk.column\[0\].row\[9\].yc/lempty blk.column\[0\].row\[9\].yc/lin[0] blk.column\[0\].row\[9\].yc/lin[1]
+ blk.column\[1\].row\[9\].yc/rin[0] blk.column\[1\].row\[9\].yc/rin[1] _444_/HI blk.column\[0\].row\[9\].yc/reset
+ blk.column\[0\].row\[9\].yc/reseto _509_/LO _510_/LO blk.column\[0\].row\[9\].yc/rout[0]
+ blk.column\[0\].row\[9\].yc/rout[1] blk.column\[0\].row\[9\].yc/uempty blk.column\[0\].row\[9\].yc/uin[0]
+ blk.column\[0\].row\[9\].yc/uin[1] blk.column\[0\].row\[8\].yc/din[0] blk.column\[0\].row\[8\].yc/din[1]
+ blk.column\[0\].row\[8\].yc/dempty blk.column\[0\].row\[9\].yc/vempty2 VPWR VGND
+ ycell
XFILLER_526_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_522_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_318_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_352_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_494_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_527_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_525_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_438_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_418_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_517_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_513_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[2\].yc blk.column\[14\].row\[2\].yc/cbitin blk.column\[14\].row\[3\].yc/cbitin
+ blk.column\[14\].row\[2\].yc/confclk blk.column\[14\].row\[3\].yc/confclk blk.column\[14\].row\[2\].yc/dempty
+ blk.column\[14\].row\[2\].yc/din[0] blk.column\[14\].row\[2\].yc/din[1] blk.column\[14\].row\[3\].yc/uin[0]
+ blk.column\[14\].row\[3\].yc/uin[1] blk.column\[14\].row\[2\].yc/hempty blk.column\[13\].row\[2\].yc/lempty
+ blk.column\[14\].row\[2\].yc/lempty blk.column\[14\].row\[2\].yc/lin[0] blk.column\[14\].row\[2\].yc/lin[1]
+ blk.column\[15\].row\[2\].yc/rin[0] blk.column\[15\].row\[2\].yc/rin[1] blk.column\[13\].row\[2\].yc/hempty
+ blk.column\[14\].row\[2\].yc/reset blk.column\[14\].row\[3\].yc/reset blk.column\[14\].row\[2\].yc/rin[0]
+ blk.column\[14\].row\[2\].yc/rin[1] blk.column\[13\].row\[2\].yc/lin[0] blk.column\[13\].row\[2\].yc/lin[1]
+ blk.column\[14\].row\[2\].yc/uempty blk.column\[14\].row\[2\].yc/uin[0] blk.column\[14\].row\[2\].yc/uin[1]
+ blk.column\[14\].row\[1\].yc/din[0] blk.column\[14\].row\[1\].yc/din[1] blk.column\[14\].row\[1\].yc/dempty
+ blk.column\[14\].row\[3\].yc/uempty VPWR VGND ycell
XPHY_11324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_296_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_2967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_10645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[14\].yc blk.column\[15\].row\[14\].yc/cbitin blk.column\[15\].row\[15\].yc/cbitin
+ blk.column\[15\].row\[14\].yc/confclk blk.column\[15\].row\[15\].yc/confclk blk.column\[15\].row\[14\].yc/dempty
+ blk.column\[15\].row\[14\].yc/din[0] blk.column\[15\].row\[14\].yc/din[1] blk.column\[15\].row\[15\].yc/uin[0]
+ blk.column\[15\].row\[15\].yc/uin[1] blk.column\[15\].row\[14\].yc/hempty blk.column\[14\].row\[14\].yc/lempty
+ _455_/HI _537_/LO _538_/LO blk.column\[15\].row\[14\].yc/lout[0] blk.column\[15\].row\[14\].yc/lout[1]
+ blk.column\[14\].row\[14\].yc/hempty blk.column\[15\].row\[14\].yc/reset blk.column\[15\].row\[15\].yc/reset
+ blk.column\[15\].row\[14\].yc/rin[0] blk.column\[15\].row\[14\].yc/rin[1] blk.column\[14\].row\[14\].yc/lin[0]
+ blk.column\[14\].row\[14\].yc/lin[1] blk.column\[15\].row\[14\].yc/uempty blk.column\[15\].row\[14\].yc/uin[0]
+ blk.column\[15\].row\[14\].yc/uin[1] blk.column\[15\].row\[13\].yc/din[0] blk.column\[15\].row\[13\].yc/din[1]
+ blk.column\[15\].row\[13\].yc/dempty blk.column\[15\].row\[15\].yc/uempty VPWR VGND
+ ycell
XPHY_10667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_421_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_525_ VGND VGND VPWR VPWR _525_/HI _525_/LO sky130_fd_sc_hd__conb_1
XPHY_5296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[3\].yc blk.column\[5\].row\[3\].yc/cbitin blk.column\[5\].row\[4\].yc/cbitin
+ blk.column\[5\].row\[3\].yc/confclk blk.column\[5\].row\[4\].yc/confclk blk.column\[5\].row\[3\].yc/dempty
+ blk.column\[5\].row\[3\].yc/din[0] blk.column\[5\].row\[3\].yc/din[1] blk.column\[5\].row\[4\].yc/uin[0]
+ blk.column\[5\].row\[4\].yc/uin[1] blk.column\[5\].row\[3\].yc/hempty blk.column\[4\].row\[3\].yc/lempty
+ blk.column\[5\].row\[3\].yc/lempty blk.column\[5\].row\[3\].yc/lin[0] blk.column\[5\].row\[3\].yc/lin[1]
+ blk.column\[6\].row\[3\].yc/rin[0] blk.column\[6\].row\[3\].yc/rin[1] blk.column\[4\].row\[3\].yc/hempty
+ blk.column\[5\].row\[3\].yc/reset blk.column\[5\].row\[4\].yc/reset blk.column\[5\].row\[3\].yc/rin[0]
+ blk.column\[5\].row\[3\].yc/rin[1] blk.column\[4\].row\[3\].yc/lin[0] blk.column\[4\].row\[3\].yc/lin[1]
+ blk.column\[5\].row\[3\].yc/uempty blk.column\[5\].row\[3\].yc/uin[0] blk.column\[5\].row\[3\].yc/uin[1]
+ blk.column\[5\].row\[2\].yc/din[0] blk.column\[5\].row\[2\].yc/din[1] blk.column\[5\].row\[2\].yc/dempty
+ blk.column\[5\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_205_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_456_ VGND VGND VPWR VPWR _456_/HI _456_/LO sky130_fd_sc_hd__conb_1
XFILLER_321_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_376_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_387_ _384_/X wbs_dat_o[28] _780_/Q _382_/X VGND VGND VPWR VPWR _772_/D sky130_fd_sc_hd__o22a_4
XFILLER_517_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_334_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_313_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_463_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_500_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_539_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_468_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_2936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_288_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_299_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_405_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_310_ _298_/A VGND VGND VPWR VPWR _310_/X sky130_fd_sc_hd__buf_2
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_449_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_295_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_316_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_533_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_408_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_523_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_508_ VGND VGND VPWR VPWR _508_/HI _508_/LO sky130_fd_sc_hd__conb_1
XPHY_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_394_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_439_ VGND VGND VPWR VPWR _439_/HI _439_/LO sky130_fd_sc_hd__conb_1
XFILLER_536_2706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_347_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_520_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_348_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_541_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_251_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_498_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1018 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_359_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_472_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_790_ wb_clk_i _790_/D VGND VGND VPWR VPWR _790_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_491_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_215_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_430_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_431_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_286_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_380_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[13\].yc blk.column\[3\].row\[13\].yc/cbitin blk.column\[3\].row\[14\].yc/cbitin
+ blk.column\[3\].row\[13\].yc/confclk blk.column\[3\].row\[14\].yc/confclk blk.column\[3\].row\[13\].yc/dempty
+ blk.column\[3\].row\[13\].yc/din[0] blk.column\[3\].row\[13\].yc/din[1] blk.column\[3\].row\[14\].yc/uin[0]
+ blk.column\[3\].row\[14\].yc/uin[1] blk.column\[3\].row\[13\].yc/hempty blk.column\[2\].row\[13\].yc/lempty
+ blk.column\[3\].row\[13\].yc/lempty blk.column\[3\].row\[13\].yc/lin[0] blk.column\[3\].row\[13\].yc/lin[1]
+ blk.column\[4\].row\[13\].yc/rin[0] blk.column\[4\].row\[13\].yc/rin[1] blk.column\[2\].row\[13\].yc/hempty
+ blk.column\[3\].row\[13\].yc/reset blk.column\[3\].row\[14\].yc/reset blk.column\[3\].row\[13\].yc/rin[0]
+ blk.column\[3\].row\[13\].yc/rin[1] blk.column\[2\].row\[13\].yc/lin[0] blk.column\[2\].row\[13\].yc/lin[1]
+ blk.column\[3\].row\[13\].yc/uempty blk.column\[3\].row\[13\].yc/uin[0] blk.column\[3\].row\[13\].yc/uin[1]
+ blk.column\[3\].row\[12\].yc/din[0] blk.column\[3\].row\[12\].yc/din[1] blk.column\[3\].row\[12\].yc/dempty
+ blk.column\[3\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_536_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_517_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_528_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_256_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[15\].row\[4\].yc blk.column\[15\].row\[4\].yc/cbitin blk.column\[15\].row\[5\].yc/cbitin
+ blk.column\[15\].row\[4\].yc/confclk blk.column\[15\].row\[5\].yc/confclk blk.column\[15\].row\[4\].yc/dempty
+ blk.column\[15\].row\[4\].yc/din[0] blk.column\[15\].row\[4\].yc/din[1] blk.column\[15\].row\[5\].yc/uin[0]
+ blk.column\[15\].row\[5\].yc/uin[1] blk.column\[15\].row\[4\].yc/hempty blk.column\[14\].row\[4\].yc/lempty
+ _461_/HI _549_/LO _550_/LO blk.column\[15\].row\[4\].yc/lout[0] blk.column\[15\].row\[4\].yc/lout[1]
+ blk.column\[14\].row\[4\].yc/hempty blk.column\[15\].row\[4\].yc/reset blk.column\[15\].row\[5\].yc/reset
+ blk.column\[15\].row\[4\].yc/rin[0] blk.column\[15\].row\[4\].yc/rin[1] blk.column\[14\].row\[4\].yc/lin[0]
+ blk.column\[14\].row\[4\].yc/lin[1] blk.column\[15\].row\[4\].yc/uempty blk.column\[15\].row\[4\].yc/uin[0]
+ blk.column\[15\].row\[4\].yc/uin[1] blk.column\[15\].row\[3\].yc/din[0] blk.column\[15\].row\[3\].yc/din[1]
+ blk.column\[15\].row\[3\].yc/dempty blk.column\[15\].row\[5\].yc/uempty VPWR VGND
+ ycell
XFILLER_159_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_368_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_380_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[5\].yc blk.column\[6\].row\[5\].yc/cbitin blk.column\[6\].row\[6\].yc/cbitin
+ blk.column\[6\].row\[5\].yc/confclk blk.column\[6\].row\[6\].yc/confclk blk.column\[6\].row\[5\].yc/dempty
+ blk.column\[6\].row\[5\].yc/din[0] blk.column\[6\].row\[5\].yc/din[1] blk.column\[6\].row\[6\].yc/uin[0]
+ blk.column\[6\].row\[6\].yc/uin[1] blk.column\[6\].row\[5\].yc/hempty blk.column\[5\].row\[5\].yc/lempty
+ blk.column\[6\].row\[5\].yc/lempty blk.column\[6\].row\[5\].yc/lin[0] blk.column\[6\].row\[5\].yc/lin[1]
+ blk.column\[7\].row\[5\].yc/rin[0] blk.column\[7\].row\[5\].yc/rin[1] blk.column\[5\].row\[5\].yc/hempty
+ blk.column\[6\].row\[5\].yc/reset blk.column\[6\].row\[6\].yc/reset blk.column\[6\].row\[5\].yc/rin[0]
+ blk.column\[6\].row\[5\].yc/rin[1] blk.column\[5\].row\[5\].yc/lin[0] blk.column\[5\].row\[5\].yc/lin[1]
+ blk.column\[6\].row\[5\].yc/uempty blk.column\[6\].row\[5\].yc/uin[0] blk.column\[6\].row\[5\].yc/uin[1]
+ blk.column\[6\].row\[4\].yc/din[0] blk.column\[6\].row\[4\].yc/din[1] blk.column\[6\].row\[4\].yc/dempty
+ blk.column\[6\].row\[6\].yc/uempty VPWR VGND ycell
XPHY_8499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_773_ wb_clk_i _386_/X VGND VGND VPWR VPWR wbs_dat_o[29] sky130_fd_sc_hd__dfxtp_4
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_262_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_420_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_531_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_518_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_391_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_317_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_529_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_442_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_514_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_331_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_510_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_445_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_404_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_301_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_521_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_495_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[15\].yc blk.column\[10\].row\[15\].yc/cbitin la_data_out[42]
+ blk.column\[10\].row\[15\].yc/confclk blk.column\[10\].row\[15\].yc/confclko _445_/HI
+ _512_/LO _513_/LO blk.column\[10\].row\[15\].yc/dout[0] blk.column\[10\].row\[15\].yc/dout[1]
+ blk.column\[10\].row\[15\].yc/hempty blk.column\[9\].row\[15\].yc/lempty blk.column\[10\].row\[15\].yc/lempty
+ blk.column\[10\].row\[15\].yc/lin[0] blk.column\[10\].row\[15\].yc/lin[1] blk.column\[11\].row\[15\].yc/rin[0]
+ blk.column\[11\].row\[15\].yc/rin[1] blk.column\[9\].row\[15\].yc/hempty blk.column\[10\].row\[15\].yc/reset
+ blk.column\[10\].row\[15\].yc/reseto blk.column\[9\].row\[15\].yc/lout[0] blk.column\[9\].row\[15\].yc/lout[1]
+ blk.column\[9\].row\[15\].yc/lin[0] blk.column\[9\].row\[15\].yc/lin[1] blk.column\[10\].row\[15\].yc/uempty
+ blk.column\[10\].row\[15\].yc/uin[0] blk.column\[10\].row\[15\].yc/uin[1] blk.column\[10\].row\[14\].yc/din[0]
+ blk.column\[10\].row\[14\].yc/din[1] blk.column\[10\].row\[14\].yc/dempty blk.column\[10\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_314_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_532_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_342_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_756_ wb_clk_i _756_/D VGND VGND VPWR VPWR wbs_dat_o[12] sky130_fd_sc_hd__dfxtp_4
XPHY_6872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_687_ VGND VGND VPWR VPWR _687_/HI la_data_out[71] sky130_fd_sc_hd__conb_1
XFILLER_160_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_379_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_455_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_220_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_271_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_313_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_397_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_529_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_610_ VGND VGND VPWR VPWR _610_/HI io_oeb[22] sky130_fd_sc_hd__conb_1
XPHY_6146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_291_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_541_ VGND VGND VPWR VPWR _541_/HI _541_/LO sky130_fd_sc_hd__conb_1
XPHY_5456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_472_ VGND VGND VPWR VPWR _472_/HI _472_/LO sky130_fd_sc_hd__conb_1
XFILLER_433_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2090 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_343_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_519_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_270_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_255_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_808_ wb_clk_i _808_/D VGND VGND VPWR VPWR wbs_ack_o sky130_fd_sc_hd__dfxtp_4
XFILLER_166_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_307_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_739_ VGND VGND VPWR VPWR _739_/HI la_data_out[123] sky130_fd_sc_hd__conb_1
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_507_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_537_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_514_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_511_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_273_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_505_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_227_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_415_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_307_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_368_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_383_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_254_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[7\].yc blk.column\[7\].row\[7\].yc/cbitin blk.column\[7\].row\[8\].yc/cbitin
+ blk.column\[7\].row\[7\].yc/confclk blk.column\[7\].row\[8\].yc/confclk blk.column\[7\].row\[7\].yc/dempty
+ blk.column\[7\].row\[7\].yc/din[0] blk.column\[7\].row\[7\].yc/din[1] blk.column\[7\].row\[8\].yc/uin[0]
+ blk.column\[7\].row\[8\].yc/uin[1] blk.column\[7\].row\[7\].yc/hempty blk.column\[6\].row\[7\].yc/lempty
+ blk.column\[7\].row\[7\].yc/lempty blk.column\[7\].row\[7\].yc/lin[0] blk.column\[7\].row\[7\].yc/lin[1]
+ blk.column\[8\].row\[7\].yc/rin[0] blk.column\[8\].row\[7\].yc/rin[1] blk.column\[6\].row\[7\].yc/hempty
+ blk.column\[7\].row\[7\].yc/reset blk.column\[7\].row\[8\].yc/reset blk.column\[7\].row\[7\].yc/rin[0]
+ blk.column\[7\].row\[7\].yc/rin[1] blk.column\[6\].row\[7\].yc/lin[0] blk.column\[6\].row\[7\].yc/lin[1]
+ blk.column\[7\].row\[7\].yc/uempty blk.column\[7\].row\[7\].yc/uin[0] blk.column\[7\].row\[7\].yc/uin[1]
+ blk.column\[7\].row\[6\].yc/din[0] blk.column\[7\].row\[6\].yc/din[1] blk.column\[7\].row\[6\].yc/dempty
+ blk.column\[7\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_307_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_351_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_314_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_524_ VGND VGND VPWR VPWR _524_/HI _524_/LO sky130_fd_sc_hd__conb_1
XPHY_5286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ VGND VGND VPWR VPWR _455_/HI _455_/LO sky130_fd_sc_hd__conb_1
XFILLER_35_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_386_ _384_/X wbs_dat_o[29] _365_/A _382_/X VGND VGND VPWR VPWR _386_/X sky130_fd_sc_hd__o22a_4
XFILLER_185_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_491_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_348_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_495_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_506_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_270_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_522_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[10\].yc blk.column\[12\].row\[9\].yc/cbitout blk.column\[12\].row\[11\].yc/cbitin
+ blk.column\[12\].row\[9\].yc/confclko blk.column\[12\].row\[11\].yc/confclk blk.column\[12\].row\[10\].yc/dempty
+ blk.column\[12\].row\[10\].yc/din[0] blk.column\[12\].row\[10\].yc/din[1] blk.column\[12\].row\[11\].yc/uin[0]
+ blk.column\[12\].row\[11\].yc/uin[1] blk.column\[12\].row\[10\].yc/hempty blk.column\[11\].row\[10\].yc/lempty
+ blk.column\[12\].row\[10\].yc/lempty blk.column\[12\].row\[10\].yc/lin[0] blk.column\[12\].row\[10\].yc/lin[1]
+ blk.column\[13\].row\[10\].yc/rin[0] blk.column\[13\].row\[10\].yc/rin[1] blk.column\[11\].row\[10\].yc/hempty
+ blk.column\[12\].row\[9\].yc/reseto blk.column\[12\].row\[11\].yc/reset blk.column\[12\].row\[10\].yc/rin[0]
+ blk.column\[12\].row\[10\].yc/rin[1] blk.column\[11\].row\[10\].yc/lin[0] blk.column\[11\].row\[10\].yc/lin[1]
+ blk.column\[12\].row\[9\].yc/vempty2 blk.column\[12\].row\[9\].yc/dout[0] blk.column\[12\].row\[9\].yc/dout[1]
+ blk.column\[12\].row\[9\].yc/din[0] blk.column\[12\].row\[9\].yc/din[1] blk.column\[12\].row\[9\].yc/dempty
+ blk.column\[12\].row\[11\].yc/uempty VPWR VGND ycell
XFILLER_533_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_504_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_299_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_318_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_512_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_10454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_252_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_507_ VGND VGND VPWR VPWR _507_/HI _507_/LO sky130_fd_sc_hd__conb_1
XPHY_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_438_ VGND VGND VPWR VPWR _438_/HI _438_/LO sky130_fd_sc_hd__conb_1
XFILLER_394_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_369_ _368_/Y _366_/X wbs_dat_i[28] _366_/X VGND VGND VPWR VPWR _369_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_11_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_228_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xblk.column\[2\].row\[0\].yc la_data_in[98] blk.column\[2\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[2\].row\[1\].yc/confclk blk.column\[2\].row\[0\].yc/dempty blk.column\[2\].row\[0\].yc/din[0]
+ blk.column\[2\].row\[0\].yc/din[1] blk.column\[2\].row\[1\].yc/uin[0] blk.column\[2\].row\[1\].yc/uin[1]
+ blk.column\[2\].row\[0\].yc/hempty blk.column\[1\].row\[0\].yc/lempty blk.column\[2\].row\[0\].yc/lempty
+ blk.column\[2\].row\[0\].yc/lin[0] blk.column\[2\].row\[0\].yc/lin[1] blk.column\[3\].row\[0\].yc/rin[0]
+ blk.column\[3\].row\[0\].yc/rin[1] blk.column\[1\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[2\].row\[1\].yc/reset blk.column\[2\].row\[0\].yc/rin[0] blk.column\[2\].row\[0\].yc/rin[1]
+ blk.column\[1\].row\[0\].yc/lin[0] blk.column\[1\].row\[0\].yc/lin[1] _564_/LO la_data_in[68]
+ la_data_in[69] la_data_out[4] la_data_out[5] blk.column\[2\].row\[0\].yc/vempty
+ blk.column\[2\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_408_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_397_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_224_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_355_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[11\].yc blk.column\[9\].row\[11\].yc/cbitin blk.column\[9\].row\[12\].yc/cbitin
+ blk.column\[9\].row\[11\].yc/confclk blk.column\[9\].row\[12\].yc/confclk blk.column\[9\].row\[11\].yc/dempty
+ blk.column\[9\].row\[11\].yc/din[0] blk.column\[9\].row\[11\].yc/din[1] blk.column\[9\].row\[12\].yc/uin[0]
+ blk.column\[9\].row\[12\].yc/uin[1] blk.column\[9\].row\[11\].yc/hempty blk.column\[8\].row\[11\].yc/lempty
+ blk.column\[9\].row\[11\].yc/lempty blk.column\[9\].row\[11\].yc/lin[0] blk.column\[9\].row\[11\].yc/lin[1]
+ blk.column\[9\].row\[11\].yc/lout[0] blk.column\[9\].row\[11\].yc/lout[1] blk.column\[8\].row\[11\].yc/hempty
+ blk.column\[9\].row\[11\].yc/reset blk.column\[9\].row\[12\].yc/reset blk.column\[9\].row\[11\].yc/rin[0]
+ blk.column\[9\].row\[11\].yc/rin[1] blk.column\[8\].row\[11\].yc/lin[0] blk.column\[8\].row\[11\].yc/lin[1]
+ blk.column\[9\].row\[11\].yc/uempty blk.column\[9\].row\[11\].yc/uin[0] blk.column\[9\].row\[11\].yc/uin[1]
+ blk.column\[9\].row\[10\].yc/din[0] blk.column\[9\].row\[10\].yc/din[1] blk.column\[9\].row\[10\].yc/dempty
+ blk.column\[9\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_14_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_535_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_216_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_415_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_320_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_376_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_423_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_373_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_488_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_488_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_414_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_379_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_540_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_458_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_533_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_315_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_437_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[9\].yc blk.column\[8\].row\[9\].yc/cbitin blk.column\[8\].row\[9\].yc/cbitout
+ blk.column\[8\].row\[9\].yc/confclk blk.column\[8\].row\[9\].yc/confclko blk.column\[8\].row\[9\].yc/dempty
+ blk.column\[8\].row\[9\].yc/din[0] blk.column\[8\].row\[9\].yc/din[1] blk.column\[8\].row\[9\].yc/dout[0]
+ blk.column\[8\].row\[9\].yc/dout[1] blk.column\[8\].row\[9\].yc/hempty blk.column\[7\].row\[9\].yc/lempty
+ blk.column\[8\].row\[9\].yc/lempty blk.column\[8\].row\[9\].yc/lin[0] blk.column\[8\].row\[9\].yc/lin[1]
+ blk.column\[9\].row\[9\].yc/rin[0] blk.column\[9\].row\[9\].yc/rin[1] blk.column\[7\].row\[9\].yc/hempty
+ blk.column\[8\].row\[9\].yc/reset blk.column\[8\].row\[9\].yc/reseto blk.column\[8\].row\[9\].yc/rin[0]
+ blk.column\[8\].row\[9\].yc/rin[1] blk.column\[7\].row\[9\].yc/lin[0] blk.column\[7\].row\[9\].yc/lin[1]
+ blk.column\[8\].row\[9\].yc/uempty blk.column\[8\].row\[9\].yc/uin[0] blk.column\[8\].row\[9\].yc/uin[1]
+ blk.column\[8\].row\[8\].yc/din[0] blk.column\[8\].row\[8\].yc/din[1] blk.column\[8\].row\[8\].yc/dempty
+ blk.column\[8\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_220_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_535_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_368_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_772_ wb_clk_i _772_/D VGND VGND VPWR VPWR wbs_dat_o[28] sky130_fd_sc_hd__dfxtp_4
XFILLER_492_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_501_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_487_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_455_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_384_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_506_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_269_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_446_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_345_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_444_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_499_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_308_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_477_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_282_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_331_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_512_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_404_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_220_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_490_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_755_ wb_clk_i _411_/X VGND VGND VPWR VPWR wbs_dat_o[11] sky130_fd_sc_hd__dfxtp_4
XFILLER_526_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_507_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_686_ VGND VGND VPWR VPWR _686_/HI la_data_out[70] sky130_fd_sc_hd__conb_1
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[1\].yc blk.column\[12\].row\[1\].yc/cbitin blk.column\[12\].row\[2\].yc/cbitin
+ blk.column\[12\].row\[1\].yc/confclk blk.column\[12\].row\[2\].yc/confclk blk.column\[12\].row\[1\].yc/dempty
+ blk.column\[12\].row\[1\].yc/din[0] blk.column\[12\].row\[1\].yc/din[1] blk.column\[12\].row\[2\].yc/uin[0]
+ blk.column\[12\].row\[2\].yc/uin[1] blk.column\[12\].row\[1\].yc/hempty blk.column\[11\].row\[1\].yc/lempty
+ blk.column\[12\].row\[1\].yc/lempty blk.column\[12\].row\[1\].yc/lin[0] blk.column\[12\].row\[1\].yc/lin[1]
+ blk.column\[13\].row\[1\].yc/rin[0] blk.column\[13\].row\[1\].yc/rin[1] blk.column\[11\].row\[1\].yc/hempty
+ blk.column\[12\].row\[1\].yc/reset blk.column\[12\].row\[2\].yc/reset blk.column\[12\].row\[1\].yc/rin[0]
+ blk.column\[12\].row\[1\].yc/rin[1] blk.column\[11\].row\[1\].yc/lin[0] blk.column\[11\].row\[1\].yc/lin[1]
+ blk.column\[12\].row\[1\].yc/uempty blk.column\[12\].row\[1\].yc/uin[0] blk.column\[12\].row\[1\].yc/uin[1]
+ blk.column\[12\].row\[0\].yc/din[0] blk.column\[12\].row\[0\].yc/din[1] blk.column\[12\].row\[0\].yc/dempty
+ blk.column\[12\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_188_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_507_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_455_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[2\].yc blk.column\[3\].row\[2\].yc/cbitin blk.column\[3\].row\[3\].yc/cbitin
+ blk.column\[3\].row\[2\].yc/confclk blk.column\[3\].row\[3\].yc/confclk blk.column\[3\].row\[2\].yc/dempty
+ blk.column\[3\].row\[2\].yc/din[0] blk.column\[3\].row\[2\].yc/din[1] blk.column\[3\].row\[3\].yc/uin[0]
+ blk.column\[3\].row\[3\].yc/uin[1] blk.column\[3\].row\[2\].yc/hempty blk.column\[2\].row\[2\].yc/lempty
+ blk.column\[3\].row\[2\].yc/lempty blk.column\[3\].row\[2\].yc/lin[0] blk.column\[3\].row\[2\].yc/lin[1]
+ blk.column\[4\].row\[2\].yc/rin[0] blk.column\[4\].row\[2\].yc/rin[1] blk.column\[2\].row\[2\].yc/hempty
+ blk.column\[3\].row\[2\].yc/reset blk.column\[3\].row\[3\].yc/reset blk.column\[3\].row\[2\].yc/rin[0]
+ blk.column\[3\].row\[2\].yc/rin[1] blk.column\[2\].row\[2\].yc/lin[0] blk.column\[2\].row\[2\].yc/lin[1]
+ blk.column\[3\].row\[2\].yc/uempty blk.column\[3\].row\[2\].yc/uin[0] blk.column\[3\].row\[2\].yc/uin[1]
+ blk.column\[3\].row\[1\].yc/din[0] blk.column\[3\].row\[1\].yc/din[1] blk.column\[3\].row\[1\].yc/dempty
+ blk.column\[3\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_316_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_522_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_323_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_499_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_358_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_520_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_520_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_276_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_493_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_406_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_291_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_540_ VGND VGND VPWR VPWR _540_/HI _540_/LO sky130_fd_sc_hd__conb_1
XPHY_5457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_478_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_471_ VGND VGND VPWR VPWR _471_/HI _471_/LO sky130_fd_sc_hd__conb_1
XFILLER_263_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_439_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_489_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_485_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_266_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_807_ wb_clk_i _299_/X VGND VGND VPWR VPWR _807_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_7382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_307_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_738_ VGND VGND VPWR VPWR _738_/HI la_data_out[122] sky130_fd_sc_hd__conb_1
XFILLER_526_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_669_ VGND VGND VPWR VPWR _669_/HI la_data_out[53] sky130_fd_sc_hd__conb_1
XFILLER_507_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_528_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_259_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_258_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_540_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[12\].yc blk.column\[4\].row\[12\].yc/cbitin blk.column\[4\].row\[13\].yc/cbitin
+ blk.column\[4\].row\[12\].yc/confclk blk.column\[4\].row\[13\].yc/confclk blk.column\[4\].row\[12\].yc/dempty
+ blk.column\[4\].row\[12\].yc/din[0] blk.column\[4\].row\[12\].yc/din[1] blk.column\[4\].row\[13\].yc/uin[0]
+ blk.column\[4\].row\[13\].yc/uin[1] blk.column\[4\].row\[12\].yc/hempty blk.column\[3\].row\[12\].yc/lempty
+ blk.column\[4\].row\[12\].yc/lempty blk.column\[4\].row\[12\].yc/lin[0] blk.column\[4\].row\[12\].yc/lin[1]
+ blk.column\[5\].row\[12\].yc/rin[0] blk.column\[5\].row\[12\].yc/rin[1] blk.column\[3\].row\[12\].yc/hempty
+ blk.column\[4\].row\[12\].yc/reset blk.column\[4\].row\[13\].yc/reset blk.column\[4\].row\[12\].yc/rin[0]
+ blk.column\[4\].row\[12\].yc/rin[1] blk.column\[3\].row\[12\].yc/lin[0] blk.column\[3\].row\[12\].yc/lin[1]
+ blk.column\[4\].row\[12\].yc/uempty blk.column\[4\].row\[12\].yc/uin[0] blk.column\[4\].row\[12\].yc/uin[1]
+ blk.column\[4\].row\[11\].yc/din[0] blk.column\[4\].row\[11\].yc/din[1] blk.column\[4\].row\[11\].yc/dempty
+ blk.column\[4\].row\[13\].yc/uempty VPWR VGND ycell
XFILLER_260_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_368_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_314_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_351_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_464_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_261_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_453_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_523_ VGND VGND VPWR VPWR _523_/HI _523_/LO sky130_fd_sc_hd__conb_1
XPHY_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_454_ VGND VGND VPWR VPWR _454_/HI _454_/LO sky130_fd_sc_hd__conb_1
XFILLER_360_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_385_ _384_/X wbs_dat_o[30] _363_/A _382_/X VGND VGND VPWR VPWR _385_/X sky130_fd_sc_hd__o22a_4
XFILLER_14_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_534_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_320_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_306_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_520_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_221_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_505_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_535_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_531_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_412_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[13\].row\[3\].yc blk.column\[13\].row\[3\].yc/cbitin blk.column\[13\].row\[4\].yc/cbitin
+ blk.column\[13\].row\[3\].yc/confclk blk.column\[13\].row\[4\].yc/confclk blk.column\[13\].row\[3\].yc/dempty
+ blk.column\[13\].row\[3\].yc/din[0] blk.column\[13\].row\[3\].yc/din[1] blk.column\[13\].row\[4\].yc/uin[0]
+ blk.column\[13\].row\[4\].yc/uin[1] blk.column\[13\].row\[3\].yc/hempty blk.column\[12\].row\[3\].yc/lempty
+ blk.column\[13\].row\[3\].yc/lempty blk.column\[13\].row\[3\].yc/lin[0] blk.column\[13\].row\[3\].yc/lin[1]
+ blk.column\[14\].row\[3\].yc/rin[0] blk.column\[14\].row\[3\].yc/rin[1] blk.column\[12\].row\[3\].yc/hempty
+ blk.column\[13\].row\[3\].yc/reset blk.column\[13\].row\[4\].yc/reset blk.column\[13\].row\[3\].yc/rin[0]
+ blk.column\[13\].row\[3\].yc/rin[1] blk.column\[12\].row\[3\].yc/lin[0] blk.column\[12\].row\[3\].yc/lin[1]
+ blk.column\[13\].row\[3\].yc/uempty blk.column\[13\].row\[3\].yc/uin[0] blk.column\[13\].row\[3\].yc/uin[1]
+ blk.column\[13\].row\[2\].yc/din[0] blk.column\[13\].row\[2\].yc/din[1] blk.column\[13\].row\[2\].yc/dempty
+ blk.column\[13\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_426_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_304_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_430_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_506_ VGND VGND VPWR VPWR _506_/HI _506_/LO sky130_fd_sc_hd__conb_1
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_437_ VGND VGND VPWR VPWR _437_/HI _437_/LO sky130_fd_sc_hd__conb_1
XFILLER_399_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xblk.column\[4\].row\[4\].yc blk.column\[4\].row\[4\].yc/cbitin blk.column\[4\].row\[5\].yc/cbitin
+ blk.column\[4\].row\[4\].yc/confclk blk.column\[4\].row\[5\].yc/confclk blk.column\[4\].row\[4\].yc/dempty
+ blk.column\[4\].row\[4\].yc/din[0] blk.column\[4\].row\[4\].yc/din[1] blk.column\[4\].row\[5\].yc/uin[0]
+ blk.column\[4\].row\[5\].yc/uin[1] blk.column\[4\].row\[4\].yc/hempty blk.column\[3\].row\[4\].yc/lempty
+ blk.column\[4\].row\[4\].yc/lempty blk.column\[4\].row\[4\].yc/lin[0] blk.column\[4\].row\[4\].yc/lin[1]
+ blk.column\[5\].row\[4\].yc/rin[0] blk.column\[5\].row\[4\].yc/rin[1] blk.column\[3\].row\[4\].yc/hempty
+ blk.column\[4\].row\[4\].yc/reset blk.column\[4\].row\[5\].yc/reset blk.column\[4\].row\[4\].yc/rin[0]
+ blk.column\[4\].row\[4\].yc/rin[1] blk.column\[3\].row\[4\].yc/lin[0] blk.column\[3\].row\[4\].yc/lin[1]
+ blk.column\[4\].row\[4\].yc/uempty blk.column\[4\].row\[4\].yc/uin[0] blk.column\[4\].row\[4\].yc/uin[1]
+ blk.column\[4\].row\[3\].yc/din[0] blk.column\[4\].row\[3\].yc/din[1] blk.column\[4\].row\[3\].yc/dempty
+ blk.column\[4\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_537_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_368_ _780_/Q VGND VGND VPWR VPWR _368_/Y sky130_fd_sc_hd__inv_2
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xblk.column\[11\].row\[14\].yc blk.column\[11\].row\[14\].yc/cbitin blk.column\[11\].row\[15\].yc/cbitin
+ blk.column\[11\].row\[14\].yc/confclk blk.column\[11\].row\[15\].yc/confclk blk.column\[11\].row\[14\].yc/dempty
+ blk.column\[11\].row\[14\].yc/din[0] blk.column\[11\].row\[14\].yc/din[1] blk.column\[11\].row\[15\].yc/uin[0]
+ blk.column\[11\].row\[15\].yc/uin[1] blk.column\[11\].row\[14\].yc/hempty blk.column\[10\].row\[14\].yc/lempty
+ blk.column\[11\].row\[14\].yc/lempty blk.column\[11\].row\[14\].yc/lin[0] blk.column\[11\].row\[14\].yc/lin[1]
+ blk.column\[12\].row\[14\].yc/rin[0] blk.column\[12\].row\[14\].yc/rin[1] blk.column\[10\].row\[14\].yc/hempty
+ blk.column\[11\].row\[14\].yc/reset blk.column\[11\].row\[15\].yc/reset blk.column\[11\].row\[14\].yc/rin[0]
+ blk.column\[11\].row\[14\].yc/rin[1] blk.column\[10\].row\[14\].yc/lin[0] blk.column\[10\].row\[14\].yc/lin[1]
+ blk.column\[11\].row\[14\].yc/uempty blk.column\[11\].row\[14\].yc/uin[0] blk.column\[11\].row\[14\].yc/uin[1]
+ blk.column\[11\].row\[13\].yc/din[0] blk.column\[11\].row\[13\].yc/din[1] blk.column\[11\].row\[13\].yc/dempty
+ blk.column\[11\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_89_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_493_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_530_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_517_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_299_ _294_/Y _298_/X wbs_dat_i[7] _298_/X VGND VGND VPWR VPWR _299_/X sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_534_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_315_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_330_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_283_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_244_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_435_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_216_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_366_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_527_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_388_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_476_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_329_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_453_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_265_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_536_1804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[8\].row\[15\].yc blk.column\[8\].row\[15\].yc/cbitin la_data_out[40]
+ blk.column\[8\].row\[15\].yc/confclk blk.column\[8\].row\[15\].yc/confclko _474_/HI
+ _583_/LO _584_/LO blk.column\[8\].row\[15\].yc/dout[0] blk.column\[8\].row\[15\].yc/dout[1]
+ blk.column\[8\].row\[15\].yc/hempty blk.column\[7\].row\[15\].yc/lempty blk.column\[8\].row\[15\].yc/lempty
+ blk.column\[8\].row\[15\].yc/lin[0] blk.column\[8\].row\[15\].yc/lin[1] blk.column\[9\].row\[15\].yc/rin[0]
+ blk.column\[9\].row\[15\].yc/rin[1] blk.column\[7\].row\[15\].yc/hempty blk.column\[8\].row\[15\].yc/reset
+ blk.column\[8\].row\[15\].yc/reseto blk.column\[8\].row\[15\].yc/rin[0] blk.column\[8\].row\[15\].yc/rin[1]
+ blk.column\[7\].row\[15\].yc/lin[0] blk.column\[7\].row\[15\].yc/lin[1] blk.column\[8\].row\[15\].yc/uempty
+ blk.column\[8\].row\[15\].yc/uin[0] blk.column\[8\].row\[15\].yc/uin[1] blk.column\[8\].row\[14\].yc/din[0]
+ blk.column\[8\].row\[14\].yc/din[1] blk.column\[8\].row\[14\].yc/dempty blk.column\[8\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XFILLER_11_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_514_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_528_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_502_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_212_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_402_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_222_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_257_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_539_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_535_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_531_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_517_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_315_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_771_ wb_clk_i _388_/X VGND VGND VPWR VPWR wbs_dat_o[27] sky130_fd_sc_hd__dfxtp_4
XFILLER_247_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_331_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_230_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_396_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_531_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_332_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_513_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_345_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_221_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_510_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_493_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_460_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[14\].row\[5\].yc blk.column\[14\].row\[5\].yc/cbitin blk.column\[14\].row\[6\].yc/cbitin
+ blk.column\[14\].row\[5\].yc/confclk blk.column\[14\].row\[6\].yc/confclk blk.column\[14\].row\[5\].yc/dempty
+ blk.column\[14\].row\[5\].yc/din[0] blk.column\[14\].row\[5\].yc/din[1] blk.column\[14\].row\[6\].yc/uin[0]
+ blk.column\[14\].row\[6\].yc/uin[1] blk.column\[14\].row\[5\].yc/hempty blk.column\[13\].row\[5\].yc/lempty
+ blk.column\[14\].row\[5\].yc/lempty blk.column\[14\].row\[5\].yc/lin[0] blk.column\[14\].row\[5\].yc/lin[1]
+ blk.column\[15\].row\[5\].yc/rin[0] blk.column\[15\].row\[5\].yc/rin[1] blk.column\[13\].row\[5\].yc/hempty
+ blk.column\[14\].row\[5\].yc/reset blk.column\[14\].row\[6\].yc/reset blk.column\[14\].row\[5\].yc/rin[0]
+ blk.column\[14\].row\[5\].yc/rin[1] blk.column\[13\].row\[5\].yc/lin[0] blk.column\[13\].row\[5\].yc/lin[1]
+ blk.column\[14\].row\[5\].yc/uempty blk.column\[14\].row\[5\].yc/uin[0] blk.column\[14\].row\[5\].yc/uin[1]
+ blk.column\[14\].row\[4\].yc/din[0] blk.column\[14\].row\[4\].yc/din[1] blk.column\[14\].row\[4\].yc/dempty
+ blk.column\[14\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_314_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_530_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_754_ wb_clk_i _754_/D VGND VGND VPWR VPWR wbs_dat_o[10] sky130_fd_sc_hd__dfxtp_4
XPHY_7597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_451_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_344_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_685_ VGND VGND VPWR VPWR _685_/HI la_data_out[69] sky130_fd_sc_hd__conb_1
Xblk.column\[5\].row\[6\].yc blk.column\[5\].row\[6\].yc/cbitin blk.column\[5\].row\[7\].yc/cbitin
+ blk.column\[5\].row\[6\].yc/confclk blk.column\[5\].row\[7\].yc/confclk blk.column\[5\].row\[6\].yc/dempty
+ blk.column\[5\].row\[6\].yc/din[0] blk.column\[5\].row\[6\].yc/din[1] blk.column\[5\].row\[7\].yc/uin[0]
+ blk.column\[5\].row\[7\].yc/uin[1] blk.column\[5\].row\[6\].yc/hempty blk.column\[4\].row\[6\].yc/lempty
+ blk.column\[5\].row\[6\].yc/lempty blk.column\[5\].row\[6\].yc/lin[0] blk.column\[5\].row\[6\].yc/lin[1]
+ blk.column\[6\].row\[6\].yc/rin[0] blk.column\[6\].row\[6\].yc/rin[1] blk.column\[4\].row\[6\].yc/hempty
+ blk.column\[5\].row\[6\].yc/reset blk.column\[5\].row\[7\].yc/reset blk.column\[5\].row\[6\].yc/rin[0]
+ blk.column\[5\].row\[6\].yc/rin[1] blk.column\[4\].row\[6\].yc/lin[0] blk.column\[4\].row\[6\].yc/lin[1]
+ blk.column\[5\].row\[6\].yc/uempty blk.column\[5\].row\[6\].yc/uin[0] blk.column\[5\].row\[6\].yc/uin[1]
+ blk.column\[5\].row\[5\].yc/din[0] blk.column\[5\].row\[5\].yc/din[1] blk.column\[5\].row\[5\].yc/dempty
+ blk.column\[5\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_235_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_455_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_517_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_370_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_351_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_474_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_252_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_522_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_526_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_495_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_525_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_427_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_513_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_11508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_10807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_465_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_478_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_470_ VGND VGND VPWR VPWR _470_/HI _470_/LO sky130_fd_sc_hd__conb_1
XPHY_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_298_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_519_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_515_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_806_ wb_clk_i _806_/D VGND VGND VPWR VPWR _806_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_7372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_737_ VGND VGND VPWR VPWR _737_/HI la_data_out[121] sky130_fd_sc_hd__conb_1
XPHY_6682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_668_ VGND VGND VPWR VPWR _668_/HI la_data_out[52] sky130_fd_sc_hd__conb_1
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_539_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_412_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_599_ VGND VGND VPWR VPWR _599_/HI io_oeb[11] sky130_fd_sc_hd__conb_1
XFILLER_496_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_0 _338_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_522_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_511_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_440_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_503_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_328_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_516_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_497_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_522_ VGND VGND VPWR VPWR _522_/HI _522_/LO sky130_fd_sc_hd__conb_1
XPHY_5266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_453_ VGND VGND VPWR VPWR _453_/HI _453_/LO sky130_fd_sc_hd__conb_1
XFILLER_306_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_359_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_360_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_384_ _391_/A VGND VGND VPWR VPWR _384_/X sky130_fd_sc_hd__buf_2
XFILLER_13_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_532_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_313_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_429_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_498_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_253_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_424_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_299_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_295_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xblk.column\[15\].row\[7\].yc blk.column\[15\].row\[7\].yc/cbitin blk.column\[15\].row\[8\].yc/cbitin
+ blk.column\[15\].row\[7\].yc/confclk blk.column\[15\].row\[8\].yc/confclk blk.column\[15\].row\[7\].yc/dempty
+ blk.column\[15\].row\[7\].yc/din[0] blk.column\[15\].row\[7\].yc/din[1] blk.column\[15\].row\[8\].yc/uin[0]
+ blk.column\[15\].row\[8\].yc/uin[1] blk.column\[15\].row\[7\].yc/hempty blk.column\[14\].row\[7\].yc/lempty
+ _464_/HI _555_/LO _556_/LO blk.column\[15\].row\[7\].yc/lout[0] blk.column\[15\].row\[7\].yc/lout[1]
+ blk.column\[14\].row\[7\].yc/hempty blk.column\[15\].row\[7\].yc/reset blk.column\[15\].row\[8\].yc/reset
+ blk.column\[15\].row\[7\].yc/rin[0] blk.column\[15\].row\[7\].yc/rin[1] blk.column\[14\].row\[7\].yc/lin[0]
+ blk.column\[14\].row\[7\].yc/lin[1] blk.column\[15\].row\[7\].yc/uempty blk.column\[15\].row\[7\].yc/uin[0]
+ blk.column\[15\].row\[7\].yc/uin[1] blk.column\[15\].row\[6\].yc/din[0] blk.column\[15\].row\[6\].yc/din[1]
+ blk.column\[15\].row\[6\].yc/dempty blk.column\[15\].row\[8\].yc/uempty VPWR VGND
+ ycell
XFILLER_503_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_312_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_334_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_396_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[6\].row\[8\].yc blk.column\[6\].row\[8\].yc/cbitin blk.column\[6\].row\[9\].yc/cbitin
+ blk.column\[6\].row\[8\].yc/confclk blk.column\[6\].row\[9\].yc/confclk blk.column\[6\].row\[8\].yc/dempty
+ blk.column\[6\].row\[8\].yc/din[0] blk.column\[6\].row\[8\].yc/din[1] blk.column\[6\].row\[9\].yc/uin[0]
+ blk.column\[6\].row\[9\].yc/uin[1] blk.column\[6\].row\[8\].yc/hempty blk.column\[5\].row\[8\].yc/lempty
+ blk.column\[6\].row\[8\].yc/lempty blk.column\[6\].row\[8\].yc/lin[0] blk.column\[6\].row\[8\].yc/lin[1]
+ blk.column\[7\].row\[8\].yc/rin[0] blk.column\[7\].row\[8\].yc/rin[1] blk.column\[5\].row\[8\].yc/hempty
+ blk.column\[6\].row\[8\].yc/reset blk.column\[6\].row\[9\].yc/reset blk.column\[6\].row\[8\].yc/rin[0]
+ blk.column\[6\].row\[8\].yc/rin[1] blk.column\[5\].row\[8\].yc/lin[0] blk.column\[5\].row\[8\].yc/lin[1]
+ blk.column\[6\].row\[8\].yc/uempty blk.column\[6\].row\[8\].yc/uin[0] blk.column\[6\].row\[8\].yc/uin[1]
+ blk.column\[6\].row\[7\].yc/din[0] blk.column\[6\].row\[7\].yc/din[1] blk.column\[6\].row\[7\].yc/dempty
+ blk.column\[6\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_510_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_447_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_542_2927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_292_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_505_ VGND VGND VPWR VPWR _505_/HI _505_/LO sky130_fd_sc_hd__conb_1
XFILLER_505_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_436_ VGND VGND VPWR VPWR _436_/HI _436_/LO sky130_fd_sc_hd__conb_1
XPHY_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_399_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_367_ _365_/Y _361_/X wbs_dat_i[29] _366_/X VGND VGND VPWR VPWR _781_/D sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_534_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_298_ _298_/A VGND VGND VPWR VPWR _298_/X sky130_fd_sc_hd__buf_2
XFILLER_493_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_525_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_476_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_348_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_428_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_419_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_290_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_331_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_361_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_530_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_311_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_524_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_388_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_299_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_329_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_506_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_531_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_501_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_312_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_454_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_419_ _419_/A VGND VGND VPWR VPWR _419_/X sky130_fd_sc_hd__buf_2
XFILLER_11_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_509_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[10\].row\[0\].yc la_data_in[106] blk.column\[10\].row\[1\].yc/cbitin
+ la_data_in[112] blk.column\[10\].row\[1\].yc/confclk blk.column\[10\].row\[0\].yc/dempty
+ blk.column\[10\].row\[0\].yc/din[0] blk.column\[10\].row\[0\].yc/din[1] blk.column\[10\].row\[1\].yc/uin[0]
+ blk.column\[10\].row\[1\].yc/uin[1] blk.column\[10\].row\[0\].yc/hempty blk.column\[9\].row\[0\].yc/lempty
+ blk.column\[10\].row\[0\].yc/lempty blk.column\[10\].row\[0\].yc/lin[0] blk.column\[10\].row\[0\].yc/lin[1]
+ blk.column\[11\].row\[0\].yc/rin[0] blk.column\[11\].row\[0\].yc/rin[1] blk.column\[9\].row\[0\].yc/hempty
+ la_data_in[113] blk.column\[10\].row\[1\].yc/reset blk.column\[9\].row\[0\].yc/lout[0]
+ blk.column\[9\].row\[0\].yc/lout[1] blk.column\[9\].row\[0\].yc/lin[0] blk.column\[9\].row\[0\].yc/lin[1]
+ _511_/LO la_data_in[84] la_data_in[85] la_data_out[20] la_data_out[21] blk.column\[10\].row\[0\].yc/vempty
+ blk.column\[10\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_83_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_520_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_457_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_361_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[1\].yc blk.column\[1\].row\[1\].yc/cbitin blk.column\[1\].row\[2\].yc/cbitin
+ blk.column\[1\].row\[1\].yc/confclk blk.column\[1\].row\[2\].yc/confclk blk.column\[1\].row\[1\].yc/dempty
+ blk.column\[1\].row\[1\].yc/din[0] blk.column\[1\].row\[1\].yc/din[1] blk.column\[1\].row\[2\].yc/uin[0]
+ blk.column\[1\].row\[2\].yc/uin[1] blk.column\[1\].row\[1\].yc/hempty blk.column\[0\].row\[1\].yc/lempty
+ blk.column\[1\].row\[1\].yc/lempty blk.column\[1\].row\[1\].yc/lin[0] blk.column\[1\].row\[1\].yc/lin[1]
+ blk.column\[2\].row\[1\].yc/rin[0] blk.column\[2\].row\[1\].yc/rin[1] blk.column\[0\].row\[1\].yc/hempty
+ blk.column\[1\].row\[1\].yc/reset blk.column\[1\].row\[2\].yc/reset blk.column\[1\].row\[1\].yc/rin[0]
+ blk.column\[1\].row\[1\].yc/rin[1] blk.column\[0\].row\[1\].yc/lin[0] blk.column\[0\].row\[1\].yc/lin[1]
+ blk.column\[1\].row\[1\].yc/uempty blk.column\[1\].row\[1\].yc/uin[0] blk.column\[1\].row\[1\].yc/uin[1]
+ blk.column\[1\].row\[0\].yc/din[0] blk.column\[1\].row\[0\].yc/din[1] blk.column\[1\].row\[0\].yc/dempty
+ blk.column\[1\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_506_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_437_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_385_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_517_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_770_ wb_clk_i _770_/D VGND VGND VPWR VPWR wbs_dat_o[26] sky130_fd_sc_hd__dfxtp_4
XPHY_7757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_487_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_492_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[11\].yc blk.column\[5\].row\[11\].yc/cbitin blk.column\[5\].row\[12\].yc/cbitin
+ blk.column\[5\].row\[11\].yc/confclk blk.column\[5\].row\[12\].yc/confclk blk.column\[5\].row\[11\].yc/dempty
+ blk.column\[5\].row\[11\].yc/din[0] blk.column\[5\].row\[11\].yc/din[1] blk.column\[5\].row\[12\].yc/uin[0]
+ blk.column\[5\].row\[12\].yc/uin[1] blk.column\[5\].row\[11\].yc/hempty blk.column\[4\].row\[11\].yc/lempty
+ blk.column\[5\].row\[11\].yc/lempty blk.column\[5\].row\[11\].yc/lin[0] blk.column\[5\].row\[11\].yc/lin[1]
+ blk.column\[6\].row\[11\].yc/rin[0] blk.column\[6\].row\[11\].yc/rin[1] blk.column\[4\].row\[11\].yc/hempty
+ blk.column\[5\].row\[11\].yc/reset blk.column\[5\].row\[12\].yc/reset blk.column\[5\].row\[11\].yc/rin[0]
+ blk.column\[5\].row\[11\].yc/rin[1] blk.column\[4\].row\[11\].yc/lin[0] blk.column\[4\].row\[11\].yc/lin[1]
+ blk.column\[5\].row\[11\].yc/uempty blk.column\[5\].row\[11\].yc/uin[0] blk.column\[5\].row\[11\].yc/uin[1]
+ blk.column\[5\].row\[10\].yc/din[0] blk.column\[5\].row\[10\].yc/din[1] blk.column\[5\].row\[10\].yc/dempty
+ blk.column\[5\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_227_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_261_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_349_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_494_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_396_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_238_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_483_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_454_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_253_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_3037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_501_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_524_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_432_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_215_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_284_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_528_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_506_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_322_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_468_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_526_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_342_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_485_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_753_ wb_clk_i _753_/D VGND VGND VPWR VPWR wbs_dat_o[9] sky130_fd_sc_hd__dfxtp_4
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_524_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_684_ VGND VGND VPWR VPWR _684_/HI la_data_out[68] sky130_fd_sc_hd__conb_1
XPHY_6897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_349_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_519_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_518_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_509_2758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_525_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_503_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_332_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_503_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[12\].row\[13\].yc blk.column\[12\].row\[13\].yc/cbitin blk.column\[12\].row\[14\].yc/cbitin
+ blk.column\[12\].row\[13\].yc/confclk blk.column\[12\].row\[14\].yc/confclk blk.column\[12\].row\[13\].yc/dempty
+ blk.column\[12\].row\[13\].yc/din[0] blk.column\[12\].row\[13\].yc/din[1] blk.column\[12\].row\[14\].yc/uin[0]
+ blk.column\[12\].row\[14\].yc/uin[1] blk.column\[12\].row\[13\].yc/hempty blk.column\[11\].row\[13\].yc/lempty
+ blk.column\[12\].row\[13\].yc/lempty blk.column\[12\].row\[13\].yc/lin[0] blk.column\[12\].row\[13\].yc/lin[1]
+ blk.column\[13\].row\[13\].yc/rin[0] blk.column\[13\].row\[13\].yc/rin[1] blk.column\[11\].row\[13\].yc/hempty
+ blk.column\[12\].row\[13\].yc/reset blk.column\[12\].row\[14\].yc/reset blk.column\[12\].row\[13\].yc/rin[0]
+ blk.column\[12\].row\[13\].yc/rin[1] blk.column\[11\].row\[13\].yc/lin[0] blk.column\[11\].row\[13\].yc/lin[1]
+ blk.column\[12\].row\[13\].yc/uempty blk.column\[12\].row\[13\].yc/uin[0] blk.column\[12\].row\[13\].yc/uin[1]
+ blk.column\[12\].row\[12\].yc/din[0] blk.column\[12\].row\[12\].yc/din[1] blk.column\[12\].row\[12\].yc/dempty
+ blk.column\[12\].row\[14\].yc/uempty VPWR VGND ycell
XFILLER_526_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_497_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_480_3106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_386_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_465_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_217_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_517_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_337_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_532_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_503_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_353_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_310_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_805_ wb_clk_i _304_/X VGND VGND VPWR VPWR _805_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_248_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_526_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_736_ VGND VGND VPWR VPWR _736_/HI la_data_out[120] sky130_fd_sc_hd__conb_1
XFILLER_75_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_422_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_667_ VGND VGND VPWR VPWR _667_/HI la_data_out[51] sky130_fd_sc_hd__conb_1
XFILLER_524_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_598_ VGND VGND VPWR VPWR _598_/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XFILLER_496_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_378_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[2\].yc blk.column\[11\].row\[2\].yc/cbitin blk.column\[11\].row\[3\].yc/cbitin
+ blk.column\[11\].row\[2\].yc/confclk blk.column\[11\].row\[3\].yc/confclk blk.column\[11\].row\[2\].yc/dempty
+ blk.column\[11\].row\[2\].yc/din[0] blk.column\[11\].row\[2\].yc/din[1] blk.column\[11\].row\[3\].yc/uin[0]
+ blk.column\[11\].row\[3\].yc/uin[1] blk.column\[11\].row\[2\].yc/hempty blk.column\[10\].row\[2\].yc/lempty
+ blk.column\[11\].row\[2\].yc/lempty blk.column\[11\].row\[2\].yc/lin[0] blk.column\[11\].row\[2\].yc/lin[1]
+ blk.column\[12\].row\[2\].yc/rin[0] blk.column\[12\].row\[2\].yc/rin[1] blk.column\[10\].row\[2\].yc/hempty
+ blk.column\[11\].row\[2\].yc/reset blk.column\[11\].row\[3\].yc/reset blk.column\[11\].row\[2\].yc/rin[0]
+ blk.column\[11\].row\[2\].yc/rin[1] blk.column\[10\].row\[2\].yc/lin[0] blk.column\[10\].row\[2\].yc/lin[1]
+ blk.column\[11\].row\[2\].yc/uempty blk.column\[11\].row\[2\].yc/uin[0] blk.column\[11\].row\[2\].yc/uin[1]
+ blk.column\[11\].row\[1\].yc/din[0] blk.column\[11\].row\[1\].yc/din[1] blk.column\[11\].row\[1\].yc/dempty
+ blk.column\[11\].row\[3\].yc/uempty VPWR VGND ycell
XFILLER_520_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_479_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_301_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[3\].yc blk.column\[2\].row\[3\].yc/cbitin blk.column\[2\].row\[4\].yc/cbitin
+ blk.column\[2\].row\[3\].yc/confclk blk.column\[2\].row\[4\].yc/confclk blk.column\[2\].row\[3\].yc/dempty
+ blk.column\[2\].row\[3\].yc/din[0] blk.column\[2\].row\[3\].yc/din[1] blk.column\[2\].row\[4\].yc/uin[0]
+ blk.column\[2\].row\[4\].yc/uin[1] blk.column\[2\].row\[3\].yc/hempty blk.column\[1\].row\[3\].yc/lempty
+ blk.column\[2\].row\[3\].yc/lempty blk.column\[2\].row\[3\].yc/lin[0] blk.column\[2\].row\[3\].yc/lin[1]
+ blk.column\[3\].row\[3\].yc/rin[0] blk.column\[3\].row\[3\].yc/rin[1] blk.column\[1\].row\[3\].yc/hempty
+ blk.column\[2\].row\[3\].yc/reset blk.column\[2\].row\[4\].yc/reset blk.column\[2\].row\[3\].yc/rin[0]
+ blk.column\[2\].row\[3\].yc/rin[1] blk.column\[1\].row\[3\].yc/lin[0] blk.column\[1\].row\[3\].yc/lin[1]
+ blk.column\[2\].row\[3\].yc/uempty blk.column\[2\].row\[3\].yc/uin[0] blk.column\[2\].row\[3\].yc/uin[1]
+ blk.column\[2\].row\[2\].yc/din[0] blk.column\[2\].row\[2\].yc/din[1] blk.column\[2\].row\[2\].yc/dempty
+ blk.column\[2\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_7_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_447_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_462_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_214_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_520_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_368_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_438_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[14\].yc blk.column\[9\].row\[14\].yc/cbitin blk.column\[9\].row\[15\].yc/cbitin
+ blk.column\[9\].row\[14\].yc/confclk blk.column\[9\].row\[15\].yc/confclk blk.column\[9\].row\[14\].yc/dempty
+ blk.column\[9\].row\[14\].yc/din[0] blk.column\[9\].row\[14\].yc/din[1] blk.column\[9\].row\[15\].yc/uin[0]
+ blk.column\[9\].row\[15\].yc/uin[1] blk.column\[9\].row\[14\].yc/hempty blk.column\[8\].row\[14\].yc/lempty
+ blk.column\[9\].row\[14\].yc/lempty blk.column\[9\].row\[14\].yc/lin[0] blk.column\[9\].row\[14\].yc/lin[1]
+ blk.column\[9\].row\[14\].yc/lout[0] blk.column\[9\].row\[14\].yc/lout[1] blk.column\[8\].row\[14\].yc/hempty
+ blk.column\[9\].row\[14\].yc/reset blk.column\[9\].row\[15\].yc/reset blk.column\[9\].row\[14\].yc/rin[0]
+ blk.column\[9\].row\[14\].yc/rin[1] blk.column\[8\].row\[14\].yc/lin[0] blk.column\[8\].row\[14\].yc/lin[1]
+ blk.column\[9\].row\[14\].yc/uempty blk.column\[9\].row\[14\].yc/uin[0] blk.column\[9\].row\[14\].yc/uin[1]
+ blk.column\[9\].row\[13\].yc/din[0] blk.column\[9\].row\[13\].yc/din[1] blk.column\[9\].row\[13\].yc/dempty
+ blk.column\[9\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_328_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_500_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_534_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_2949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_470_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_445_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_265_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_521_ VGND VGND VPWR VPWR _521_/HI _521_/LO sky130_fd_sc_hd__conb_1
XFILLER_406_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_452_ VGND VGND VPWR VPWR _452_/HI _452_/LO sky130_fd_sc_hd__conb_1
XPHY_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_360_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_383_ wbs_dat_o[31] _391_/A _358_/A _382_/X VGND VGND VPWR VPWR _775_/D sky130_fd_sc_hd__o22a_4
XPHY_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_374_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_352_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_429_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_283_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_506_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_719_ VGND VGND VPWR VPWR _719_/HI la_data_out[103] sky130_fd_sc_hd__conb_1
XFILLER_480_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_504_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_365_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_475_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_249_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_440_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_475_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_503_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_538_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_516_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_431_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xblk.column\[0\].row\[12\].yc blk.column\[0\].row\[12\].yc/cbitin blk.column\[0\].row\[13\].yc/cbitin
+ blk.column\[0\].row\[12\].yc/confclk blk.column\[0\].row\[13\].yc/confclk blk.column\[0\].row\[12\].yc/dempty
+ blk.column\[0\].row\[12\].yc/din[0] blk.column\[0\].row\[12\].yc/din[1] blk.column\[0\].row\[13\].yc/uin[0]
+ blk.column\[0\].row\[13\].yc/uin[1] blk.column\[0\].row\[12\].yc/hempty blk.column\[0\].row\[12\].yc/hempty2
+ blk.column\[0\].row\[12\].yc/lempty blk.column\[0\].row\[12\].yc/lin[0] blk.column\[0\].row\[12\].yc/lin[1]
+ blk.column\[1\].row\[12\].yc/rin[0] blk.column\[1\].row\[12\].yc/rin[1] _431_/HI
+ blk.column\[0\].row\[12\].yc/reset blk.column\[0\].row\[13\].yc/reset _483_/LO _484_/LO
+ blk.column\[0\].row\[12\].yc/rout[0] blk.column\[0\].row\[12\].yc/rout[1] blk.column\[0\].row\[12\].yc/uempty
+ blk.column\[0\].row\[12\].yc/uin[0] blk.column\[0\].row\[12\].yc/uin[1] blk.column\[0\].row\[11\].yc/din[0]
+ blk.column\[0\].row\[11\].yc/din[1] blk.column\[0\].row\[11\].yc/dempty blk.column\[0\].row\[13\].yc/uempty
+ VPWR VGND ycell
XFILLER_312_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_11158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_426_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_482_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_480_2032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_504_ VGND VGND VPWR VPWR _504_/HI _504_/LO sky130_fd_sc_hd__conb_1
XPHY_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_430_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_505_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_504_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_435_ VGND VGND VPWR VPWR _435_/HI _435_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_366_ _361_/A VGND VGND VPWR VPWR _366_/X sky130_fd_sc_hd__buf_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_536_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_509_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_347_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_538_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_297_ _297_/A VGND VGND VPWR VPWR _298_/A sky130_fd_sc_hd__buf_2
XFILLER_13_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_541_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_228_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_428_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_397_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_361_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_321_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_259_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_451_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_408_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_509_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_446_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_522_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_250_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_303_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_396_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_476_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_527_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_516_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_361_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_454_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_361_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_425_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_308_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[4\].yc blk.column\[12\].row\[4\].yc/cbitin blk.column\[12\].row\[5\].yc/cbitin
+ blk.column\[12\].row\[4\].yc/confclk blk.column\[12\].row\[5\].yc/confclk blk.column\[12\].row\[4\].yc/dempty
+ blk.column\[12\].row\[4\].yc/din[0] blk.column\[12\].row\[4\].yc/din[1] blk.column\[12\].row\[5\].yc/uin[0]
+ blk.column\[12\].row\[5\].yc/uin[1] blk.column\[12\].row\[4\].yc/hempty blk.column\[11\].row\[4\].yc/lempty
+ blk.column\[12\].row\[4\].yc/lempty blk.column\[12\].row\[4\].yc/lin[0] blk.column\[12\].row\[4\].yc/lin[1]
+ blk.column\[13\].row\[4\].yc/rin[0] blk.column\[13\].row\[4\].yc/rin[1] blk.column\[11\].row\[4\].yc/hempty
+ blk.column\[12\].row\[4\].yc/reset blk.column\[12\].row\[5\].yc/reset blk.column\[12\].row\[4\].yc/rin[0]
+ blk.column\[12\].row\[4\].yc/rin[1] blk.column\[11\].row\[4\].yc/lin[0] blk.column\[11\].row\[4\].yc/lin[1]
+ blk.column\[12\].row\[4\].yc/uempty blk.column\[12\].row\[4\].yc/uin[0] blk.column\[12\].row\[4\].yc/uin[1]
+ blk.column\[12\].row\[3\].yc/din[0] blk.column\[12\].row\[3\].yc/din[1] blk.column\[12\].row\[3\].yc/dempty
+ blk.column\[12\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_501_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_379_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_523_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_477_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_419_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_418_ _412_/X wbs_dat_o[6] _806_/Q _417_/X VGND VGND VPWR VPWR _418_/X sky130_fd_sc_hd__o22a_4
XFILLER_499_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_497_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_438_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_349_ _349_/A VGND VGND VPWR VPWR _349_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[5\].yc blk.column\[3\].row\[5\].yc/cbitin blk.column\[3\].row\[6\].yc/cbitin
+ blk.column\[3\].row\[5\].yc/confclk blk.column\[3\].row\[6\].yc/confclk blk.column\[3\].row\[5\].yc/dempty
+ blk.column\[3\].row\[5\].yc/din[0] blk.column\[3\].row\[5\].yc/din[1] blk.column\[3\].row\[6\].yc/uin[0]
+ blk.column\[3\].row\[6\].yc/uin[1] blk.column\[3\].row\[5\].yc/hempty blk.column\[2\].row\[5\].yc/lempty
+ blk.column\[3\].row\[5\].yc/lempty blk.column\[3\].row\[5\].yc/lin[0] blk.column\[3\].row\[5\].yc/lin[1]
+ blk.column\[4\].row\[5\].yc/rin[0] blk.column\[4\].row\[5\].yc/rin[1] blk.column\[2\].row\[5\].yc/hempty
+ blk.column\[3\].row\[5\].yc/reset blk.column\[3\].row\[6\].yc/reset blk.column\[3\].row\[5\].yc/rin[0]
+ blk.column\[3\].row\[5\].yc/rin[1] blk.column\[2\].row\[5\].yc/lin[0] blk.column\[2\].row\[5\].yc/lin[1]
+ blk.column\[3\].row\[5\].yc/uempty blk.column\[3\].row\[5\].yc/uin[0] blk.column\[3\].row\[5\].yc/uin[1]
+ blk.column\[3\].row\[4\].yc/din[0] blk.column\[3\].row\[4\].yc/din[1] blk.column\[3\].row\[4\].yc/dempty
+ blk.column\[3\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_534_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_343_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_246_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_326_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_501_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_506_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_437_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_239_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_389_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_302_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_2356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_411_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_502_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_357_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_518_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_396_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_418_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_356_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_325_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_297_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_333_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_285_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_509_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_349_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_425_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_399_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_321_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_245_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_321_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_301_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_252_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_332_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_528_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[15\].yc blk.column\[4\].row\[15\].yc/cbitin la_data_out[36]
+ blk.column\[4\].row\[15\].yc/confclk blk.column\[4\].row\[15\].yc/confclko _470_/HI
+ _571_/LO _572_/LO blk.column\[4\].row\[15\].yc/dout[0] blk.column\[4\].row\[15\].yc/dout[1]
+ blk.column\[4\].row\[15\].yc/hempty blk.column\[3\].row\[15\].yc/lempty blk.column\[4\].row\[15\].yc/lempty
+ blk.column\[4\].row\[15\].yc/lin[0] blk.column\[4\].row\[15\].yc/lin[1] blk.column\[5\].row\[15\].yc/rin[0]
+ blk.column\[5\].row\[15\].yc/rin[1] blk.column\[3\].row\[15\].yc/hempty blk.column\[4\].row\[15\].yc/reset
+ blk.column\[4\].row\[15\].yc/reseto blk.column\[4\].row\[15\].yc/rin[0] blk.column\[4\].row\[15\].yc/rin[1]
+ blk.column\[3\].row\[15\].yc/lin[0] blk.column\[3\].row\[15\].yc/lin[1] blk.column\[4\].row\[15\].yc/uempty
+ blk.column\[4\].row\[15\].yc/uin[0] blk.column\[4\].row\[15\].yc/uin[1] blk.column\[4\].row\[14\].yc/din[0]
+ blk.column\[4\].row\[14\].yc/din[1] blk.column\[4\].row\[14\].yc/dempty blk.column\[4\].row\[15\].yc/vempty2
+ VPWR VGND ycell
XPHY_4907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_541_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_519_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_752_ wb_clk_i _752_/D VGND VGND VPWR VPWR wbs_dat_o[8] sky130_fd_sc_hd__dfxtp_4
XPHY_7577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_469_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_683_ VGND VGND VPWR VPWR _683_/HI la_data_out[67] sky130_fd_sc_hd__conb_1
XFILLER_508_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_483_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_379_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_538_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_372_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_515_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_511_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_286_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_299_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_536_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_236_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_287_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_367_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_3118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_386_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_341_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_224_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[13\].row\[6\].yc blk.column\[13\].row\[6\].yc/cbitin blk.column\[13\].row\[7\].yc/cbitin
+ blk.column\[13\].row\[6\].yc/confclk blk.column\[13\].row\[7\].yc/confclk blk.column\[13\].row\[6\].yc/dempty
+ blk.column\[13\].row\[6\].yc/din[0] blk.column\[13\].row\[6\].yc/din[1] blk.column\[13\].row\[7\].yc/uin[0]
+ blk.column\[13\].row\[7\].yc/uin[1] blk.column\[13\].row\[6\].yc/hempty blk.column\[12\].row\[6\].yc/lempty
+ blk.column\[13\].row\[6\].yc/lempty blk.column\[13\].row\[6\].yc/lin[0] blk.column\[13\].row\[6\].yc/lin[1]
+ blk.column\[14\].row\[6\].yc/rin[0] blk.column\[14\].row\[6\].yc/rin[1] blk.column\[12\].row\[6\].yc/hempty
+ blk.column\[13\].row\[6\].yc/reset blk.column\[13\].row\[7\].yc/reset blk.column\[13\].row\[6\].yc/rin[0]
+ blk.column\[13\].row\[6\].yc/rin[1] blk.column\[12\].row\[6\].yc/lin[0] blk.column\[12\].row\[6\].yc/lin[1]
+ blk.column\[13\].row\[6\].yc/uempty blk.column\[13\].row\[6\].yc/uin[0] blk.column\[13\].row\[6\].yc/uin[1]
+ blk.column\[13\].row\[5\].yc/din[0] blk.column\[13\].row\[5\].yc/din[1] blk.column\[13\].row\[5\].yc/dempty
+ blk.column\[13\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_510_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_267_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_804_ wb_clk_i _306_/X VGND VGND VPWR VPWR _305_/A sky130_fd_sc_hd__dfxtp_4
XPHY_8097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_346_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_735_ VGND VGND VPWR VPWR _735_/HI la_data_out[119] sky130_fd_sc_hd__conb_1
XFILLER_507_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_263_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_666_ VGND VGND VPWR VPWR _666_/HI la_data_out[50] sky130_fd_sc_hd__conb_1
XFILLER_1_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_441_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_597_ VGND VGND VPWR VPWR _597_/HI io_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_539_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[4\].row\[7\].yc blk.column\[4\].row\[7\].yc/cbitin blk.column\[4\].row\[8\].yc/cbitin
+ blk.column\[4\].row\[7\].yc/confclk blk.column\[4\].row\[8\].yc/confclk blk.column\[4\].row\[7\].yc/dempty
+ blk.column\[4\].row\[7\].yc/din[0] blk.column\[4\].row\[7\].yc/din[1] blk.column\[4\].row\[8\].yc/uin[0]
+ blk.column\[4\].row\[8\].yc/uin[1] blk.column\[4\].row\[7\].yc/hempty blk.column\[3\].row\[7\].yc/lempty
+ blk.column\[4\].row\[7\].yc/lempty blk.column\[4\].row\[7\].yc/lin[0] blk.column\[4\].row\[7\].yc/lin[1]
+ blk.column\[5\].row\[7\].yc/rin[0] blk.column\[5\].row\[7\].yc/rin[1] blk.column\[3\].row\[7\].yc/hempty
+ blk.column\[4\].row\[7\].yc/reset blk.column\[4\].row\[8\].yc/reset blk.column\[4\].row\[7\].yc/rin[0]
+ blk.column\[4\].row\[7\].yc/rin[1] blk.column\[3\].row\[7\].yc/lin[0] blk.column\[3\].row\[7\].yc/lin[1]
+ blk.column\[4\].row\[7\].yc/uempty blk.column\[4\].row\[7\].yc/uin[0] blk.column\[4\].row\[7\].yc/uin[1]
+ blk.column\[4\].row\[6\].yc/din[0] blk.column\[4\].row\[6\].yc/din[1] blk.column\[4\].row\[6\].yc/dempty
+ blk.column\[4\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_378_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_318_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_508_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_518_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_503_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_415_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_516_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_495_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_513_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_249_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_264_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_520_ VGND VGND VPWR VPWR _520_/HI _520_/LO sky130_fd_sc_hd__conb_1
XFILLER_527_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_451_ VGND VGND VPWR VPWR _451_/HI _451_/LO sky130_fd_sc_hd__conb_1
XPHY_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_382_ _382_/A VGND VGND VPWR VPWR _382_/X sky130_fd_sc_hd__buf_2
XFILLER_496_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_348_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_536_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[9\].row\[1\].yc blk.column\[9\].row\[1\].yc/cbitin blk.column\[9\].row\[2\].yc/cbitin
+ blk.column\[9\].row\[1\].yc/confclk blk.column\[9\].row\[2\].yc/confclk blk.column\[9\].row\[1\].yc/dempty
+ blk.column\[9\].row\[1\].yc/din[0] blk.column\[9\].row\[1\].yc/din[1] blk.column\[9\].row\[2\].yc/uin[0]
+ blk.column\[9\].row\[2\].yc/uin[1] blk.column\[9\].row\[1\].yc/hempty blk.column\[8\].row\[1\].yc/lempty
+ blk.column\[9\].row\[1\].yc/lempty blk.column\[9\].row\[1\].yc/lin[0] blk.column\[9\].row\[1\].yc/lin[1]
+ blk.column\[9\].row\[1\].yc/lout[0] blk.column\[9\].row\[1\].yc/lout[1] blk.column\[8\].row\[1\].yc/hempty
+ blk.column\[9\].row\[1\].yc/reset blk.column\[9\].row\[2\].yc/reset blk.column\[9\].row\[1\].yc/rin[0]
+ blk.column\[9\].row\[1\].yc/rin[1] blk.column\[8\].row\[1\].yc/lin[0] blk.column\[8\].row\[1\].yc/lin[1]
+ blk.column\[9\].row\[1\].yc/uempty blk.column\[9\].row\[1\].yc/uin[0] blk.column\[9\].row\[1\].yc/uin[1]
+ blk.column\[9\].row\[0\].yc/din[0] blk.column\[9\].row\[0\].yc/din[1] blk.column\[9\].row\[0\].yc/dempty
+ blk.column\[9\].row\[2\].yc/uempty VPWR VGND ycell
XFILLER_185_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_491_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_519_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_534_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[6\].row\[10\].yc blk.column\[6\].row\[9\].yc/cbitout blk.column\[6\].row\[11\].yc/cbitin
+ blk.column\[6\].row\[9\].yc/confclko blk.column\[6\].row\[11\].yc/confclk blk.column\[6\].row\[10\].yc/dempty
+ blk.column\[6\].row\[10\].yc/din[0] blk.column\[6\].row\[10\].yc/din[1] blk.column\[6\].row\[11\].yc/uin[0]
+ blk.column\[6\].row\[11\].yc/uin[1] blk.column\[6\].row\[10\].yc/hempty blk.column\[5\].row\[10\].yc/lempty
+ blk.column\[6\].row\[10\].yc/lempty blk.column\[6\].row\[10\].yc/lin[0] blk.column\[6\].row\[10\].yc/lin[1]
+ blk.column\[7\].row\[10\].yc/rin[0] blk.column\[7\].row\[10\].yc/rin[1] blk.column\[5\].row\[10\].yc/hempty
+ blk.column\[6\].row\[9\].yc/reseto blk.column\[6\].row\[11\].yc/reset blk.column\[6\].row\[10\].yc/rin[0]
+ blk.column\[6\].row\[10\].yc/rin[1] blk.column\[5\].row\[10\].yc/lin[0] blk.column\[5\].row\[10\].yc/lin[1]
+ blk.column\[6\].row\[9\].yc/vempty2 blk.column\[6\].row\[9\].yc/dout[0] blk.column\[6\].row\[9\].yc/dout[1]
+ blk.column\[6\].row\[9\].yc/din[0] blk.column\[6\].row\[9\].yc/din[1] blk.column\[6\].row\[9\].yc/dempty
+ blk.column\[6\].row\[11\].yc/uempty VPWR VGND ycell
XPHY_7171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_460_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_718_ VGND VGND VPWR VPWR _718_/HI la_data_out[102] sky130_fd_sc_hd__conb_1
XPHY_6492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_324_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_649_ VGND VGND VPWR VPWR _649_/HI io_out[23] sky130_fd_sc_hd__conb_1
XPHY_5791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_496_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_496_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_365_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_523_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_479_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_325_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_383_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_370_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_260_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_396_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_449_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_295_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_538_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_516_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_320_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_510_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_382_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_280_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_434_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_451_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_423_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_2077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_503_ VGND VGND VPWR VPWR _503_/HI _503_/LO sky130_fd_sc_hd__conb_1
XPHY_5087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_359_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_434_ VGND VGND VPWR VPWR _434_/HI _434_/LO sky130_fd_sc_hd__conb_1
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_365_ _365_/A VGND VGND VPWR VPWR _365_/Y sky130_fd_sc_hd__inv_2
XPHY_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_347_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_296_ _295_/Y wbs_we_i wbs_sel_i[0] VGND VGND VPWR VPWR _297_/A sky130_fd_sc_hd__and3_4
XFILLER_517_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_510_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_387_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_457_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_268_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_248_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_251_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_400_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_269_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_398_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_290_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_350_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_2685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_491_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_502_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_505_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_377_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xblk.column\[13\].row\[12\].yc blk.column\[13\].row\[12\].yc/cbitin blk.column\[13\].row\[13\].yc/cbitin
+ blk.column\[13\].row\[12\].yc/confclk blk.column\[13\].row\[13\].yc/confclk blk.column\[13\].row\[12\].yc/dempty
+ blk.column\[13\].row\[12\].yc/din[0] blk.column\[13\].row\[12\].yc/din[1] blk.column\[13\].row\[13\].yc/uin[0]
+ blk.column\[13\].row\[13\].yc/uin[1] blk.column\[13\].row\[12\].yc/hempty blk.column\[12\].row\[12\].yc/lempty
+ blk.column\[13\].row\[12\].yc/lempty blk.column\[13\].row\[12\].yc/lin[0] blk.column\[13\].row\[12\].yc/lin[1]
+ blk.column\[14\].row\[12\].yc/rin[0] blk.column\[14\].row\[12\].yc/rin[1] blk.column\[12\].row\[12\].yc/hempty
+ blk.column\[13\].row\[12\].yc/reset blk.column\[13\].row\[13\].yc/reset blk.column\[13\].row\[12\].yc/rin[0]
+ blk.column\[13\].row\[12\].yc/rin[1] blk.column\[12\].row\[12\].yc/lin[0] blk.column\[12\].row\[12\].yc/lin[1]
+ blk.column\[13\].row\[12\].yc/uempty blk.column\[13\].row\[12\].yc/uin[0] blk.column\[13\].row\[12\].yc/uin[1]
+ blk.column\[13\].row\[11\].yc/din[0] blk.column\[13\].row\[11\].yc/din[1] blk.column\[13\].row\[11\].yc/dempty
+ blk.column\[13\].row\[13\].yc/uempty VPWR VGND ycell
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_230_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_497_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_338_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_273_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_344_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[14\].row\[8\].yc blk.column\[14\].row\[8\].yc/cbitin blk.column\[14\].row\[9\].yc/cbitin
+ blk.column\[14\].row\[8\].yc/confclk blk.column\[14\].row\[9\].yc/confclk blk.column\[14\].row\[8\].yc/dempty
+ blk.column\[14\].row\[8\].yc/din[0] blk.column\[14\].row\[8\].yc/din[1] blk.column\[14\].row\[9\].yc/uin[0]
+ blk.column\[14\].row\[9\].yc/uin[1] blk.column\[14\].row\[8\].yc/hempty blk.column\[13\].row\[8\].yc/lempty
+ blk.column\[14\].row\[8\].yc/lempty blk.column\[14\].row\[8\].yc/lin[0] blk.column\[14\].row\[8\].yc/lin[1]
+ blk.column\[15\].row\[8\].yc/rin[0] blk.column\[15\].row\[8\].yc/rin[1] blk.column\[13\].row\[8\].yc/hempty
+ blk.column\[14\].row\[8\].yc/reset blk.column\[14\].row\[9\].yc/reset blk.column\[14\].row\[8\].yc/rin[0]
+ blk.column\[14\].row\[8\].yc/rin[1] blk.column\[13\].row\[8\].yc/lin[0] blk.column\[13\].row\[8\].yc/lin[1]
+ blk.column\[14\].row\[8\].yc/uempty blk.column\[14\].row\[8\].yc/uin[0] blk.column\[14\].row\[8\].yc/uin[1]
+ blk.column\[14\].row\[7\].yc/din[0] blk.column\[14\].row\[7\].yc/din[1] blk.column\[14\].row\[7\].yc/dempty
+ blk.column\[14\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_534_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_502_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_439_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_361_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_425_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_308_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[9\].yc blk.column\[5\].row\[9\].yc/cbitin blk.column\[5\].row\[9\].yc/cbitout
+ blk.column\[5\].row\[9\].yc/confclk blk.column\[5\].row\[9\].yc/confclko blk.column\[5\].row\[9\].yc/dempty
+ blk.column\[5\].row\[9\].yc/din[0] blk.column\[5\].row\[9\].yc/din[1] blk.column\[5\].row\[9\].yc/dout[0]
+ blk.column\[5\].row\[9\].yc/dout[1] blk.column\[5\].row\[9\].yc/hempty blk.column\[4\].row\[9\].yc/lempty
+ blk.column\[5\].row\[9\].yc/lempty blk.column\[5\].row\[9\].yc/lin[0] blk.column\[5\].row\[9\].yc/lin[1]
+ blk.column\[6\].row\[9\].yc/rin[0] blk.column\[6\].row\[9\].yc/rin[1] blk.column\[4\].row\[9\].yc/hempty
+ blk.column\[5\].row\[9\].yc/reset blk.column\[5\].row\[9\].yc/reseto blk.column\[5\].row\[9\].yc/rin[0]
+ blk.column\[5\].row\[9\].yc/rin[1] blk.column\[4\].row\[9\].yc/lin[0] blk.column\[4\].row\[9\].yc/lin[1]
+ blk.column\[5\].row\[9\].yc/uempty blk.column\[5\].row\[9\].yc/uin[0] blk.column\[5\].row\[9\].yc/uin[1]
+ blk.column\[5\].row\[8\].yc/din[0] blk.column\[5\].row\[8\].yc/din[1] blk.column\[5\].row\[8\].yc/dempty
+ blk.column\[5\].row\[9\].yc/vempty2 VPWR VGND ycell
XFILLER_265_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_379_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_458_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_394_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_417_ wb_rst_i VGND VGND VPWR VPWR _417_/X sky130_fd_sc_hd__buf_2
XFILLER_19_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_501_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_375_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_348_ _347_/Y _345_/X wbs_dat_i[20] _345_/X VGND VGND VPWR VPWR _788_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_386_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_536_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_315_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_517_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_255_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_271_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_457_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_3125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_460_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_1666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_212_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_496_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_446_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_326_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_381_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_333_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_524_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_462_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_463_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_420_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_522_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_519_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_507_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_414_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_356_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_418_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_529_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_300_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_388_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_305_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_454_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_2512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_284_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_442_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_507_1953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_261_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_395_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_493_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_266_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_525_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_436_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_291_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_252_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_346_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_282_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_477_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_445_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_2142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_443_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_506_1496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[0\].row\[2\].yc blk.column\[0\].row\[2\].yc/cbitin blk.column\[0\].row\[3\].yc/cbitin
+ blk.column\[0\].row\[2\].yc/confclk blk.column\[0\].row\[3\].yc/confclk blk.column\[0\].row\[2\].yc/dempty
+ blk.column\[0\].row\[2\].yc/din[0] blk.column\[0\].row\[2\].yc/din[1] blk.column\[0\].row\[3\].yc/uin[0]
+ blk.column\[0\].row\[3\].yc/uin[1] blk.column\[0\].row\[2\].yc/hempty blk.column\[0\].row\[2\].yc/hempty2
+ blk.column\[0\].row\[2\].yc/lempty blk.column\[0\].row\[2\].yc/lin[0] blk.column\[0\].row\[2\].yc/lin[1]
+ blk.column\[1\].row\[2\].yc/rin[0] blk.column\[1\].row\[2\].yc/rin[1] _437_/HI blk.column\[0\].row\[2\].yc/reset
+ blk.column\[0\].row\[3\].yc/reset _495_/LO _496_/LO blk.column\[0\].row\[2\].yc/rout[0]
+ blk.column\[0\].row\[2\].yc/rout[1] blk.column\[0\].row\[2\].yc/uempty blk.column\[0\].row\[2\].yc/uin[0]
+ blk.column\[0\].row\[2\].yc/uin[1] blk.column\[0\].row\[1\].yc/din[0] blk.column\[0\].row\[1\].yc/din[1]
+ blk.column\[0\].row\[1\].yc/dempty blk.column\[0\].row\[3\].yc/uempty VPWR VGND
+ ycell
XFILLER_519_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_296_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_354_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_532_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_489_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_279_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_512_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_513_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_409_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_751_ wb_clk_i _416_/X VGND VGND VPWR VPWR wbs_dat_o[7] sky130_fd_sc_hd__dfxtp_4
XFILLER_125_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_428_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_682_ VGND VGND VPWR VPWR _682_/HI la_data_out[66] sky130_fd_sc_hd__conb_1
XPHY_6877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_383_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_424_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_344_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_537_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_367_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_494_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_236_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_345_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_316_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_522_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[11\].yc blk.column\[1\].row\[11\].yc/cbitin blk.column\[1\].row\[12\].yc/cbitin
+ blk.column\[1\].row\[11\].yc/confclk blk.column\[1\].row\[12\].yc/confclk blk.column\[1\].row\[11\].yc/dempty
+ blk.column\[1\].row\[11\].yc/din[0] blk.column\[1\].row\[11\].yc/din[1] blk.column\[1\].row\[12\].yc/uin[0]
+ blk.column\[1\].row\[12\].yc/uin[1] blk.column\[1\].row\[11\].yc/hempty blk.column\[0\].row\[11\].yc/lempty
+ blk.column\[1\].row\[11\].yc/lempty blk.column\[1\].row\[11\].yc/lin[0] blk.column\[1\].row\[11\].yc/lin[1]
+ blk.column\[2\].row\[11\].yc/rin[0] blk.column\[2\].row\[11\].yc/rin[1] blk.column\[0\].row\[11\].yc/hempty
+ blk.column\[1\].row\[11\].yc/reset blk.column\[1\].row\[12\].yc/reset blk.column\[1\].row\[11\].yc/rin[0]
+ blk.column\[1\].row\[11\].yc/rin[1] blk.column\[0\].row\[11\].yc/lin[0] blk.column\[0\].row\[11\].yc/lin[1]
+ blk.column\[1\].row\[11\].yc/uempty blk.column\[1\].row\[11\].yc/uin[0] blk.column\[1\].row\[11\].yc/uin[1]
+ blk.column\[1\].row\[10\].yc/din[0] blk.column\[1\].row\[10\].yc/din[1] blk.column\[1\].row\[10\].yc/dempty
+ blk.column\[1\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_474_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_427_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_427_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_3032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_529_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_241_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_229_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_538_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_277_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_541_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_540_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_443_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_276_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_257_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2040 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_282_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_225_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_240_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_519_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_299_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_417_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_353_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_532_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_330_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_481_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_803_ wb_clk_i _308_/X VGND VGND VPWR VPWR _307_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_381_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_471_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_275_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_734_ VGND VGND VPWR VPWR _734_/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_208_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_290_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_665_ VGND VGND VPWR VPWR _665_/HI la_data_out[49] sky130_fd_sc_hd__conb_1
XFILLER_5_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_596_ VGND VGND VPWR VPWR _596_/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_504_2679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_441_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_441_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_458_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_392_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_537_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_298_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_2123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_542_2183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_411_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_503_1477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_293_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_391_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_541_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_369_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_494_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_438_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_534_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_230_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_2569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_453_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_486_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_272_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_403_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_380_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_527_1989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_525_2392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_450_ VGND VGND VPWR VPWR _450_/HI _450_/LO sky130_fd_sc_hd__conb_1
XPHY_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_2977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_341_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_414_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_381_ wb_rst_i VGND VGND VPWR VPWR _382_/A sky130_fd_sc_hd__buf_2
XPHY_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_421_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_538_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_364_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_444_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_437_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_244_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_717_ VGND VGND VPWR VPWR _717_/HI la_data_out[101] sky130_fd_sc_hd__conb_1
XFILLER_127_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_452_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_500_3008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_412_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_397_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_648_ VGND VGND VPWR VPWR _648_/HI io_out[22] sky130_fd_sc_hd__conb_1
XPHY_5792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_226_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_579_ VGND VGND VPWR VPWR _579_/HI _579_/LO sky130_fd_sc_hd__conb_1
XFILLER_18_2655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[10\].row\[3\].yc blk.column\[10\].row\[3\].yc/cbitin blk.column\[10\].row\[4\].yc/cbitin
+ blk.column\[10\].row\[3\].yc/confclk blk.column\[10\].row\[4\].yc/confclk blk.column\[10\].row\[3\].yc/dempty
+ blk.column\[10\].row\[3\].yc/din[0] blk.column\[10\].row\[3\].yc/din[1] blk.column\[10\].row\[4\].yc/uin[0]
+ blk.column\[10\].row\[4\].yc/uin[1] blk.column\[10\].row\[3\].yc/hempty blk.column\[9\].row\[3\].yc/lempty
+ blk.column\[10\].row\[3\].yc/lempty blk.column\[10\].row\[3\].yc/lin[0] blk.column\[10\].row\[3\].yc/lin[1]
+ blk.column\[11\].row\[3\].yc/rin[0] blk.column\[11\].row\[3\].yc/rin[1] blk.column\[9\].row\[3\].yc/hempty
+ blk.column\[10\].row\[3\].yc/reset blk.column\[10\].row\[4\].yc/reset blk.column\[9\].row\[3\].yc/lout[0]
+ blk.column\[9\].row\[3\].yc/lout[1] blk.column\[9\].row\[3\].yc/lin[0] blk.column\[9\].row\[3\].yc/lin[1]
+ blk.column\[10\].row\[3\].yc/uempty blk.column\[10\].row\[3\].yc/uin[0] blk.column\[10\].row\[3\].yc/uin[1]
+ blk.column\[10\].row\[2\].yc/din[0] blk.column\[10\].row\[2\].yc/din[1] blk.column\[10\].row\[2\].yc/dempty
+ blk.column\[10\].row\[4\].yc/uempty VPWR VGND ycell
XFILLER_138_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_511_3148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_214_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_435_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_364_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_329_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[1\].row\[4\].yc blk.column\[1\].row\[4\].yc/cbitin blk.column\[1\].row\[5\].yc/cbitin
+ blk.column\[1\].row\[4\].yc/confclk blk.column\[1\].row\[5\].yc/confclk blk.column\[1\].row\[4\].yc/dempty
+ blk.column\[1\].row\[4\].yc/din[0] blk.column\[1\].row\[4\].yc/din[1] blk.column\[1\].row\[5\].yc/uin[0]
+ blk.column\[1\].row\[5\].yc/uin[1] blk.column\[1\].row\[4\].yc/hempty blk.column\[0\].row\[4\].yc/lempty
+ blk.column\[1\].row\[4\].yc/lempty blk.column\[1\].row\[4\].yc/lin[0] blk.column\[1\].row\[4\].yc/lin[1]
+ blk.column\[2\].row\[4\].yc/rin[0] blk.column\[2\].row\[4\].yc/rin[1] blk.column\[0\].row\[4\].yc/hempty
+ blk.column\[1\].row\[4\].yc/reset blk.column\[1\].row\[5\].yc/reset blk.column\[1\].row\[4\].yc/rin[0]
+ blk.column\[1\].row\[4\].yc/rin[1] blk.column\[0\].row\[4\].yc/lin[0] blk.column\[0\].row\[4\].yc/lin[1]
+ blk.column\[1\].row\[4\].yc/uempty blk.column\[1\].row\[4\].yc/uin[0] blk.column\[1\].row\[4\].yc/uin[1]
+ blk.column\[1\].row\[3\].yc/din[0] blk.column\[1\].row\[3\].yc/din[1] blk.column\[1\].row\[3\].yc/dempty
+ blk.column\[1\].row\[5\].yc/uempty VPWR VGND ycell
XFILLER_23_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_1867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_424_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_479_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_449_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_500_2874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_356_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_320_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_371_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_2325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_470_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_412_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_431_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_232_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_514_2093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_264_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[5\].row\[14\].yc blk.column\[5\].row\[14\].yc/cbitin blk.column\[5\].row\[15\].yc/cbitin
+ blk.column\[5\].row\[14\].yc/confclk blk.column\[5\].row\[15\].yc/confclk blk.column\[5\].row\[14\].yc/dempty
+ blk.column\[5\].row\[14\].yc/din[0] blk.column\[5\].row\[14\].yc/din[1] blk.column\[5\].row\[15\].yc/uin[0]
+ blk.column\[5\].row\[15\].yc/uin[1] blk.column\[5\].row\[14\].yc/hempty blk.column\[4\].row\[14\].yc/lempty
+ blk.column\[5\].row\[14\].yc/lempty blk.column\[5\].row\[14\].yc/lin[0] blk.column\[5\].row\[14\].yc/lin[1]
+ blk.column\[6\].row\[14\].yc/rin[0] blk.column\[6\].row\[14\].yc/rin[1] blk.column\[4\].row\[14\].yc/hempty
+ blk.column\[5\].row\[14\].yc/reset blk.column\[5\].row\[15\].yc/reset blk.column\[5\].row\[14\].yc/rin[0]
+ blk.column\[5\].row\[14\].yc/rin[1] blk.column\[4\].row\[14\].yc/lin[0] blk.column\[4\].row\[14\].yc/lin[1]
+ blk.column\[5\].row\[14\].yc/uempty blk.column\[5\].row\[14\].yc/uin[0] blk.column\[5\].row\[14\].yc/uin[1]
+ blk.column\[5\].row\[13\].yc/din[0] blk.column\[5\].row\[13\].yc/din[1] blk.column\[5\].row\[13\].yc/dempty
+ blk.column\[5\].row\[15\].yc/uempty VPWR VGND ycell
XFILLER_382_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_493_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_2465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_419_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_277_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_499_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_423_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_502_ VGND VGND VPWR VPWR _502_/HI _502_/LO sky130_fd_sc_hd__conb_1
XFILLER_497_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_480_2089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_444_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_433_ VGND VGND VPWR VPWR _433_/HI _433_/LO sky130_fd_sc_hd__conb_1
XFILLER_260_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_2075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_497_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_364_ _363_/Y _361_/X wbs_dat_i[30] _361_/X VGND VGND VPWR VPWR _782_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_536_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_295_ wb_rst_i VGND VGND VPWR VPWR _295_/Y sky130_fd_sc_hd__inv_2
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_375_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_534_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_375_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_355_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_256_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_491_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_520_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_387_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_467_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_506_3228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_485_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_428_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_283_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_506_1837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_397_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_440_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_338_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_536_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_530_2801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_1977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_448_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_515_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_407_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_509_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_3099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_2026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_416_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_524_1959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_2947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_400_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_342_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_498_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_279_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_539_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_337_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_409_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_352_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_502_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_216_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_940 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_2130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_394_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_466_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_267_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_486_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_10256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_361_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_482_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_366_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_308_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_218_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_3130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_501_3136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_407_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_2484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_458_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_505_1892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_416_ _412_/X wbs_dat_o[7] _807_/Q _410_/X VGND VGND VPWR VPWR _416_/X sky130_fd_sc_hd__o22a_4
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_394_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_1745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_2794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_537_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_375_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_347_ _347_/A VGND VGND VPWR VPWR _347_/Y sky130_fd_sc_hd__inv_2
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_493_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_466_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_315_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_3232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_512_2520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_469_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_303_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_335_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_465_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_1874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_250_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_486_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_271_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_3069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_472_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_326_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_406_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_402_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_2660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_421_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_2111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_476_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_292_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_319_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_413_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_530_2642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_533_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_462_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_245_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_487_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_247_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_262_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_246_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_481_2184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_285_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_227_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_420_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_502_2777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_537_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_3191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_396_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_535_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_357_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_372_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_407_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_273_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_238_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_292_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_234_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_314_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_3014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_502_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_372_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_297_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_340_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_9696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_300_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_278_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_388_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_384_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_529_1623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_439_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_542_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_10075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_293_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_464_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_452_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_507_2611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_3209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_454_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_280_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_425_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_507_1965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_527_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_245_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_450_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_340_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_501_2221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_321_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[11\].row\[5\].yc blk.column\[11\].row\[5\].yc/cbitin blk.column\[11\].row\[6\].yc/cbitin
+ blk.column\[11\].row\[5\].yc/confclk blk.column\[11\].row\[6\].yc/confclk blk.column\[11\].row\[5\].yc/dempty
+ blk.column\[11\].row\[5\].yc/din[0] blk.column\[11\].row\[5\].yc/din[1] blk.column\[11\].row\[6\].yc/uin[0]
+ blk.column\[11\].row\[6\].yc/uin[1] blk.column\[11\].row\[5\].yc/hempty blk.column\[10\].row\[5\].yc/lempty
+ blk.column\[11\].row\[5\].yc/lempty blk.column\[11\].row\[5\].yc/lin[0] blk.column\[11\].row\[5\].yc/lin[1]
+ blk.column\[12\].row\[5\].yc/rin[0] blk.column\[12\].row\[5\].yc/rin[1] blk.column\[10\].row\[5\].yc/hempty
+ blk.column\[11\].row\[5\].yc/reset blk.column\[11\].row\[6\].yc/reset blk.column\[11\].row\[5\].yc/rin[0]
+ blk.column\[11\].row\[5\].yc/rin[1] blk.column\[10\].row\[5\].yc/lin[0] blk.column\[10\].row\[5\].yc/lin[1]
+ blk.column\[11\].row\[5\].yc/uempty blk.column\[11\].row\[5\].yc/uin[0] blk.column\[11\].row\[5\].yc/uin[1]
+ blk.column\[11\].row\[4\].yc/din[0] blk.column\[11\].row\[4\].yc/din[1] blk.column\[11\].row\[4\].yc/dempty
+ blk.column\[11\].row\[6\].yc/uempty VPWR VGND ycell
XFILLER_538_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_221_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_340_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_395_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_375_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_471_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_291_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_331_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_282_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[2\].row\[6\].yc blk.column\[2\].row\[6\].yc/cbitin blk.column\[2\].row\[7\].yc/cbitin
+ blk.column\[2\].row\[6\].yc/confclk blk.column\[2\].row\[7\].yc/confclk blk.column\[2\].row\[6\].yc/dempty
+ blk.column\[2\].row\[6\].yc/din[0] blk.column\[2\].row\[6\].yc/din[1] blk.column\[2\].row\[7\].yc/uin[0]
+ blk.column\[2\].row\[7\].yc/uin[1] blk.column\[2\].row\[6\].yc/hempty blk.column\[1\].row\[6\].yc/lempty
+ blk.column\[2\].row\[6\].yc/lempty blk.column\[2\].row\[6\].yc/lin[0] blk.column\[2\].row\[6\].yc/lin[1]
+ blk.column\[3\].row\[6\].yc/rin[0] blk.column\[3\].row\[6\].yc/rin[1] blk.column\[1\].row\[6\].yc/hempty
+ blk.column\[2\].row\[6\].yc/reset blk.column\[2\].row\[7\].yc/reset blk.column\[2\].row\[6\].yc/rin[0]
+ blk.column\[2\].row\[6\].yc/rin[1] blk.column\[1\].row\[6\].yc/lin[0] blk.column\[1\].row\[6\].yc/lin[1]
+ blk.column\[2\].row\[6\].yc/uempty blk.column\[2\].row\[6\].yc/uin[0] blk.column\[2\].row\[6\].yc/uin[1]
+ blk.column\[2\].row\[5\].yc/din[0] blk.column\[2\].row\[5\].yc/din[1] blk.column\[2\].row\[5\].yc/dempty
+ blk.column\[2\].row\[7\].yc/uempty VPWR VGND ycell
XFILLER_332_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_477_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_328_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_362_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_269_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_215_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_229_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_2880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_2001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_244_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_506_2154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_478_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_2288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_398_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_358_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_401_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_1276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_296_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_381_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_2937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_317_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_2294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_2136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_489_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_279_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_530_2472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_496_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_448_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_322_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_213_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_294_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_467_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_268_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_526_2508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_750_ wb_clk_i _418_/X VGND VGND VPWR VPWR wbs_dat_o[6] sky130_fd_sc_hd__dfxtp_4
XPHY_7557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_483_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_229_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_2177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_436_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_363_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_681_ VGND VGND VPWR VPWR _681_/HI la_data_out[65] sky130_fd_sc_hd__conb_1
XFILLER_422_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_309_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_305_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_2276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_389_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_432_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_404_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_524_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_455_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_502_1862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_240_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_2925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_275_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_535_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_518_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_534_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_372_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_316_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_390_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_360_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_531_2258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_383_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_313_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_459_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_466_3134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_488_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_411_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_474_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_2807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[7\].row\[0\].yc la_data_in[103] blk.column\[7\].row\[1\].yc/cbitin la_data_in[112]
+ blk.column\[7\].row\[1\].yc/confclk blk.column\[7\].row\[0\].yc/dempty blk.column\[7\].row\[0\].yc/din[0]
+ blk.column\[7\].row\[0\].yc/din[1] blk.column\[7\].row\[1\].yc/uin[0] blk.column\[7\].row\[1\].yc/uin[1]
+ blk.column\[7\].row\[0\].yc/hempty blk.column\[6\].row\[0\].yc/lempty blk.column\[7\].row\[0\].yc/lempty
+ blk.column\[7\].row\[0\].yc/lin[0] blk.column\[7\].row\[0\].yc/lin[1] blk.column\[8\].row\[0\].yc/rin[0]
+ blk.column\[8\].row\[0\].yc/rin[1] blk.column\[6\].row\[0\].yc/hempty la_data_in[113]
+ blk.column\[7\].row\[1\].yc/reset blk.column\[7\].row\[0\].yc/rin[0] blk.column\[7\].row\[0\].yc/rin[1]
+ blk.column\[6\].row\[0\].yc/lin[0] blk.column\[6\].row\[0\].yc/lin[1] _579_/LO la_data_in[78]
+ la_data_in[79] la_data_out[14] la_data_out[15] blk.column\[7\].row\[0\].yc/vempty
+ blk.column\[7\].row\[1\].yc/uempty VPWR VGND ycell
XFILLER_78_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_3221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_226_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_3197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_482_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_323_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_2575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_2630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_1675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_501_2062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_1574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_395_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_277_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_379_2961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_2125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_363_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_536_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_3179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_275_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_217_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_330_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_507_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_410_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_236_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_304_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_1788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_2191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_276_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_2691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_484_2533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_367_3054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_257_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_2987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_3017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_408_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_2563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_484_1898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_521_2416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_228_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_414_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_282_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_224_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_2916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_386_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_519_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_243_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_1196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_323_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_3183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_3036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_339_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_393_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_393_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_354_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_434_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_274_3170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_3112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_473_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_3066 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_270_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_2672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xblk.column\[0\].row\[15\].yc blk.column\[0\].row\[15\].yc/cbitin la_data_out[32]
+ blk.column\[0\].row\[15\].yc/confclk blk.column\[0\].row\[15\].yc/confclko _434_/HI
+ _489_/LO _490_/LO blk.column\[0\].row\[15\].yc/dout[0] blk.column\[0\].row\[15\].yc/dout[1]
+ blk.column\[0\].row\[15\].yc/hempty blk.column\[0\].row\[15\].yc/hempty2 blk.column\[0\].row\[15\].yc/lempty
+ blk.column\[0\].row\[15\].yc/lin[0] blk.column\[0\].row\[15\].yc/lin[1] blk.column\[1\].row\[15\].yc/rin[0]
+ blk.column\[1\].row\[15\].yc/rin[1] _435_/HI blk.column\[0\].row\[15\].yc/reset
+ blk.column\[0\].row\[15\].yc/reseto _491_/LO _492_/LO blk.column\[0\].row\[15\].yc/rout[0]
+ blk.column\[0\].row\[15\].yc/rout[1] blk.column\[0\].row\[15\].yc/uempty blk.column\[0\].row\[15\].yc/uin[0]
+ blk.column\[0\].row\[15\].yc/uin[1] blk.column\[0\].row\[14\].yc/din[0] blk.column\[0\].row\[14\].yc/din[1]
+ blk.column\[0\].row\[14\].yc/dempty blk.column\[0\].row\[15\].yc/vempty2 VPWR VGND
+ ycell
XFILLER_342_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_235_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_310_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_1721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_311_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_489_2477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_511_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_2319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_456_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_330_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_802_ wb_clk_i _311_/X VGND VGND VPWR VPWR _802_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_433_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_8099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_385_3176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_474_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_733_ VGND VGND VPWR VPWR _733_/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XPHY_7387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_492_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_461_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_2087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_2862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_426_3195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_664_ VGND VGND VPWR VPWR _664_/HI la_data_out[48] sky130_fd_sc_hd__conb_1
XPHY_6697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_480_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_281_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_263_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_302_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_422_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xblk.column\[14\].row\[11\].yc blk.column\[14\].row\[11\].yc/cbitin blk.column\[14\].row\[12\].yc/cbitin
+ blk.column\[14\].row\[11\].yc/confclk blk.column\[14\].row\[12\].yc/confclk blk.column\[14\].row\[11\].yc/dempty
+ blk.column\[14\].row\[11\].yc/din[0] blk.column\[14\].row\[11\].yc/din[1] blk.column\[14\].row\[12\].yc/uin[0]
+ blk.column\[14\].row\[12\].yc/uin[1] blk.column\[14\].row\[11\].yc/hempty blk.column\[13\].row\[11\].yc/lempty
+ blk.column\[14\].row\[11\].yc/lempty blk.column\[14\].row\[11\].yc/lin[0] blk.column\[14\].row\[11\].yc/lin[1]
+ blk.column\[15\].row\[11\].yc/rin[0] blk.column\[15\].row\[11\].yc/rin[1] blk.column\[13\].row\[11\].yc/hempty
+ blk.column\[14\].row\[11\].yc/reset blk.column\[14\].row\[12\].yc/reset blk.column\[14\].row\[11\].yc/rin[0]
+ blk.column\[14\].row\[11\].yc/rin[1] blk.column\[13\].row\[11\].yc/lin[0] blk.column\[13\].row\[11\].yc/lin[1]
+ blk.column\[14\].row\[11\].yc/uempty blk.column\[14\].row\[11\].yc/uin[0] blk.column\[14\].row\[11\].yc/uin[1]
+ blk.column\[14\].row\[10\].yc/din[0] blk.column\[14\].row\[10\].yc/din[1] blk.column\[14\].row\[10\].yc/dempty
+ blk.column\[14\].row\[12\].yc/uempty VPWR VGND ycell
XFILLER_17_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_595_ VGND VGND VPWR VPWR _595_/HI io_oeb[7] sky130_fd_sc_hd__conb_1
XFILLER_524_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_242_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_378_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_231_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_502_3094 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_377_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_259_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_318_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_345_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_2594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_392_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_1733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_2447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_515_2721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_494_1471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_518_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2069 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_433_3188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_474_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_2099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_1928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_530_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_258_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_485_2831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_509_2514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_1264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_343_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_239_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_286_3085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_254_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_2648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_2587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_405_3213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_2703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_415_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_529_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_509_1879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_212_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_507_2282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_525_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_430_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_542_2195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_499_2050 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_368_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_301_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_307_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_288_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_411_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_223_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_503_1489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_2922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_1508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_492_2813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_538_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_495_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_457_2966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_525_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_451_3200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_418_2939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_219_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_336_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_537_2990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_293_3078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_533_2843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_540_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_3091 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_498_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_2581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_391_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_324_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_351_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_541_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_514_2264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_510_2106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_384_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_289_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_237_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_334_3097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_11309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_522_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_369_3127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_486_2606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_438_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_253_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_230_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_470_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_253_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_2020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_493_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_265_3103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_527_2636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_2374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_5215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_508_2057 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_461_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_306_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_403_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_540_2825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_3073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_360_2913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_260_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_521_1501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_401_2910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_380_ _419_/A VGND VGND VPWR VPWR _391_/A sky130_fd_sc_hd__buf_2
XPHY_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_497_2746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_3109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_495_3160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_359_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_491_3002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_456_3122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_374_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_2892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_517_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_327_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_3030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_534_2618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_417_3139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_222_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_3021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_1611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_2197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_519_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_505_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_491_2367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_2963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_516_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_488_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_294_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_1630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_532_2386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_469_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_219_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_512_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_513_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_497_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_2014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_484_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_350_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_489_1562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_295_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_485_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_485_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_380_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_289_2958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_463_3115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_289_2969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_2935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_283_3225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_2716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_3012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_369_2993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[12\].row\[7\].yc blk.column\[12\].row\[7\].yc/cbitin blk.column\[12\].row\[8\].yc/cbitin
+ blk.column\[12\].row\[7\].yc/confclk blk.column\[12\].row\[8\].yc/confclk blk.column\[12\].row\[7\].yc/dempty
+ blk.column\[12\].row\[7\].yc/din[0] blk.column\[12\].row\[7\].yc/din[1] blk.column\[12\].row\[8\].yc/uin[0]
+ blk.column\[12\].row\[8\].yc/uin[1] blk.column\[12\].row\[7\].yc/hempty blk.column\[11\].row\[7\].yc/lempty
+ blk.column\[12\].row\[7\].yc/lempty blk.column\[12\].row\[7\].yc/lin[0] blk.column\[12\].row\[7\].yc/lin[1]
+ blk.column\[13\].row\[7\].yc/rin[0] blk.column\[13\].row\[7\].yc/rin[1] blk.column\[11\].row\[7\].yc/hempty
+ blk.column\[12\].row\[7\].yc/reset blk.column\[12\].row\[8\].yc/reset blk.column\[12\].row\[7\].yc/rin[0]
+ blk.column\[12\].row\[7\].yc/rin[1] blk.column\[11\].row\[7\].yc/lin[0] blk.column\[11\].row\[7\].yc/lin[1]
+ blk.column\[12\].row\[7\].yc/uempty blk.column\[12\].row\[7\].yc/uin[0] blk.column\[12\].row\[7\].yc/uin[1]
+ blk.column\[12\].row\[6\].yc/din[0] blk.column\[12\].row\[6\].yc/din[1] blk.column\[12\].row\[6\].yc/dempty
+ blk.column\[12\].row\[8\].yc/uempty VPWR VGND ycell
XFILLER_236_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_6450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_7195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_716_ VGND VGND VPWR VPWR _716_/HI la_data_out[100] sky130_fd_sc_hd__conb_1
XFILLER_185_2934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_526_2179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_2411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_460_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_6494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_313_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_3167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_483_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_647_ VGND VGND VPWR VPWR _647_/HI io_out[21] sky130_fd_sc_hd__conb_1
XFILLER_412_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_578_ VGND VGND VPWR VPWR _578_/HI _578_/LO sky130_fd_sc_hd__conb_1
XFILLER_226_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_524_1191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_1776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_520_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_500_1618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_2667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_220_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_1806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_539_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_2289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_496_1544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_357_3042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xblk.column\[3\].row\[8\].yc blk.column\[3\].row\[8\].yc/cbitin blk.column\[3\].row\[9\].yc/cbitin
+ blk.column\[3\].row\[8\].yc/confclk blk.column\[3\].row\[9\].yc/confclk blk.column\[3\].row\[8\].yc/dempty
+ blk.column\[3\].row\[8\].yc/din[0] blk.column\[3\].row\[8\].yc/din[1] blk.column\[3\].row\[9\].yc/uin[0]
+ blk.column\[3\].row\[9\].yc/uin[1] blk.column\[3\].row\[8\].yc/hempty blk.column\[2\].row\[8\].yc/lempty
+ blk.column\[3\].row\[8\].yc/lempty blk.column\[3\].row\[8\].yc/lin[0] blk.column\[3\].row\[8\].yc/lin[1]
+ blk.column\[4\].row\[8\].yc/rin[0] blk.column\[4\].row\[8\].yc/rin[1] blk.column\[2\].row\[8\].yc/hempty
+ blk.column\[3\].row\[8\].yc/reset blk.column\[3\].row\[9\].yc/reset blk.column\[3\].row\[8\].yc/rin[0]
+ blk.column\[3\].row\[8\].yc/rin[1] blk.column\[2\].row\[8\].yc/lin[0] blk.column\[2\].row\[8\].yc/lin[1]
+ blk.column\[3\].row\[8\].yc/uempty blk.column\[3\].row\[8\].yc/uin[0] blk.column\[3\].row\[8\].yc/uin[1]
+ blk.column\[3\].row\[7\].yc/din[0] blk.column\[3\].row\[7\].yc/din[1] blk.column\[3\].row\[7\].yc/dempty
+ blk.column\[3\].row\[9\].yc/uempty VPWR VGND ycell
XFILLER_507_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_3207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_3152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_376_2975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_318_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_508_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_535_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_522_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_370_3231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_537_1585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_533_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_373_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_333_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_306_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_511_2404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_523_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_490_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_272_2951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_214_3024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_487_2904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_504_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_468_3048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_233_2946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_2868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_531_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_288_3158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_290_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_3124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_528_2923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_313_2981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3063 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_475_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

