magic
tech sky130A
magscale 1 2
timestamp 1608218641
<< locali >>
rect 9505 6647 9539 6817
<< viali >>
rect 7665 12733 7699 12767
rect 7757 12597 7791 12631
rect 3433 11713 3467 11747
rect 3709 11645 3743 11679
rect 4813 11509 4847 11543
rect 7573 10761 7607 10795
rect 6837 10625 6871 10659
rect 5917 10557 5951 10591
rect 6377 10557 6411 10591
rect 6929 10557 6963 10591
rect 7481 10557 7515 10591
rect 7389 10489 7423 10523
rect 6009 10421 6043 10455
rect 6469 10421 6503 10455
rect 5733 10217 5767 10251
rect 5365 10081 5399 10115
rect 5641 10081 5675 10115
rect 5917 10081 5951 10115
rect 6607 10081 6641 10115
rect 6745 10081 6779 10115
rect 7021 10081 7055 10115
rect 7849 10081 7883 10115
rect 8125 10081 8159 10115
rect 6469 10013 6503 10047
rect 7389 10013 7423 10047
rect 7665 10013 7699 10047
rect 8217 9945 8251 9979
rect 5457 9877 5491 9911
rect 7159 9877 7193 9911
rect 7297 9877 7331 9911
rect 7941 9877 7975 9911
rect 4978 9673 5012 9707
rect 5089 9605 5123 9639
rect 3433 9537 3467 9571
rect 3985 9537 4019 9571
rect 5181 9537 5215 9571
rect 6193 9537 6227 9571
rect 7389 9537 7423 9571
rect 1961 9469 1995 9503
rect 3525 9469 3559 9503
rect 4261 9469 4295 9503
rect 4629 9469 4663 9503
rect 4813 9469 4847 9503
rect 6469 9469 6503 9503
rect 6653 9469 6687 9503
rect 7665 9469 7699 9503
rect 7849 9469 7883 9503
rect 8033 9469 8067 9503
rect 8401 9469 8435 9503
rect 8769 9469 8803 9503
rect 5641 9401 5675 9435
rect 6837 9401 6871 9435
rect 2053 9333 2087 9367
rect 5457 9333 5491 9367
rect 8033 9333 8067 9367
rect 8861 9333 8895 9367
rect 7573 9129 7607 9163
rect 3157 8993 3191 9027
rect 4077 8993 4111 9027
rect 5457 8993 5491 9027
rect 5733 8993 5767 9027
rect 6285 8993 6319 9027
rect 6469 8993 6503 9027
rect 6561 8993 6595 9027
rect 7941 8993 7975 9027
rect 8309 8993 8343 9027
rect 8585 8993 8619 9027
rect 9229 8993 9263 9027
rect 4261 8925 4295 8959
rect 4629 8925 4663 8959
rect 5181 8925 5215 8959
rect 5641 8925 5675 8959
rect 6929 8925 6963 8959
rect 7113 8925 7147 8959
rect 7849 8925 7883 8959
rect 8217 8925 8251 8959
rect 3249 8789 3283 8823
rect 8677 8789 8711 8823
rect 3157 8585 3191 8619
rect 10333 8585 10367 8619
rect 8677 8517 8711 8551
rect 9827 8517 9861 8551
rect 9965 8517 9999 8551
rect 4629 8449 4663 8483
rect 8217 8449 8251 8483
rect 8861 8449 8895 8483
rect 10057 8449 10091 8483
rect 3065 8381 3099 8415
rect 3801 8381 3835 8415
rect 3985 8381 4019 8415
rect 4353 8381 4387 8415
rect 6285 8381 6319 8415
rect 6653 8381 6687 8415
rect 7297 8381 7331 8415
rect 7481 8381 7515 8415
rect 7757 8381 7791 8415
rect 7941 8381 7975 8415
rect 9045 8381 9079 8415
rect 9413 8381 9447 8415
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 10517 8381 10551 8415
rect 2881 8313 2915 8347
rect 4261 8313 4295 8347
rect 6101 8313 6135 8347
rect 6837 8313 6871 8347
rect 10609 8313 10643 8347
rect 5733 8245 5767 8279
rect 2697 8041 2731 8075
rect 8585 8041 8619 8075
rect 9137 8041 9171 8075
rect 9781 8041 9815 8075
rect 10701 8041 10735 8075
rect 2421 7973 2455 8007
rect 4077 7973 4111 8007
rect 4629 7973 4663 8007
rect 8861 7973 8895 8007
rect 11253 7973 11287 8007
rect 2329 7905 2363 7939
rect 3249 7905 3283 7939
rect 3617 7905 3651 7939
rect 4261 7905 4295 7939
rect 5273 7905 5307 7939
rect 5549 7905 5583 7939
rect 6285 7905 6319 7939
rect 6469 7905 6503 7939
rect 6745 7905 6779 7939
rect 7297 7905 7331 7939
rect 7573 7905 7607 7939
rect 7665 7905 7699 7939
rect 8033 7905 8067 7939
rect 8125 7905 8159 7939
rect 9045 7905 9079 7939
rect 9689 7905 9723 7939
rect 10149 7905 10183 7939
rect 10517 7905 10551 7939
rect 10885 7905 10919 7939
rect 11161 7905 11195 7939
rect 3341 7837 3375 7871
rect 3525 7837 3559 7871
rect 4721 7837 4755 7871
rect 5733 7837 5767 7871
rect 5825 7837 5859 7871
rect 6929 7837 6963 7871
rect 10977 7701 11011 7735
rect 2053 7429 2087 7463
rect 1777 7361 1811 7395
rect 3157 7361 3191 7395
rect 3709 7361 3743 7395
rect 4353 7361 4387 7395
rect 6561 7361 6595 7395
rect 8217 7361 8251 7395
rect 8861 7361 8895 7395
rect 9413 7361 9447 7395
rect 10103 7361 10137 7395
rect 1685 7293 1719 7327
rect 1961 7293 1995 7327
rect 2513 7293 2547 7327
rect 2697 7293 2731 7327
rect 3053 7293 3087 7327
rect 3341 7293 3375 7327
rect 4537 7293 4571 7327
rect 4905 7293 4939 7327
rect 5089 7293 5123 7327
rect 5181 7293 5215 7327
rect 5641 7293 5675 7327
rect 5917 7293 5951 7327
rect 6101 7293 6135 7327
rect 6469 7293 6503 7327
rect 7297 7293 7331 7327
rect 7481 7293 7515 7327
rect 7849 7293 7883 7327
rect 7941 7293 7975 7327
rect 8769 7293 8803 7327
rect 9137 7293 9171 7327
rect 9321 7293 9355 7327
rect 9965 7293 9999 7327
rect 10241 7293 10275 7327
rect 10517 7293 10551 7327
rect 10609 7293 10643 7327
rect 10793 7293 10827 7327
rect 11345 7293 11379 7327
rect 2329 7157 2363 7191
rect 4169 7157 4203 7191
rect 7113 7157 7147 7191
rect 10977 7157 11011 7191
rect 11437 7157 11471 7191
rect 2513 6817 2547 6851
rect 2697 6817 2731 6851
rect 3157 6817 3191 6851
rect 3525 6817 3559 6851
rect 3893 6817 3927 6851
rect 6561 6817 6595 6851
rect 6653 6817 6687 6851
rect 6929 6817 6963 6851
rect 8033 6817 8067 6851
rect 8217 6817 8251 6851
rect 8493 6817 8527 6851
rect 9137 6817 9171 6851
rect 9505 6817 9539 6851
rect 9689 6817 9723 6851
rect 10517 6817 10551 6851
rect 10701 6817 10735 6851
rect 4261 6749 4295 6783
rect 4537 6749 4571 6783
rect 5641 6749 5675 6783
rect 6009 6749 6043 6783
rect 7113 6749 7147 6783
rect 7389 6749 7423 6783
rect 7573 6749 7607 6783
rect 8677 6749 8711 6783
rect 8953 6749 8987 6783
rect 10057 6749 10091 6783
rect 10149 6681 10183 6715
rect 2789 6613 2823 6647
rect 9321 6613 9355 6647
rect 9505 6613 9539 6647
rect 9827 6613 9861 6647
rect 9965 6613 9999 6647
rect 10793 6613 10827 6647
rect 3874 6409 3908 6443
rect 4169 6409 4203 6443
rect 3985 6341 4019 6375
rect 4077 6273 4111 6307
rect 5641 6273 5675 6307
rect 7941 6273 7975 6307
rect 8217 6273 8251 6307
rect 8953 6273 8987 6307
rect 3433 6205 3467 6239
rect 5089 6205 5123 6239
rect 5365 6205 5399 6239
rect 5549 6205 5583 6239
rect 6193 6205 6227 6239
rect 6469 6205 6503 6239
rect 6653 6205 6687 6239
rect 7297 6205 7331 6239
rect 7573 6205 7607 6239
rect 7757 6205 7791 6239
rect 8401 6205 8435 6239
rect 9137 6205 9171 6239
rect 9597 6205 9631 6239
rect 9873 6205 9907 6239
rect 10333 6205 10367 6239
rect 3709 6137 3743 6171
rect 4537 6137 4571 6171
rect 6837 6137 6871 6171
rect 8769 6137 8803 6171
rect 3525 6069 3559 6103
rect 7573 5865 7607 5899
rect 4261 5729 4295 5763
rect 4445 5729 4479 5763
rect 5089 5729 5123 5763
rect 5917 5729 5951 5763
rect 6837 5729 6871 5763
rect 7205 5729 7239 5763
rect 7757 5729 7791 5763
rect 8033 5729 8067 5763
rect 8953 5729 8987 5763
rect 9321 5729 9355 5763
rect 9689 5729 9723 5763
rect 5641 5661 5675 5695
rect 6101 5661 6135 5695
rect 6653 5661 6687 5695
rect 7113 5661 7147 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 9781 5661 9815 5695
rect 6469 5593 6503 5627
rect 4537 5525 4571 5559
rect 8585 5525 8619 5559
rect 7757 5253 7791 5287
rect 6653 5185 6687 5219
rect 8401 5185 8435 5219
rect 4997 5117 5031 5151
rect 5273 5117 5307 5151
rect 5733 5117 5767 5151
rect 6009 5117 6043 5151
rect 6286 5117 6320 5151
rect 7113 5117 7147 5151
rect 7389 5117 7423 5151
rect 7665 5117 7699 5151
rect 7941 5117 7975 5151
rect 6101 5049 6135 5083
rect 4813 4981 4847 5015
rect 6929 4981 6963 5015
rect 5733 4777 5767 4811
rect 10885 4777 10919 4811
rect 5365 4641 5399 4675
rect 5641 4641 5675 4675
rect 5917 4641 5951 4675
rect 6009 4641 6043 4675
rect 6193 4641 6227 4675
rect 6469 4641 6503 4675
rect 7021 4641 7055 4675
rect 7113 4641 7147 4675
rect 7297 4641 7331 4675
rect 8401 4641 8435 4675
rect 8585 4641 8619 4675
rect 8953 4641 8987 4675
rect 9045 4641 9079 4675
rect 9137 4641 9171 4675
rect 9873 4641 9907 4675
rect 10333 4641 10367 4675
rect 10425 4641 10459 4675
rect 6653 4573 6687 4607
rect 7757 4573 7791 4607
rect 9781 4573 9815 4607
rect 6285 4505 6319 4539
rect 5457 4437 5491 4471
rect 6561 4233 6595 4267
rect 6929 4233 6963 4267
rect 8493 4233 8527 4267
rect 8953 4097 8987 4131
rect 9137 4097 9171 4131
rect 6469 4029 6503 4063
rect 6837 4029 6871 4063
rect 8861 4029 8895 4063
rect 9229 4029 9263 4063
rect 1409 3553 1443 3587
rect 2421 3553 2455 3587
rect 1593 3349 1627 3383
rect 2605 3349 2639 3383
rect 7665 2941 7699 2975
rect 7849 2805 7883 2839
rect 7021 2465 7055 2499
rect 7113 2261 7147 2295
<< metal1 >>
rect 1104 13082 11960 13104
rect 1104 13030 2791 13082
rect 2843 13030 2855 13082
rect 2907 13030 2919 13082
rect 2971 13030 2983 13082
rect 3035 13030 6410 13082
rect 6462 13030 6474 13082
rect 6526 13030 6538 13082
rect 6590 13030 6602 13082
rect 6654 13030 10028 13082
rect 10080 13030 10092 13082
rect 10144 13030 10156 13082
rect 10208 13030 10220 13082
rect 10272 13030 11960 13082
rect 1104 13008 11960 13030
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 7834 12764 7840 12776
rect 7699 12736 7840 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7745 12631 7803 12637
rect 7745 12628 7757 12631
rect 6972 12600 7757 12628
rect 6972 12588 6978 12600
rect 7745 12597 7757 12600
rect 7791 12597 7803 12631
rect 7745 12591 7803 12597
rect 1104 12538 11960 12560
rect 1104 12486 4600 12538
rect 4652 12486 4664 12538
rect 4716 12486 4728 12538
rect 4780 12486 4792 12538
rect 4844 12486 8219 12538
rect 8271 12486 8283 12538
rect 8335 12486 8347 12538
rect 8399 12486 8411 12538
rect 8463 12486 11960 12538
rect 1104 12464 11960 12486
rect 1104 11994 11960 12016
rect 1104 11942 2791 11994
rect 2843 11942 2855 11994
rect 2907 11942 2919 11994
rect 2971 11942 2983 11994
rect 3035 11942 6410 11994
rect 6462 11942 6474 11994
rect 6526 11942 6538 11994
rect 6590 11942 6602 11994
rect 6654 11942 10028 11994
rect 10080 11942 10092 11994
rect 10144 11942 10156 11994
rect 10208 11942 10220 11994
rect 10272 11942 11960 11994
rect 1104 11920 11960 11942
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 3421 11747 3479 11753
rect 3421 11744 3433 11747
rect 2096 11716 3433 11744
rect 2096 11704 2102 11716
rect 3421 11713 3433 11716
rect 3467 11744 3479 11747
rect 4338 11744 4344 11756
rect 3467 11716 4344 11744
rect 3467 11713 3479 11716
rect 3421 11707 3479 11713
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 4982 11704 4988 11756
rect 5040 11744 5046 11756
rect 7098 11744 7104 11756
rect 5040 11716 7104 11744
rect 5040 11704 5046 11716
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 3510 11636 3516 11688
rect 3568 11676 3574 11688
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 3568 11648 3709 11676
rect 3568 11636 3574 11648
rect 3697 11645 3709 11648
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4212 11512 4813 11540
rect 4212 11500 4218 11512
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 4801 11503 4859 11509
rect 1104 11450 11960 11472
rect 1104 11398 4600 11450
rect 4652 11398 4664 11450
rect 4716 11398 4728 11450
rect 4780 11398 4792 11450
rect 4844 11398 8219 11450
rect 8271 11398 8283 11450
rect 8335 11398 8347 11450
rect 8399 11398 8411 11450
rect 8463 11398 11960 11450
rect 1104 11376 11960 11398
rect 658 11024 664 11076
rect 716 11064 722 11076
rect 5350 11064 5356 11076
rect 716 11036 5356 11064
rect 716 11024 722 11036
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 12250 11064 12256 11076
rect 10560 11036 12256 11064
rect 10560 11024 10566 11036
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 1104 10906 11960 10928
rect 1104 10854 2791 10906
rect 2843 10854 2855 10906
rect 2907 10854 2919 10906
rect 2971 10854 2983 10906
rect 3035 10854 6410 10906
rect 6462 10854 6474 10906
rect 6526 10854 6538 10906
rect 6590 10854 6602 10906
rect 6654 10854 10028 10906
rect 10080 10854 10092 10906
rect 10144 10854 10156 10906
rect 10208 10854 10220 10906
rect 10272 10854 11960 10906
rect 1104 10832 11960 10854
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 9306 10792 9312 10804
rect 7607 10764 9312 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 8662 10724 8668 10736
rect 5920 10696 8668 10724
rect 5920 10597 5948 10696
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6788 10628 6837 10656
rect 6788 10616 6794 10628
rect 6825 10625 6837 10628
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 5905 10591 5963 10597
rect 5905 10557 5917 10591
rect 5951 10557 5963 10591
rect 6362 10588 6368 10600
rect 6323 10560 6368 10588
rect 5905 10551 5963 10557
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 6914 10588 6920 10600
rect 6827 10560 6920 10588
rect 6914 10548 6920 10560
rect 6972 10588 6978 10600
rect 7190 10588 7196 10600
rect 6972 10560 7196 10588
rect 6972 10548 6978 10560
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7374 10520 7380 10532
rect 7335 10492 7380 10520
rect 7374 10480 7380 10492
rect 7432 10480 7438 10532
rect 5997 10455 6055 10461
rect 5997 10421 6009 10455
rect 6043 10452 6055 10455
rect 6178 10452 6184 10464
rect 6043 10424 6184 10452
rect 6043 10421 6055 10424
rect 5997 10415 6055 10421
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6270 10412 6276 10464
rect 6328 10452 6334 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 6328 10424 6469 10452
rect 6328 10412 6334 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 7484 10452 7512 10551
rect 6788 10424 7512 10452
rect 6788 10412 6794 10424
rect 1104 10362 11960 10384
rect 1104 10310 4600 10362
rect 4652 10310 4664 10362
rect 4716 10310 4728 10362
rect 4780 10310 4792 10362
rect 4844 10310 8219 10362
rect 8271 10310 8283 10362
rect 8335 10310 8347 10362
rect 8399 10310 8411 10362
rect 8463 10310 11960 10362
rect 1104 10288 11960 10310
rect 5721 10251 5779 10257
rect 5721 10217 5733 10251
rect 5767 10248 5779 10251
rect 8018 10248 8024 10260
rect 5767 10220 8024 10248
rect 5767 10217 5779 10220
rect 5721 10211 5779 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 7926 10180 7932 10192
rect 7340 10152 7932 10180
rect 7340 10140 7346 10152
rect 7926 10140 7932 10152
rect 7984 10180 7990 10192
rect 7984 10152 8156 10180
rect 7984 10140 7990 10152
rect 5350 10112 5356 10124
rect 5311 10084 5356 10112
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6362 10112 6368 10124
rect 5951 10084 6368 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 5166 10004 5172 10056
rect 5224 10044 5230 10056
rect 5644 10044 5672 10075
rect 6362 10072 6368 10084
rect 6420 10112 6426 10124
rect 6595 10115 6653 10121
rect 6595 10112 6607 10115
rect 6420 10084 6607 10112
rect 6420 10072 6426 10084
rect 6595 10081 6607 10084
rect 6641 10081 6653 10115
rect 6595 10075 6653 10081
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 6914 10112 6920 10124
rect 6779 10084 6920 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 7742 10112 7748 10124
rect 7055 10084 7748 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 8128 10121 8156 10152
rect 7837 10115 7895 10121
rect 7837 10081 7849 10115
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 5224 10016 5672 10044
rect 5224 10004 5230 10016
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6236 10016 6469 10044
rect 6236 10004 6242 10016
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 6880 10016 7389 10044
rect 6880 10004 6886 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7650 10044 7656 10056
rect 7611 10016 7656 10044
rect 7377 10007 7435 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 7852 10044 7880 10075
rect 8754 10044 8760 10056
rect 7852 10016 8760 10044
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 7006 9936 7012 9988
rect 7064 9976 7070 9988
rect 8205 9979 8263 9985
rect 8205 9976 8217 9979
rect 7064 9948 8217 9976
rect 7064 9936 7070 9948
rect 8205 9945 8217 9948
rect 8251 9945 8263 9979
rect 8205 9939 8263 9945
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9908 5503 9911
rect 5626 9908 5632 9920
rect 5491 9880 5632 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 7147 9911 7205 9917
rect 7147 9908 7159 9911
rect 6144 9880 7159 9908
rect 6144 9868 6150 9880
rect 7147 9877 7159 9880
rect 7193 9877 7205 9911
rect 7147 9871 7205 9877
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 7466 9908 7472 9920
rect 7331 9880 7472 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7929 9911 7987 9917
rect 7929 9908 7941 9911
rect 7616 9880 7941 9908
rect 7616 9868 7622 9880
rect 7929 9877 7941 9880
rect 7975 9877 7987 9911
rect 7929 9871 7987 9877
rect 1104 9818 11960 9840
rect 1104 9766 2791 9818
rect 2843 9766 2855 9818
rect 2907 9766 2919 9818
rect 2971 9766 2983 9818
rect 3035 9766 6410 9818
rect 6462 9766 6474 9818
rect 6526 9766 6538 9818
rect 6590 9766 6602 9818
rect 6654 9766 10028 9818
rect 10080 9766 10092 9818
rect 10144 9766 10156 9818
rect 10208 9766 10220 9818
rect 10272 9766 11960 9818
rect 1104 9744 11960 9766
rect 4966 9707 5024 9713
rect 4966 9704 4978 9707
rect 4908 9676 4978 9704
rect 3418 9568 3424 9580
rect 3379 9540 3424 9568
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9568 4031 9571
rect 4908 9568 4936 9676
rect 4966 9673 4978 9676
rect 5012 9704 5024 9707
rect 5012 9676 5212 9704
rect 5012 9673 5024 9676
rect 4966 9667 5024 9673
rect 5074 9636 5080 9648
rect 5035 9608 5080 9636
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5184 9636 5212 9676
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 7650 9704 7656 9716
rect 7432 9676 7656 9704
rect 7432 9664 7438 9676
rect 7650 9664 7656 9676
rect 7708 9664 7714 9716
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 7926 9704 7932 9716
rect 7800 9676 7932 9704
rect 7800 9664 7806 9676
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 5534 9636 5540 9648
rect 5184 9608 5540 9636
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 9674 9636 9680 9648
rect 7392 9608 9680 9636
rect 5166 9568 5172 9580
rect 4019 9540 4936 9568
rect 5127 9540 5172 9568
rect 4019 9537 4031 9540
rect 3973 9531 4031 9537
rect 5166 9528 5172 9540
rect 5224 9528 5230 9580
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 6178 9568 6184 9580
rect 5316 9540 6184 9568
rect 5316 9528 5322 9540
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 7392 9577 7420 9608
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 9858 9568 9864 9580
rect 8260 9540 9864 9568
rect 8260 9528 8266 9540
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 3292 9472 3525 9500
rect 3292 9460 3298 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 4246 9500 4252 9512
rect 4207 9472 4252 9500
rect 3513 9463 3571 9469
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9500 4675 9503
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4663 9472 4813 9500
rect 4663 9469 4675 9472
rect 4617 9463 4675 9469
rect 4801 9469 4813 9472
rect 4847 9500 4859 9503
rect 5442 9500 5448 9512
rect 4847 9472 5448 9500
rect 4847 9469 4859 9472
rect 4801 9463 4859 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6454 9500 6460 9512
rect 6415 9472 6460 9500
rect 6454 9460 6460 9472
rect 6512 9460 6518 9512
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 7282 9500 7288 9512
rect 6687 9472 7288 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 5629 9435 5687 9441
rect 5629 9401 5641 9435
rect 5675 9432 5687 9435
rect 6656 9432 6684 9463
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 7650 9500 7656 9512
rect 7611 9472 7656 9500
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 7837 9503 7895 9509
rect 7837 9469 7849 9503
rect 7883 9469 7895 9503
rect 8018 9500 8024 9512
rect 7979 9472 8024 9500
rect 7837 9463 7895 9469
rect 5675 9404 6684 9432
rect 6825 9435 6883 9441
rect 5675 9401 5687 9404
rect 5629 9395 5687 9401
rect 6825 9401 6837 9435
rect 6871 9432 6883 9435
rect 7852 9432 7880 9463
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 8168 9472 8401 9500
rect 8168 9460 8174 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9030 9500 9036 9512
rect 8803 9472 9036 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 9030 9460 9036 9472
rect 9088 9500 9094 9512
rect 10778 9500 10784 9512
rect 9088 9472 10784 9500
rect 9088 9460 9094 9472
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 7926 9432 7932 9444
rect 6871 9404 7932 9432
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 3602 9364 3608 9376
rect 2087 9336 3608 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 3694 9324 3700 9376
rect 3752 9364 3758 9376
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 3752 9336 5457 9364
rect 3752 9324 3758 9336
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 8021 9367 8079 9373
rect 8021 9364 8033 9367
rect 6972 9336 8033 9364
rect 6972 9324 6978 9336
rect 8021 9333 8033 9336
rect 8067 9333 8079 9367
rect 8846 9364 8852 9376
rect 8807 9336 8852 9364
rect 8021 9327 8079 9333
rect 8846 9324 8852 9336
rect 8904 9324 8910 9376
rect 1104 9274 11960 9296
rect 1104 9222 4600 9274
rect 4652 9222 4664 9274
rect 4716 9222 4728 9274
rect 4780 9222 4792 9274
rect 4844 9222 8219 9274
rect 8271 9222 8283 9274
rect 8335 9222 8347 9274
rect 8399 9222 8411 9274
rect 8463 9222 11960 9274
rect 1104 9200 11960 9222
rect 7561 9163 7619 9169
rect 7561 9129 7573 9163
rect 7607 9160 7619 9163
rect 9582 9160 9588 9172
rect 7607 9132 9588 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 9582 9120 9588 9132
rect 9640 9160 9646 9172
rect 10410 9160 10416 9172
rect 9640 9132 10416 9160
rect 9640 9120 9646 9132
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 5626 9052 5632 9104
rect 5684 9092 5690 9104
rect 5684 9064 6592 9092
rect 5684 9052 5690 9064
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3510 9024 3516 9036
rect 3191 8996 3516 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4154 9024 4160 9036
rect 4111 8996 4160 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 5442 9024 5448 9036
rect 5403 8996 5448 9024
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5718 9024 5724 9036
rect 5679 8996 5724 9024
rect 5718 8984 5724 8996
rect 5776 8984 5782 9036
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 8993 6331 9027
rect 6454 9024 6460 9036
rect 6415 8996 6460 9024
rect 6273 8987 6331 8993
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4617 8959 4675 8965
rect 4617 8925 4629 8959
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 4264 8888 4292 8919
rect 4120 8860 4292 8888
rect 4632 8888 4660 8919
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5626 8956 5632 8968
rect 5587 8928 5632 8956
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 6288 8956 6316 8987
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 6564 9033 6592 9064
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 7190 9092 7196 9104
rect 6972 9064 7196 9092
rect 6972 9052 6978 9064
rect 7190 9052 7196 9064
rect 7248 9052 7254 9104
rect 7852 9064 8064 9092
rect 6549 9027 6607 9033
rect 6549 8993 6561 9027
rect 6595 8993 6607 9027
rect 7558 9024 7564 9036
rect 6549 8987 6607 8993
rect 6656 8996 7564 9024
rect 6656 8956 6684 8996
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 7852 9024 7880 9064
rect 7668 8996 7880 9024
rect 7929 9027 7987 9033
rect 6914 8956 6920 8968
rect 6288 8928 6684 8956
rect 6875 8928 6920 8956
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7098 8956 7104 8968
rect 7059 8928 7104 8956
rect 7098 8916 7104 8928
rect 7156 8916 7162 8968
rect 7190 8916 7196 8968
rect 7248 8956 7254 8968
rect 7668 8956 7696 8996
rect 7929 8993 7941 9027
rect 7975 8993 7987 9027
rect 7929 8987 7987 8993
rect 7834 8956 7840 8968
rect 7248 8928 7696 8956
rect 7795 8928 7840 8956
rect 7248 8916 7254 8928
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 5644 8888 5672 8916
rect 4632 8860 5672 8888
rect 7944 8888 7972 8987
rect 8036 8956 8064 9064
rect 8110 9052 8116 9104
rect 8168 9092 8174 9104
rect 8168 9064 8616 9092
rect 8168 9052 8174 9064
rect 8588 9033 8616 9064
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 8573 9027 8631 9033
rect 8573 8993 8585 9027
rect 8619 8993 8631 9027
rect 8573 8987 8631 8993
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 8036 8928 8217 8956
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8312 8956 8340 8987
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 9180 8996 9229 9024
rect 9180 8984 9186 8996
rect 9217 8993 9229 8996
rect 9263 9024 9275 9027
rect 9766 9024 9772 9036
rect 9263 8996 9772 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 8938 8956 8944 8968
rect 8312 8928 8944 8956
rect 8205 8919 8263 8925
rect 8938 8916 8944 8928
rect 8996 8916 9002 8968
rect 8570 8888 8576 8900
rect 7944 8860 8576 8888
rect 4120 8848 4126 8860
rect 3234 8820 3240 8832
rect 3195 8792 3240 8820
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4632 8820 4660 8860
rect 8570 8848 8576 8860
rect 8628 8848 8634 8900
rect 8754 8848 8760 8900
rect 8812 8888 8818 8900
rect 10318 8888 10324 8900
rect 8812 8860 10324 8888
rect 8812 8848 8818 8860
rect 10318 8848 10324 8860
rect 10376 8848 10382 8900
rect 4028 8792 4660 8820
rect 4028 8780 4034 8792
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 7190 8820 7196 8832
rect 5592 8792 7196 8820
rect 5592 8780 5598 8792
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 8665 8823 8723 8829
rect 8665 8820 8677 8823
rect 7340 8792 8677 8820
rect 7340 8780 7346 8792
rect 8665 8789 8677 8792
rect 8711 8789 8723 8823
rect 8665 8783 8723 8789
rect 1104 8730 11960 8752
rect 1104 8678 2791 8730
rect 2843 8678 2855 8730
rect 2907 8678 2919 8730
rect 2971 8678 2983 8730
rect 3035 8678 6410 8730
rect 6462 8678 6474 8730
rect 6526 8678 6538 8730
rect 6590 8678 6602 8730
rect 6654 8678 10028 8730
rect 10080 8678 10092 8730
rect 10144 8678 10156 8730
rect 10208 8678 10220 8730
rect 10272 8678 11960 8730
rect 1104 8656 11960 8678
rect 3145 8619 3203 8625
rect 3145 8585 3157 8619
rect 3191 8616 3203 8619
rect 3786 8616 3792 8628
rect 3191 8588 3792 8616
rect 3191 8585 3203 8588
rect 3145 8579 3203 8585
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 8938 8616 8944 8628
rect 7248 8588 8944 8616
rect 7248 8576 7254 8588
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 10318 8616 10324 8628
rect 9088 8588 9536 8616
rect 10279 8588 10324 8616
rect 9088 8576 9094 8588
rect 5442 8508 5448 8560
rect 5500 8548 5506 8560
rect 8665 8551 8723 8557
rect 5500 8520 8248 8548
rect 5500 8508 5506 8520
rect 4154 8480 4160 8492
rect 3068 8452 4160 8480
rect 3068 8421 3096 8452
rect 4154 8440 4160 8452
rect 4212 8480 4218 8492
rect 4617 8483 4675 8489
rect 4617 8480 4629 8483
rect 4212 8452 4629 8480
rect 4212 8440 4218 8452
rect 4617 8449 4629 8452
rect 4663 8449 4675 8483
rect 4617 8443 4675 8449
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 8220 8489 8248 8520
rect 8665 8517 8677 8551
rect 8711 8548 8723 8551
rect 9122 8548 9128 8560
rect 8711 8520 9128 8548
rect 8711 8517 8723 8520
rect 8665 8511 8723 8517
rect 9122 8508 9128 8520
rect 9180 8508 9186 8560
rect 9508 8548 9536 8588
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 9815 8551 9873 8557
rect 9815 8548 9827 8551
rect 9508 8520 9827 8548
rect 9815 8517 9827 8520
rect 9861 8517 9873 8551
rect 9950 8548 9956 8560
rect 9911 8520 9956 8548
rect 9815 8511 9873 8517
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 8205 8483 8263 8489
rect 5684 8452 7512 8480
rect 5684 8440 5690 8452
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 3970 8412 3976 8424
rect 3931 8384 3976 8412
rect 3789 8375 3847 8381
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 3418 8344 3424 8356
rect 2915 8316 3424 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 3418 8304 3424 8316
rect 3476 8304 3482 8356
rect 3804 8344 3832 8375
rect 3970 8372 3976 8384
rect 4028 8372 4034 8424
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8412 4399 8415
rect 4430 8412 4436 8424
rect 4387 8384 4436 8412
rect 4387 8381 4399 8384
rect 4341 8375 4399 8381
rect 4430 8372 4436 8384
rect 4488 8372 4494 8424
rect 5810 8372 5816 8424
rect 5868 8412 5874 8424
rect 6273 8415 6331 8421
rect 6273 8412 6285 8415
rect 5868 8384 6285 8412
rect 5868 8372 5874 8384
rect 6273 8381 6285 8384
rect 6319 8381 6331 8415
rect 6273 8375 6331 8381
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7098 8412 7104 8424
rect 6687 8384 7104 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7484 8421 7512 8452
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8846 8480 8852 8492
rect 8807 8452 8852 8480
rect 8205 8443 8263 8449
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 8956 8452 10057 8480
rect 7285 8415 7343 8421
rect 7285 8412 7297 8415
rect 7248 8384 7297 8412
rect 7248 8372 7254 8384
rect 7285 8381 7297 8384
rect 7331 8381 7343 8415
rect 7285 8375 7343 8381
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8381 7527 8415
rect 7742 8412 7748 8424
rect 7703 8384 7748 8412
rect 7469 8375 7527 8381
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 7834 8372 7840 8424
rect 7892 8412 7898 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7892 8384 7941 8412
rect 7892 8372 7898 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 4154 8344 4160 8356
rect 3804 8316 4160 8344
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4249 8347 4307 8353
rect 4249 8313 4261 8347
rect 4295 8313 4307 8347
rect 4249 8307 4307 8313
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 6178 8344 6184 8356
rect 6135 8316 6184 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 4264 8276 4292 8307
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8313 6883 8347
rect 6825 8307 6883 8313
rect 4338 8276 4344 8288
rect 4264 8248 4344 8276
rect 4338 8236 4344 8248
rect 4396 8236 4402 8288
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 5721 8279 5779 8285
rect 5721 8276 5733 8279
rect 4948 8248 5733 8276
rect 4948 8236 4954 8248
rect 5721 8245 5733 8248
rect 5767 8245 5779 8279
rect 6840 8276 6868 8307
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 8956 8344 8984 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 9122 8412 9128 8424
rect 9079 8384 9128 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8381 9551 8415
rect 9493 8375 9551 8381
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10502 8412 10508 8424
rect 9723 8384 10508 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 6972 8316 8984 8344
rect 6972 8304 6978 8316
rect 7926 8276 7932 8288
rect 6840 8248 7932 8276
rect 5721 8239 5779 8245
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9416 8276 9444 8375
rect 9508 8344 9536 8375
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 9582 8344 9588 8356
rect 9495 8316 9588 8344
rect 9582 8304 9588 8316
rect 9640 8344 9646 8356
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 9640 8316 10609 8344
rect 9640 8304 9646 8316
rect 10597 8313 10609 8316
rect 10643 8313 10655 8347
rect 10597 8307 10655 8313
rect 8812 8248 9444 8276
rect 8812 8236 8818 8248
rect 9490 8236 9496 8288
rect 9548 8276 9554 8288
rect 9950 8276 9956 8288
rect 9548 8248 9956 8276
rect 9548 8236 9554 8248
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 1104 8186 11960 8208
rect 1104 8134 4600 8186
rect 4652 8134 4664 8186
rect 4716 8134 4728 8186
rect 4780 8134 4792 8186
rect 4844 8134 8219 8186
rect 8271 8134 8283 8186
rect 8335 8134 8347 8186
rect 8399 8134 8411 8186
rect 8463 8134 11960 8186
rect 1104 8112 11960 8134
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 4246 8072 4252 8084
rect 2731 8044 4252 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 5074 8072 5080 8084
rect 4540 8044 5080 8072
rect 2406 8004 2412 8016
rect 2367 7976 2412 8004
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 3694 8004 3700 8016
rect 2516 7976 3700 8004
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 2516 7936 2544 7976
rect 3694 7964 3700 7976
rect 3752 7964 3758 8016
rect 4065 8007 4123 8013
rect 4065 7973 4077 8007
rect 4111 8004 4123 8007
rect 4338 8004 4344 8016
rect 4111 7976 4344 8004
rect 4111 7973 4123 7976
rect 4065 7967 4123 7973
rect 4338 7964 4344 7976
rect 4396 8004 4402 8016
rect 4540 8004 4568 8044
rect 5074 8032 5080 8044
rect 5132 8072 5138 8084
rect 8570 8072 8576 8084
rect 5132 8044 8156 8072
rect 8531 8044 8576 8072
rect 5132 8032 5138 8044
rect 4396 7976 4568 8004
rect 4617 8007 4675 8013
rect 4396 7964 4402 7976
rect 4617 7973 4629 8007
rect 4663 8004 4675 8007
rect 4663 7976 6316 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 2363 7908 2544 7936
rect 3237 7939 3295 7945
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 3237 7905 3249 7939
rect 3283 7905 3295 7939
rect 3602 7936 3608 7948
rect 3563 7908 3608 7936
rect 3237 7899 3295 7905
rect 3252 7732 3280 7899
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 5258 7936 5264 7948
rect 4295 7908 5120 7936
rect 5219 7908 5264 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 3510 7868 3516 7880
rect 3384 7840 3429 7868
rect 3471 7840 3516 7868
rect 3384 7828 3390 7840
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4709 7871 4767 7877
rect 4709 7868 4721 7871
rect 4212 7840 4721 7868
rect 4212 7828 4218 7840
rect 4709 7837 4721 7840
rect 4755 7837 4767 7871
rect 5092 7868 5120 7908
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 5534 7936 5540 7948
rect 5495 7908 5540 7936
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 6288 7945 6316 7976
rect 6472 7976 8064 8004
rect 6273 7939 6331 7945
rect 5644 7908 5856 7936
rect 5166 7868 5172 7880
rect 5079 7840 5172 7868
rect 4709 7831 4767 7837
rect 4724 7800 4752 7831
rect 5166 7828 5172 7840
rect 5224 7868 5230 7880
rect 5644 7868 5672 7908
rect 5828 7877 5856 7908
rect 6273 7905 6285 7939
rect 6319 7905 6331 7939
rect 6273 7899 6331 7905
rect 6362 7896 6368 7948
rect 6420 7936 6426 7948
rect 6472 7945 6500 7976
rect 6457 7939 6515 7945
rect 6457 7936 6469 7939
rect 6420 7908 6469 7936
rect 6420 7896 6426 7908
rect 6457 7905 6469 7908
rect 6503 7905 6515 7939
rect 6457 7899 6515 7905
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7936 6791 7939
rect 7006 7936 7012 7948
rect 6779 7908 7012 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 7006 7896 7012 7908
rect 7064 7896 7070 7948
rect 7282 7936 7288 7948
rect 7243 7908 7288 7936
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7905 7619 7939
rect 7561 7899 7619 7905
rect 7653 7939 7711 7945
rect 7653 7905 7665 7939
rect 7699 7936 7711 7939
rect 7742 7936 7748 7948
rect 7699 7908 7748 7936
rect 7699 7905 7711 7908
rect 7653 7899 7711 7905
rect 5224 7840 5672 7868
rect 5721 7871 5779 7877
rect 5224 7828 5230 7840
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 5859 7840 6929 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 5736 7800 5764 7831
rect 7576 7800 7604 7899
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 8036 7945 8064 7976
rect 8128 7945 8156 8044
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 9125 8075 9183 8081
rect 9125 8072 9137 8075
rect 8720 8044 9137 8072
rect 8720 8032 8726 8044
rect 9125 8041 9137 8044
rect 9171 8041 9183 8075
rect 9125 8035 9183 8041
rect 9769 8075 9827 8081
rect 9769 8041 9781 8075
rect 9815 8072 9827 8075
rect 9858 8072 9864 8084
rect 9815 8044 9864 8072
rect 9815 8041 9827 8044
rect 9769 8035 9827 8041
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10686 8072 10692 8084
rect 10647 8044 10692 8072
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 8849 8007 8907 8013
rect 8849 8004 8861 8007
rect 8444 7976 8861 8004
rect 8444 7964 8450 7976
rect 8849 7973 8861 7976
rect 8895 7973 8907 8007
rect 8849 7967 8907 7973
rect 8938 7964 8944 8016
rect 8996 8004 9002 8016
rect 11241 8007 11299 8013
rect 11241 8004 11253 8007
rect 8996 7976 11253 8004
rect 8996 7964 9002 7976
rect 11241 7973 11253 7976
rect 11287 7973 11299 8007
rect 11241 7967 11299 7973
rect 8021 7939 8079 7945
rect 8021 7905 8033 7939
rect 8067 7905 8079 7939
rect 8021 7899 8079 7905
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 8202 7896 8208 7948
rect 8260 7936 8266 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8260 7908 9045 7936
rect 8260 7896 8266 7908
rect 9033 7905 9045 7908
rect 9079 7905 9091 7939
rect 9033 7899 9091 7905
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9692 7868 9720 7899
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10137 7939 10195 7945
rect 10137 7936 10149 7939
rect 9824 7908 10149 7936
rect 9824 7896 9830 7908
rect 10137 7905 10149 7908
rect 10183 7905 10195 7939
rect 10137 7899 10195 7905
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 10686 7936 10692 7948
rect 10551 7908 10692 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 10873 7939 10931 7945
rect 10873 7905 10885 7939
rect 10919 7905 10931 7939
rect 11146 7936 11152 7948
rect 11107 7908 11152 7936
rect 10873 7899 10931 7905
rect 8628 7840 9720 7868
rect 8628 7828 8634 7840
rect 4724 7772 7604 7800
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 10888 7800 10916 7899
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 7708 7772 10916 7800
rect 7708 7760 7714 7772
rect 4154 7732 4160 7744
rect 3252 7704 4160 7732
rect 4154 7692 4160 7704
rect 4212 7692 4218 7744
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 7742 7732 7748 7744
rect 4396 7704 7748 7732
rect 4396 7692 4402 7704
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 8294 7732 8300 7744
rect 8076 7704 8300 7732
rect 8076 7692 8082 7704
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9306 7732 9312 7744
rect 8720 7704 9312 7732
rect 8720 7692 8726 7704
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 1104 7642 11960 7664
rect 1104 7590 2791 7642
rect 2843 7590 2855 7642
rect 2907 7590 2919 7642
rect 2971 7590 2983 7642
rect 3035 7590 6410 7642
rect 6462 7590 6474 7642
rect 6526 7590 6538 7642
rect 6590 7590 6602 7642
rect 6654 7590 10028 7642
rect 10080 7590 10092 7642
rect 10144 7590 10156 7642
rect 10208 7590 10220 7642
rect 10272 7590 11960 7642
rect 1104 7568 11960 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 6730 7528 6736 7540
rect 2740 7500 6736 7528
rect 2740 7488 2746 7500
rect 6730 7488 6736 7500
rect 6788 7528 6794 7540
rect 9030 7528 9036 7540
rect 6788 7500 9036 7528
rect 6788 7488 6794 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 9732 7500 10548 7528
rect 9732 7488 9738 7500
rect 2041 7463 2099 7469
rect 2041 7429 2053 7463
rect 2087 7460 2099 7463
rect 2087 7432 3832 7460
rect 2087 7429 2099 7432
rect 2041 7423 2099 7429
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 3145 7395 3203 7401
rect 3145 7392 3157 7395
rect 1811 7364 3157 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 3145 7361 3157 7364
rect 3191 7392 3203 7395
rect 3510 7392 3516 7404
rect 3191 7364 3516 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 3694 7392 3700 7404
rect 3655 7364 3700 7392
rect 3694 7352 3700 7364
rect 3752 7352 3758 7404
rect 3804 7392 3832 7432
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 7190 7460 7196 7472
rect 3936 7432 7196 7460
rect 3936 7420 3942 7432
rect 7190 7420 7196 7432
rect 7248 7460 7254 7472
rect 7248 7432 7420 7460
rect 7248 7420 7254 7432
rect 4338 7392 4344 7404
rect 3804 7364 4344 7392
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 5258 7392 5264 7404
rect 4448 7364 5264 7392
rect 1670 7324 1676 7336
rect 1631 7296 1676 7324
rect 1670 7284 1676 7296
rect 1728 7284 1734 7336
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 2501 7327 2559 7333
rect 1995 7296 2452 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2314 7188 2320 7200
rect 2275 7160 2320 7188
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 2424 7188 2452 7296
rect 2501 7293 2513 7327
rect 2547 7293 2559 7327
rect 2682 7324 2688 7336
rect 2643 7296 2688 7324
rect 2501 7287 2559 7293
rect 2516 7256 2544 7287
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 3041 7327 3099 7333
rect 3041 7293 3053 7327
rect 3087 7324 3099 7327
rect 3329 7327 3387 7333
rect 3087 7296 3188 7324
rect 3087 7293 3099 7296
rect 3041 7287 3099 7293
rect 3160 7268 3188 7296
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 4062 7324 4068 7336
rect 3375 7296 4068 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 2774 7256 2780 7268
rect 2516 7228 2780 7256
rect 2774 7216 2780 7228
rect 2832 7216 2838 7268
rect 3142 7216 3148 7268
rect 3200 7216 3206 7268
rect 3344 7188 3372 7287
rect 4062 7284 4068 7296
rect 4120 7324 4126 7336
rect 4448 7324 4476 7364
rect 4120 7296 4476 7324
rect 4525 7327 4583 7333
rect 4120 7284 4126 7296
rect 4525 7293 4537 7327
rect 4571 7293 4583 7327
rect 4890 7324 4896 7336
rect 4851 7296 4896 7324
rect 4525 7287 4583 7293
rect 3510 7216 3516 7268
rect 3568 7256 3574 7268
rect 4540 7256 4568 7287
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 5092 7333 5120 7364
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5592 7364 6561 7392
rect 5592 7352 5598 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7293 5135 7327
rect 5077 7287 5135 7293
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 5626 7324 5632 7336
rect 5224 7296 5269 7324
rect 5587 7296 5632 7324
rect 5224 7284 5230 7296
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 5994 7324 6000 7336
rect 5951 7296 6000 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 5920 7256 5948 7287
rect 5994 7284 6000 7296
rect 6052 7284 6058 7336
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 6457 7327 6515 7333
rect 6457 7293 6469 7327
rect 6503 7324 6515 7327
rect 6730 7324 6736 7336
rect 6503 7296 6736 7324
rect 6503 7293 6515 7296
rect 6457 7287 6515 7293
rect 6104 7256 6132 7287
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 7098 7324 7104 7336
rect 6840 7296 7104 7324
rect 6178 7256 6184 7268
rect 3568 7228 5948 7256
rect 6091 7228 6184 7256
rect 3568 7216 3574 7228
rect 6178 7216 6184 7228
rect 6236 7256 6242 7268
rect 6840 7256 6868 7296
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 7392 7324 7420 7432
rect 7834 7420 7840 7472
rect 7892 7460 7898 7472
rect 9214 7460 9220 7472
rect 7892 7432 9220 7460
rect 7892 7420 7898 7432
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 9306 7420 9312 7472
rect 9364 7460 9370 7472
rect 9364 7432 10456 7460
rect 9364 7420 9370 7432
rect 8018 7392 8024 7404
rect 7944 7364 8024 7392
rect 7944 7333 7972 7364
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 8202 7392 8208 7404
rect 8163 7364 8208 7392
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8846 7392 8852 7404
rect 8807 7364 8852 7392
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9088 7364 9413 7392
rect 9088 7352 9094 7364
rect 9401 7361 9413 7364
rect 9447 7392 9459 7395
rect 10091 7395 10149 7401
rect 10091 7392 10103 7395
rect 9447 7364 10103 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 10091 7361 10103 7364
rect 10137 7392 10149 7395
rect 10318 7392 10324 7404
rect 10137 7364 10324 7392
rect 10137 7361 10149 7364
rect 10091 7355 10149 7361
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 7392 7296 7481 7324
rect 7469 7293 7481 7296
rect 7515 7293 7527 7327
rect 7469 7287 7527 7293
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 8754 7324 8760 7336
rect 8715 7296 8760 7324
rect 7929 7287 7987 7293
rect 6236 7228 6868 7256
rect 6236 7216 6242 7228
rect 6914 7216 6920 7268
rect 6972 7256 6978 7268
rect 7852 7256 7880 7287
rect 8754 7284 8760 7296
rect 8812 7284 8818 7336
rect 9122 7324 9128 7336
rect 9083 7296 9128 7324
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7324 9367 7327
rect 9582 7324 9588 7336
rect 9355 7296 9588 7324
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 10229 7327 10287 7333
rect 10229 7293 10241 7327
rect 10275 7324 10287 7327
rect 10428 7324 10456 7432
rect 10520 7333 10548 7500
rect 10275 7296 10456 7324
rect 10505 7327 10563 7333
rect 10275 7293 10287 7296
rect 10229 7287 10287 7293
rect 10505 7293 10517 7327
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 10778 7324 10784 7336
rect 10652 7296 10697 7324
rect 10739 7296 10784 7324
rect 10652 7284 10658 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 11330 7324 11336 7336
rect 11291 7296 11336 7324
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 6972 7228 8248 7256
rect 6972 7216 6978 7228
rect 2424 7160 3372 7188
rect 4157 7191 4215 7197
rect 4157 7157 4169 7191
rect 4203 7188 4215 7191
rect 5718 7188 5724 7200
rect 4203 7160 5724 7188
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 7101 7191 7159 7197
rect 7101 7157 7113 7191
rect 7147 7188 7159 7191
rect 8110 7188 8116 7200
rect 7147 7160 8116 7188
rect 7147 7157 7159 7160
rect 7101 7151 7159 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8220 7188 8248 7228
rect 9214 7216 9220 7268
rect 9272 7256 9278 7268
rect 11146 7256 11152 7268
rect 9272 7228 11152 7256
rect 9272 7216 9278 7228
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 10965 7191 11023 7197
rect 10965 7188 10977 7191
rect 8220 7160 10977 7188
rect 10965 7157 10977 7160
rect 11011 7157 11023 7191
rect 11422 7188 11428 7200
rect 11383 7160 11428 7188
rect 10965 7151 11023 7157
rect 11422 7148 11428 7160
rect 11480 7148 11486 7200
rect 1104 7098 11960 7120
rect 1104 7046 4600 7098
rect 4652 7046 4664 7098
rect 4716 7046 4728 7098
rect 4780 7046 4792 7098
rect 4844 7046 8219 7098
rect 8271 7046 8283 7098
rect 8335 7046 8347 7098
rect 8399 7046 8411 7098
rect 8463 7046 11960 7098
rect 1104 7024 11960 7046
rect 3528 6956 5212 6984
rect 1670 6876 1676 6928
rect 1728 6916 1734 6928
rect 1728 6888 2728 6916
rect 1728 6876 1734 6888
rect 2700 6857 2728 6888
rect 2774 6876 2780 6928
rect 2832 6916 2838 6928
rect 2832 6888 3188 6916
rect 2832 6876 2838 6888
rect 3160 6860 3188 6888
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6817 2743 6851
rect 3142 6848 3148 6860
rect 3103 6820 3148 6848
rect 2685 6811 2743 6817
rect 2516 6712 2544 6811
rect 2700 6780 2728 6811
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3528 6857 3556 6956
rect 3513 6851 3571 6857
rect 3513 6817 3525 6851
rect 3559 6817 3571 6851
rect 3878 6848 3884 6860
rect 3839 6820 3884 6848
rect 3513 6811 3571 6817
rect 3878 6808 3884 6820
rect 3936 6808 3942 6860
rect 5184 6848 5212 6956
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6822 6984 6828 6996
rect 6052 6956 6828 6984
rect 6052 6944 6058 6956
rect 6822 6944 6828 6956
rect 6880 6984 6886 6996
rect 10594 6984 10600 6996
rect 6880 6956 10600 6984
rect 6880 6944 6886 6956
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 5442 6876 5448 6928
rect 5500 6916 5506 6928
rect 6086 6916 6092 6928
rect 5500 6888 6092 6916
rect 5500 6876 5506 6888
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 6730 6916 6736 6928
rect 6564 6888 6736 6916
rect 6454 6848 6460 6860
rect 3988 6820 4568 6848
rect 5184 6820 6460 6848
rect 3988 6780 4016 6820
rect 4246 6780 4252 6792
rect 2700 6752 4016 6780
rect 4207 6752 4252 6780
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4540 6789 4568 6820
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 6564 6857 6592 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 7392 6888 9260 6916
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6817 6607 6851
rect 6549 6811 6607 6817
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 6917 6851 6975 6857
rect 6696 6820 6741 6848
rect 6696 6808 6702 6820
rect 6917 6817 6929 6851
rect 6963 6848 6975 6851
rect 7392 6848 7420 6888
rect 6963 6820 7420 6848
rect 6963 6817 6975 6820
rect 6917 6811 6975 6817
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 4890 6780 4896 6792
rect 4571 6752 4896 6780
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 4982 6740 4988 6792
rect 5040 6780 5046 6792
rect 5629 6783 5687 6789
rect 5629 6780 5641 6783
rect 5040 6752 5641 6780
rect 5040 6740 5046 6752
rect 5629 6749 5641 6752
rect 5675 6749 5687 6783
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5629 6743 5687 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6086 6740 6092 6792
rect 6144 6780 6150 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 6144 6752 7113 6780
rect 6144 6740 6150 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 3418 6712 3424 6724
rect 2516 6684 3424 6712
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 7208 6712 7236 6820
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 8021 6851 8079 6857
rect 8021 6848 8033 6851
rect 7524 6820 8033 6848
rect 7524 6808 7530 6820
rect 8021 6817 8033 6820
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 8110 6808 8116 6860
rect 8168 6848 8174 6860
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 8168 6820 8217 6848
rect 8168 6808 8174 6820
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 8205 6811 8263 6817
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6848 8539 6851
rect 8570 6848 8576 6860
rect 8527 6820 8576 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 8772 6820 9137 6848
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7558 6780 7564 6792
rect 7519 6752 7564 6780
rect 7377 6743 7435 6749
rect 5868 6684 7236 6712
rect 7392 6712 7420 6743
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 8665 6783 8723 6789
rect 8665 6780 8677 6783
rect 7800 6752 8677 6780
rect 7800 6740 7806 6752
rect 8665 6749 8677 6752
rect 8711 6749 8723 6783
rect 8665 6743 8723 6749
rect 7650 6712 7656 6724
rect 7392 6684 7656 6712
rect 5868 6672 5874 6684
rect 7650 6672 7656 6684
rect 7708 6672 7714 6724
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 5534 6644 5540 6656
rect 2823 6616 5540 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 6270 6604 6276 6656
rect 6328 6644 6334 6656
rect 8772 6644 8800 6820
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 9232 6848 9260 6888
rect 9306 6876 9312 6928
rect 9364 6916 9370 6928
rect 9582 6916 9588 6928
rect 9364 6888 9588 6916
rect 9364 6876 9370 6888
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 9950 6876 9956 6928
rect 10008 6916 10014 6928
rect 11422 6916 11428 6928
rect 10008 6888 11428 6916
rect 10008 6876 10014 6888
rect 11422 6876 11428 6888
rect 11480 6876 11486 6928
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 9232 6820 9505 6848
rect 9125 6811 9183 6817
rect 9493 6817 9505 6820
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 10505 6851 10563 6857
rect 10505 6817 10517 6851
rect 10551 6848 10563 6851
rect 10594 6848 10600 6860
rect 10551 6820 10600 6848
rect 10551 6817 10563 6820
rect 10505 6811 10563 6817
rect 8941 6783 8999 6789
rect 8941 6749 8953 6783
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 8956 6712 8984 6743
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9692 6780 9720 6811
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 10689 6851 10747 6857
rect 10689 6817 10701 6851
rect 10735 6848 10747 6851
rect 10870 6848 10876 6860
rect 10735 6820 10876 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 10042 6780 10048 6792
rect 9088 6752 9720 6780
rect 10003 6752 10048 6780
rect 9088 6740 9094 6752
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 10137 6715 10195 6721
rect 10137 6712 10149 6715
rect 8956 6684 10149 6712
rect 10137 6681 10149 6684
rect 10183 6681 10195 6715
rect 10137 6675 10195 6681
rect 9306 6644 9312 6656
rect 6328 6616 8800 6644
rect 9267 6616 9312 6644
rect 6328 6604 6334 6616
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9493 6647 9551 6653
rect 9493 6613 9505 6647
rect 9539 6644 9551 6647
rect 9815 6647 9873 6653
rect 9815 6644 9827 6647
rect 9539 6616 9827 6644
rect 9539 6613 9551 6616
rect 9493 6607 9551 6613
rect 9815 6613 9827 6616
rect 9861 6613 9873 6647
rect 9815 6607 9873 6613
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10318 6644 10324 6656
rect 9999 6616 10324 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 10778 6644 10784 6656
rect 10739 6616 10784 6644
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 1104 6554 11960 6576
rect 1104 6502 2791 6554
rect 2843 6502 2855 6554
rect 2907 6502 2919 6554
rect 2971 6502 2983 6554
rect 3035 6502 6410 6554
rect 6462 6502 6474 6554
rect 6526 6502 6538 6554
rect 6590 6502 6602 6554
rect 6654 6502 10028 6554
rect 10080 6502 10092 6554
rect 10144 6502 10156 6554
rect 10208 6502 10220 6554
rect 10272 6502 11960 6554
rect 1104 6480 11960 6502
rect 3862 6443 3920 6449
rect 3862 6409 3874 6443
rect 3908 6440 3920 6443
rect 4062 6440 4068 6452
rect 3908 6412 4068 6440
rect 3908 6409 3920 6412
rect 3862 6403 3920 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 10870 6440 10876 6452
rect 4212 6412 4257 6440
rect 6012 6412 10876 6440
rect 4212 6400 4218 6412
rect 3973 6375 4031 6381
rect 3973 6341 3985 6375
rect 4019 6372 4031 6375
rect 6012 6372 6040 6412
rect 10870 6400 10876 6412
rect 10928 6400 10934 6452
rect 10962 6372 10968 6384
rect 4019 6344 6040 6372
rect 6104 6344 7972 6372
rect 4019 6341 4031 6344
rect 3973 6335 4031 6341
rect 6104 6316 6132 6344
rect 3234 6264 3240 6316
rect 3292 6304 3298 6316
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3292 6276 4077 6304
rect 3292 6264 3298 6276
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 6086 6304 6092 6316
rect 5675 6276 6092 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 7944 6313 7972 6344
rect 8220 6344 10968 6372
rect 8220 6313 8248 6344
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 3510 6236 3516 6248
rect 3467 6208 3516 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3510 6196 3516 6208
rect 3568 6236 3574 6248
rect 4982 6236 4988 6248
rect 3568 6208 4988 6236
rect 3568 6196 3574 6208
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5350 6236 5356 6248
rect 5132 6208 5177 6236
rect 5311 6208 5356 6236
rect 5132 6196 5138 6208
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6205 5595 6239
rect 6178 6236 6184 6248
rect 6139 6208 6184 6236
rect 5537 6199 5595 6205
rect 3694 6168 3700 6180
rect 3655 6140 3700 6168
rect 3694 6128 3700 6140
rect 3752 6128 3758 6180
rect 3878 6128 3884 6180
rect 3936 6168 3942 6180
rect 4525 6171 4583 6177
rect 4525 6168 4537 6171
rect 3936 6140 4537 6168
rect 3936 6128 3942 6140
rect 4525 6137 4537 6140
rect 4571 6168 4583 6171
rect 5552 6168 5580 6199
rect 6178 6196 6184 6208
rect 6236 6196 6242 6248
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6328 6208 6469 6236
rect 6328 6196 6334 6208
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6638 6236 6644 6248
rect 6599 6208 6644 6236
rect 6457 6199 6515 6205
rect 6638 6196 6644 6208
rect 6696 6196 6702 6248
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 6788 6208 6960 6236
rect 6788 6196 6794 6208
rect 5810 6168 5816 6180
rect 4571 6140 5816 6168
rect 4571 6137 4583 6140
rect 4525 6131 4583 6137
rect 5810 6128 5816 6140
rect 5868 6128 5874 6180
rect 3513 6103 3571 6109
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 6288 6100 6316 6196
rect 6825 6171 6883 6177
rect 6825 6137 6837 6171
rect 6871 6137 6883 6171
rect 6932 6168 6960 6208
rect 7006 6196 7012 6248
rect 7064 6236 7070 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7064 6208 7297 6236
rect 7064 6196 7070 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6236 7619 6239
rect 7650 6236 7656 6248
rect 7607 6208 7656 6236
rect 7607 6205 7619 6208
rect 7561 6199 7619 6205
rect 7650 6196 7656 6208
rect 7708 6196 7714 6248
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6205 7803 6239
rect 7944 6236 7972 6267
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8904 6276 8953 6304
rect 8904 6264 8910 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 10778 6304 10784 6316
rect 8941 6267 8999 6273
rect 9876 6276 10784 6304
rect 8389 6239 8447 6245
rect 8389 6236 8401 6239
rect 7944 6208 8401 6236
rect 7745 6199 7803 6205
rect 8389 6205 8401 6208
rect 8435 6205 8447 6239
rect 8389 6199 8447 6205
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 9214 6236 9220 6248
rect 9171 6208 9220 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 7760 6168 7788 6199
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9582 6236 9588 6248
rect 9543 6208 9588 6236
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 9876 6245 9904 6276
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9732 6208 9873 6236
rect 9732 6196 9738 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 10321 6239 10379 6245
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 10410 6236 10416 6248
rect 10367 6208 10416 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 8757 6171 8815 6177
rect 8757 6168 8769 6171
rect 6932 6140 8769 6168
rect 6825 6131 6883 6137
rect 8757 6137 8769 6140
rect 8803 6137 8815 6171
rect 8757 6131 8815 6137
rect 3559 6072 6316 6100
rect 6840 6100 6868 6131
rect 7650 6100 7656 6112
rect 6840 6072 7656 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 1104 6010 11960 6032
rect 1104 5958 4600 6010
rect 4652 5958 4664 6010
rect 4716 5958 4728 6010
rect 4780 5958 4792 6010
rect 4844 5958 8219 6010
rect 8271 5958 8283 6010
rect 8335 5958 8347 6010
rect 8399 5958 8411 6010
rect 8463 5958 11960 6010
rect 1104 5936 11960 5958
rect 5350 5856 5356 5908
rect 5408 5896 5414 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 5408 5868 7573 5896
rect 5408 5856 5414 5868
rect 7561 5865 7573 5868
rect 7607 5865 7619 5899
rect 7561 5859 7619 5865
rect 5258 5828 5264 5840
rect 4448 5800 5264 5828
rect 4448 5772 4476 5800
rect 5258 5788 5264 5800
rect 5316 5828 5322 5840
rect 5442 5828 5448 5840
rect 5316 5800 5448 5828
rect 5316 5788 5322 5800
rect 5442 5788 5448 5800
rect 5500 5788 5506 5840
rect 7282 5828 7288 5840
rect 6656 5800 7288 5828
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 4028 5732 4261 5760
rect 4028 5720 4034 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4430 5760 4436 5772
rect 4343 5732 4436 5760
rect 4249 5723 4307 5729
rect 4264 5692 4292 5723
rect 4430 5720 4436 5732
rect 4488 5720 4494 5772
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 5905 5763 5963 5769
rect 5123 5732 5856 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 5626 5692 5632 5704
rect 4264 5664 4384 5692
rect 5587 5664 5632 5692
rect 4356 5624 4384 5664
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 5828 5692 5856 5732
rect 5905 5729 5917 5763
rect 5951 5760 5963 5763
rect 6270 5760 6276 5772
rect 5951 5732 6276 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 5828 5664 6101 5692
rect 6089 5661 6101 5664
rect 6135 5692 6147 5695
rect 6178 5692 6184 5704
rect 6135 5664 6184 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 6178 5652 6184 5664
rect 6236 5692 6242 5704
rect 6546 5692 6552 5704
rect 6236 5664 6552 5692
rect 6236 5652 6242 5664
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 6656 5701 6684 5800
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 8956 5800 9720 5828
rect 6730 5720 6736 5772
rect 6788 5760 6794 5772
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6788 5732 6837 5760
rect 6788 5720 6794 5732
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 7190 5760 7196 5772
rect 7151 5732 7196 5760
rect 6825 5723 6883 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 7742 5760 7748 5772
rect 7703 5732 7748 5760
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 8110 5760 8116 5772
rect 8067 5732 8116 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 8956 5769 8984 5800
rect 9692 5772 9720 5800
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 9309 5763 9367 5769
rect 9309 5729 9321 5763
rect 9355 5760 9367 5763
rect 9398 5760 9404 5772
rect 9355 5732 9404 5760
rect 9355 5729 9367 5732
rect 9309 5723 9367 5729
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 6641 5695 6699 5701
rect 6641 5661 6653 5695
rect 6687 5661 6699 5695
rect 6641 5655 6699 5661
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 6972 5664 7113 5692
rect 6972 5652 6978 5664
rect 7101 5661 7113 5664
rect 7147 5692 7159 5695
rect 7926 5692 7932 5704
rect 7147 5664 7932 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7926 5652 7932 5664
rect 7984 5692 7990 5704
rect 8846 5692 8852 5704
rect 7984 5664 8852 5692
rect 7984 5652 7990 5664
rect 8846 5652 8852 5664
rect 8904 5652 8910 5704
rect 9030 5692 9036 5704
rect 8991 5664 9036 5692
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9214 5692 9220 5704
rect 9175 5664 9220 5692
rect 9214 5652 9220 5664
rect 9272 5692 9278 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9272 5664 9781 5692
rect 9272 5652 9278 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 5810 5624 5816 5636
rect 4356 5596 5816 5624
rect 5810 5584 5816 5596
rect 5868 5584 5874 5636
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 6457 5627 6515 5633
rect 6457 5624 6469 5627
rect 6420 5596 6469 5624
rect 6420 5584 6426 5596
rect 6457 5593 6469 5596
rect 6503 5593 6515 5627
rect 6457 5587 6515 5593
rect 7190 5584 7196 5636
rect 7248 5624 7254 5636
rect 7742 5624 7748 5636
rect 7248 5596 7748 5624
rect 7248 5584 7254 5596
rect 7742 5584 7748 5596
rect 7800 5584 7806 5636
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 10594 5624 10600 5636
rect 8168 5596 10600 5624
rect 8168 5584 8174 5596
rect 10594 5584 10600 5596
rect 10652 5584 10658 5636
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 4525 5559 4583 5565
rect 4525 5556 4537 5559
rect 3752 5528 4537 5556
rect 3752 5516 3758 5528
rect 4525 5525 4537 5528
rect 4571 5556 4583 5559
rect 8018 5556 8024 5568
rect 4571 5528 8024 5556
rect 4571 5525 4583 5528
rect 4525 5519 4583 5525
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 8570 5556 8576 5568
rect 8531 5528 8576 5556
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 1104 5466 11960 5488
rect 1104 5414 2791 5466
rect 2843 5414 2855 5466
rect 2907 5414 2919 5466
rect 2971 5414 2983 5466
rect 3035 5414 6410 5466
rect 6462 5414 6474 5466
rect 6526 5414 6538 5466
rect 6590 5414 6602 5466
rect 6654 5414 10028 5466
rect 10080 5414 10092 5466
rect 10144 5414 10156 5466
rect 10208 5414 10220 5466
rect 10272 5414 11960 5466
rect 1104 5392 11960 5414
rect 6914 5352 6920 5364
rect 5000 5324 6920 5352
rect 5000 5157 5028 5324
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7098 5312 7104 5364
rect 7156 5352 7162 5364
rect 7156 5324 7972 5352
rect 7156 5312 7162 5324
rect 5902 5244 5908 5296
rect 5960 5284 5966 5296
rect 6546 5284 6552 5296
rect 5960 5256 6552 5284
rect 5960 5244 5966 5256
rect 6546 5244 6552 5256
rect 6604 5284 6610 5296
rect 6604 5256 7604 5284
rect 6604 5244 6610 5256
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 7006 5216 7012 5228
rect 6687 5188 7012 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5117 5043 5151
rect 4985 5111 5043 5117
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5117 5319 5151
rect 5718 5148 5724 5160
rect 5679 5120 5724 5148
rect 5261 5111 5319 5117
rect 3510 5040 3516 5092
rect 3568 5080 3574 5092
rect 5276 5080 5304 5111
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 5810 5108 5816 5160
rect 5868 5148 5874 5160
rect 5997 5151 6055 5157
rect 5997 5148 6009 5151
rect 5868 5120 6009 5148
rect 5868 5108 5874 5120
rect 5997 5117 6009 5120
rect 6043 5148 6055 5151
rect 6274 5151 6332 5157
rect 6043 5120 6224 5148
rect 6043 5117 6055 5120
rect 5997 5111 6055 5117
rect 3568 5052 5304 5080
rect 3568 5040 3574 5052
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 6089 5083 6147 5089
rect 6089 5080 6101 5083
rect 5592 5052 6101 5080
rect 5592 5040 5598 5052
rect 6089 5049 6101 5052
rect 6135 5049 6147 5083
rect 6196 5080 6224 5120
rect 6274 5117 6286 5151
rect 6320 5148 6332 5151
rect 6362 5148 6368 5160
rect 6320 5120 6368 5148
rect 6320 5117 6332 5120
rect 6274 5111 6332 5117
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 6730 5148 6736 5160
rect 6564 5120 6736 5148
rect 6564 5080 6592 5120
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5148 7159 5151
rect 7190 5148 7196 5160
rect 7147 5120 7196 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 7466 5148 7472 5160
rect 7423 5120 7472 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 7576 5148 7604 5256
rect 7742 5244 7748 5296
rect 7800 5284 7806 5296
rect 7800 5256 7845 5284
rect 7800 5244 7806 5256
rect 7944 5157 7972 5324
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 9122 5216 9128 5228
rect 8435 5188 9128 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7576 5120 7665 5148
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 6196 5052 6592 5080
rect 6089 5043 6147 5049
rect 3326 4972 3332 5024
rect 3384 5012 3390 5024
rect 3878 5012 3884 5024
rect 3384 4984 3884 5012
rect 3384 4972 3390 4984
rect 3878 4972 3884 4984
rect 3936 5012 3942 5024
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 3936 4984 4813 5012
rect 3936 4972 3942 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 4801 4975 4859 4981
rect 5442 4972 5448 5024
rect 5500 5012 5506 5024
rect 6454 5012 6460 5024
rect 5500 4984 6460 5012
rect 5500 4972 5506 4984
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 6914 5012 6920 5024
rect 6875 4984 6920 5012
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 7668 5012 7696 5111
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 11330 5080 11336 5092
rect 8076 5052 11336 5080
rect 8076 5040 8082 5052
rect 11330 5040 11336 5052
rect 11388 5040 11394 5092
rect 9306 5012 9312 5024
rect 7668 4984 9312 5012
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 1104 4922 11960 4944
rect 1104 4870 4600 4922
rect 4652 4870 4664 4922
rect 4716 4870 4728 4922
rect 4780 4870 4792 4922
rect 4844 4870 8219 4922
rect 8271 4870 8283 4922
rect 8335 4870 8347 4922
rect 8399 4870 8411 4922
rect 8463 4870 11960 4922
rect 1104 4848 11960 4870
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 7282 4808 7288 4820
rect 5767 4780 7288 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 7800 4780 10456 4808
rect 7800 4768 7806 4780
rect 7558 4740 7564 4752
rect 5368 4712 7564 4740
rect 5368 4681 5396 4712
rect 7558 4700 7564 4712
rect 7616 4700 7622 4752
rect 9306 4740 9312 4752
rect 8588 4712 9312 4740
rect 5353 4675 5411 4681
rect 5353 4641 5365 4675
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 5905 4675 5963 4681
rect 5675 4644 5764 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 3602 4564 3608 4616
rect 3660 4604 3666 4616
rect 4062 4604 4068 4616
rect 3660 4576 4068 4604
rect 3660 4564 3666 4576
rect 4062 4564 4068 4576
rect 4120 4604 4126 4616
rect 5736 4604 5764 4644
rect 5905 4641 5917 4675
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6181 4675 6239 4681
rect 6181 4672 6193 4675
rect 6043 4644 6193 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 6181 4641 6193 4644
rect 6227 4641 6239 4675
rect 6454 4672 6460 4684
rect 6415 4644 6460 4672
rect 6181 4635 6239 4641
rect 4120 4576 5764 4604
rect 5920 4604 5948 4635
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6604 4644 7021 4672
rect 6604 4632 6610 4644
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7098 4632 7104 4684
rect 7156 4672 7162 4684
rect 7285 4675 7343 4681
rect 7156 4644 7201 4672
rect 7156 4632 7162 4644
rect 7285 4641 7297 4675
rect 7331 4672 7343 4675
rect 7834 4672 7840 4684
rect 7331 4644 7840 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 8386 4672 8392 4684
rect 8347 4644 8392 4672
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8588 4681 8616 4712
rect 9306 4700 9312 4712
rect 9364 4740 9370 4752
rect 9490 4740 9496 4752
rect 9364 4712 9496 4740
rect 9364 4700 9370 4712
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4641 8631 4675
rect 8573 4635 8631 4641
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8904 4644 8953 4672
rect 8904 4632 8910 4644
rect 8941 4641 8953 4644
rect 8987 4672 8999 4675
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8987 4644 9045 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 10428 4681 10456 4780
rect 10502 4768 10508 4820
rect 10560 4808 10566 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 10560 4780 10885 4808
rect 10560 4768 10566 4780
rect 10873 4777 10885 4780
rect 10919 4777 10931 4811
rect 10873 4771 10931 4777
rect 9861 4675 9919 4681
rect 9861 4672 9873 4675
rect 9180 4644 9873 4672
rect 9180 4632 9186 4644
rect 9861 4641 9873 4644
rect 9907 4672 9919 4675
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 9907 4644 10333 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 6638 4604 6644 4616
rect 5920 4576 6408 4604
rect 6599 4576 6644 4604
rect 4120 4564 4126 4576
rect 5445 4471 5503 4477
rect 5445 4437 5457 4471
rect 5491 4468 5503 4471
rect 5534 4468 5540 4480
rect 5491 4440 5540 4468
rect 5491 4437 5503 4440
rect 5445 4431 5503 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5736 4468 5764 4576
rect 6086 4496 6092 4548
rect 6144 4536 6150 4548
rect 6273 4539 6331 4545
rect 6273 4536 6285 4539
rect 6144 4508 6285 4536
rect 6144 4496 6150 4508
rect 6273 4505 6285 4508
rect 6319 4505 6331 4539
rect 6380 4536 6408 4576
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 7374 4604 7380 4616
rect 6748 4576 7380 4604
rect 6748 4536 6776 4576
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 8754 4604 8760 4616
rect 7791 4576 8760 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 6380 4508 6776 4536
rect 6273 4499 6331 4505
rect 7834 4496 7840 4548
rect 7892 4536 7898 4548
rect 8386 4536 8392 4548
rect 7892 4508 8392 4536
rect 7892 4496 7898 4508
rect 8386 4496 8392 4508
rect 8444 4536 8450 4548
rect 8662 4536 8668 4548
rect 8444 4508 8668 4536
rect 8444 4496 8450 4508
rect 8662 4496 8668 4508
rect 8720 4496 8726 4548
rect 9784 4536 9812 4567
rect 12250 4536 12256 4548
rect 9784 4508 12256 4536
rect 12250 4496 12256 4508
rect 12308 4496 12314 4548
rect 8570 4468 8576 4480
rect 5736 4440 8576 4468
rect 8570 4428 8576 4440
rect 8628 4428 8634 4480
rect 1104 4378 11960 4400
rect 1104 4326 2791 4378
rect 2843 4326 2855 4378
rect 2907 4326 2919 4378
rect 2971 4326 2983 4378
rect 3035 4326 6410 4378
rect 6462 4326 6474 4378
rect 6526 4326 6538 4378
rect 6590 4326 6602 4378
rect 6654 4326 10028 4378
rect 10080 4326 10092 4378
rect 10144 4326 10156 4378
rect 10208 4326 10220 4378
rect 10272 4326 11960 4378
rect 1104 4304 11960 4326
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6328 4236 6561 4264
rect 6328 4224 6334 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 6917 4267 6975 4273
rect 6917 4233 6929 4267
rect 6963 4264 6975 4267
rect 7190 4264 7196 4276
rect 6963 4236 7196 4264
rect 6963 4233 6975 4236
rect 6917 4227 6975 4233
rect 7190 4224 7196 4236
rect 7248 4224 7254 4276
rect 8481 4267 8539 4273
rect 8481 4233 8493 4267
rect 8527 4264 8539 4267
rect 8938 4264 8944 4276
rect 8527 4236 8944 4264
rect 8527 4233 8539 4236
rect 8481 4227 8539 4233
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 5534 4156 5540 4208
rect 5592 4196 5598 4208
rect 6822 4196 6828 4208
rect 5592 4168 6828 4196
rect 5592 4156 5598 4168
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 8864 4168 9260 4196
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5994 4128 6000 4140
rect 5040 4100 6000 4128
rect 5040 4088 5046 4100
rect 5994 4088 6000 4100
rect 6052 4128 6058 4140
rect 8864 4128 8892 4168
rect 6052 4100 8892 4128
rect 8941 4131 8999 4137
rect 6052 4088 6058 4100
rect 8941 4097 8953 4131
rect 8987 4097 8999 4131
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 8941 4091 8999 4097
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 6457 4063 6515 4069
rect 6457 4060 6469 4063
rect 6236 4032 6469 4060
rect 6236 4020 6242 4032
rect 6457 4029 6469 4032
rect 6503 4029 6515 4063
rect 6822 4060 6828 4072
rect 6783 4032 6828 4060
rect 6457 4023 6515 4029
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 8846 4060 8852 4072
rect 8807 4032 8852 4060
rect 8846 4020 8852 4032
rect 8904 4020 8910 4072
rect 6086 3952 6092 4004
rect 6144 3992 6150 4004
rect 7834 3992 7840 4004
rect 6144 3964 7840 3992
rect 6144 3952 6150 3964
rect 7834 3952 7840 3964
rect 7892 3952 7898 4004
rect 8956 3992 8984 4091
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9232 4069 9260 4168
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 10778 3992 10784 4004
rect 8956 3964 10784 3992
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 1104 3834 11960 3856
rect 1104 3782 4600 3834
rect 4652 3782 4664 3834
rect 4716 3782 4728 3834
rect 4780 3782 4792 3834
rect 4844 3782 8219 3834
rect 8271 3782 8283 3834
rect 8335 3782 8347 3834
rect 8399 3782 8411 3834
rect 8463 3782 11960 3834
rect 1104 3760 11960 3782
rect 4430 3652 4436 3664
rect 1412 3624 4436 3652
rect 1412 3593 1440 3624
rect 4430 3612 4436 3624
rect 4488 3612 4494 3664
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 4246 3584 4252 3596
rect 2455 3556 4252 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 658 3340 664 3392
rect 716 3380 722 3392
rect 1581 3383 1639 3389
rect 1581 3380 1593 3383
rect 716 3352 1593 3380
rect 716 3340 722 3352
rect 1581 3349 1593 3352
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2593 3383 2651 3389
rect 2593 3380 2605 3383
rect 2096 3352 2605 3380
rect 2096 3340 2102 3352
rect 2593 3349 2605 3352
rect 2639 3349 2651 3383
rect 2593 3343 2651 3349
rect 1104 3290 11960 3312
rect 1104 3238 2791 3290
rect 2843 3238 2855 3290
rect 2907 3238 2919 3290
rect 2971 3238 2983 3290
rect 3035 3238 6410 3290
rect 6462 3238 6474 3290
rect 6526 3238 6538 3290
rect 6590 3238 6602 3290
rect 6654 3238 10028 3290
rect 10080 3238 10092 3290
rect 10144 3238 10156 3290
rect 10208 3238 10220 3290
rect 10272 3238 11960 3290
rect 1104 3216 11960 3238
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2972 7711 2975
rect 7834 2972 7840 2984
rect 7699 2944 7840 2972
rect 7699 2941 7711 2944
rect 7653 2935 7711 2941
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 7834 2836 7840 2848
rect 7795 2808 7840 2836
rect 7834 2796 7840 2808
rect 7892 2796 7898 2848
rect 1104 2746 11960 2768
rect 1104 2694 4600 2746
rect 4652 2694 4664 2746
rect 4716 2694 4728 2746
rect 4780 2694 4792 2746
rect 4844 2694 8219 2746
rect 8271 2694 8283 2746
rect 8335 2694 8347 2746
rect 8399 2694 8411 2746
rect 8463 2694 11960 2746
rect 1104 2672 11960 2694
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2496 7067 2499
rect 7650 2496 7656 2508
rect 7055 2468 7656 2496
rect 7055 2465 7067 2468
rect 7009 2459 7067 2465
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 6730 2252 6736 2304
rect 6788 2292 6794 2304
rect 7101 2295 7159 2301
rect 7101 2292 7113 2295
rect 6788 2264 7113 2292
rect 6788 2252 6794 2264
rect 7101 2261 7113 2264
rect 7147 2261 7159 2295
rect 7101 2255 7159 2261
rect 1104 2202 11960 2224
rect 1104 2150 2791 2202
rect 2843 2150 2855 2202
rect 2907 2150 2919 2202
rect 2971 2150 2983 2202
rect 3035 2150 6410 2202
rect 6462 2150 6474 2202
rect 6526 2150 6538 2202
rect 6590 2150 6602 2202
rect 6654 2150 10028 2202
rect 10080 2150 10092 2202
rect 10144 2150 10156 2202
rect 10208 2150 10220 2202
rect 10272 2150 11960 2202
rect 1104 2128 11960 2150
<< via1 >>
rect 2791 13030 2843 13082
rect 2855 13030 2907 13082
rect 2919 13030 2971 13082
rect 2983 13030 3035 13082
rect 6410 13030 6462 13082
rect 6474 13030 6526 13082
rect 6538 13030 6590 13082
rect 6602 13030 6654 13082
rect 10028 13030 10080 13082
rect 10092 13030 10144 13082
rect 10156 13030 10208 13082
rect 10220 13030 10272 13082
rect 7840 12724 7892 12776
rect 6920 12588 6972 12640
rect 4600 12486 4652 12538
rect 4664 12486 4716 12538
rect 4728 12486 4780 12538
rect 4792 12486 4844 12538
rect 8219 12486 8271 12538
rect 8283 12486 8335 12538
rect 8347 12486 8399 12538
rect 8411 12486 8463 12538
rect 2791 11942 2843 11994
rect 2855 11942 2907 11994
rect 2919 11942 2971 11994
rect 2983 11942 3035 11994
rect 6410 11942 6462 11994
rect 6474 11942 6526 11994
rect 6538 11942 6590 11994
rect 6602 11942 6654 11994
rect 10028 11942 10080 11994
rect 10092 11942 10144 11994
rect 10156 11942 10208 11994
rect 10220 11942 10272 11994
rect 2044 11704 2096 11756
rect 4344 11704 4396 11756
rect 4988 11704 5040 11756
rect 7104 11704 7156 11756
rect 3516 11636 3568 11688
rect 4160 11500 4212 11552
rect 4600 11398 4652 11450
rect 4664 11398 4716 11450
rect 4728 11398 4780 11450
rect 4792 11398 4844 11450
rect 8219 11398 8271 11450
rect 8283 11398 8335 11450
rect 8347 11398 8399 11450
rect 8411 11398 8463 11450
rect 664 11024 716 11076
rect 5356 11024 5408 11076
rect 10508 11024 10560 11076
rect 12256 11024 12308 11076
rect 2791 10854 2843 10906
rect 2855 10854 2907 10906
rect 2919 10854 2971 10906
rect 2983 10854 3035 10906
rect 6410 10854 6462 10906
rect 6474 10854 6526 10906
rect 6538 10854 6590 10906
rect 6602 10854 6654 10906
rect 10028 10854 10080 10906
rect 10092 10854 10144 10906
rect 10156 10854 10208 10906
rect 10220 10854 10272 10906
rect 9312 10752 9364 10804
rect 8668 10684 8720 10736
rect 6736 10616 6788 10668
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 7196 10548 7248 10600
rect 7380 10523 7432 10532
rect 7380 10489 7389 10523
rect 7389 10489 7423 10523
rect 7423 10489 7432 10523
rect 7380 10480 7432 10489
rect 6184 10412 6236 10464
rect 6276 10412 6328 10464
rect 6736 10412 6788 10464
rect 4600 10310 4652 10362
rect 4664 10310 4716 10362
rect 4728 10310 4780 10362
rect 4792 10310 4844 10362
rect 8219 10310 8271 10362
rect 8283 10310 8335 10362
rect 8347 10310 8399 10362
rect 8411 10310 8463 10362
rect 8024 10208 8076 10260
rect 7288 10140 7340 10192
rect 7932 10140 7984 10192
rect 5356 10115 5408 10124
rect 5356 10081 5365 10115
rect 5365 10081 5399 10115
rect 5399 10081 5408 10115
rect 5356 10072 5408 10081
rect 5172 10004 5224 10056
rect 6368 10072 6420 10124
rect 6920 10072 6972 10124
rect 7748 10072 7800 10124
rect 6184 10004 6236 10056
rect 6828 10004 6880 10056
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 8760 10004 8812 10056
rect 7012 9936 7064 9988
rect 5632 9868 5684 9920
rect 6092 9868 6144 9920
rect 7472 9868 7524 9920
rect 7564 9868 7616 9920
rect 2791 9766 2843 9818
rect 2855 9766 2907 9818
rect 2919 9766 2971 9818
rect 2983 9766 3035 9818
rect 6410 9766 6462 9818
rect 6474 9766 6526 9818
rect 6538 9766 6590 9818
rect 6602 9766 6654 9818
rect 10028 9766 10080 9818
rect 10092 9766 10144 9818
rect 10156 9766 10208 9818
rect 10220 9766 10272 9818
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 5080 9639 5132 9648
rect 5080 9605 5089 9639
rect 5089 9605 5123 9639
rect 5123 9605 5132 9639
rect 5080 9596 5132 9605
rect 7380 9664 7432 9716
rect 7656 9664 7708 9716
rect 7748 9664 7800 9716
rect 7932 9664 7984 9716
rect 5540 9596 5592 9648
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 5264 9528 5316 9580
rect 6184 9571 6236 9580
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6184 9528 6236 9537
rect 9680 9596 9732 9648
rect 8208 9528 8260 9580
rect 9864 9528 9916 9580
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 3240 9460 3292 9512
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 5448 9460 5500 9512
rect 6460 9503 6512 9512
rect 6460 9469 6469 9503
rect 6469 9469 6503 9503
rect 6503 9469 6512 9503
rect 6460 9460 6512 9469
rect 7288 9460 7340 9512
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 8116 9460 8168 9512
rect 9036 9460 9088 9512
rect 10784 9460 10836 9512
rect 7932 9392 7984 9444
rect 3608 9324 3660 9376
rect 3700 9324 3752 9376
rect 6920 9324 6972 9376
rect 8852 9367 8904 9376
rect 8852 9333 8861 9367
rect 8861 9333 8895 9367
rect 8895 9333 8904 9367
rect 8852 9324 8904 9333
rect 4600 9222 4652 9274
rect 4664 9222 4716 9274
rect 4728 9222 4780 9274
rect 4792 9222 4844 9274
rect 8219 9222 8271 9274
rect 8283 9222 8335 9274
rect 8347 9222 8399 9274
rect 8411 9222 8463 9274
rect 9588 9120 9640 9172
rect 10416 9120 10468 9172
rect 5632 9052 5684 9104
rect 3516 8984 3568 9036
rect 4160 8984 4212 9036
rect 5448 9027 5500 9036
rect 5448 8993 5457 9027
rect 5457 8993 5491 9027
rect 5491 8993 5500 9027
rect 5448 8984 5500 8993
rect 5724 9027 5776 9036
rect 5724 8993 5733 9027
rect 5733 8993 5767 9027
rect 5767 8993 5776 9027
rect 5724 8984 5776 8993
rect 6460 9027 6512 9036
rect 4068 8848 4120 8900
rect 5264 8916 5316 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 6460 8993 6469 9027
rect 6469 8993 6503 9027
rect 6503 8993 6512 9027
rect 6460 8984 6512 8993
rect 6920 9052 6972 9104
rect 7196 9052 7248 9104
rect 7564 8984 7616 9036
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7104 8916 7156 8925
rect 7196 8916 7248 8968
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 8116 9052 8168 9104
rect 9128 8984 9180 9036
rect 9772 8984 9824 9036
rect 8944 8916 8996 8968
rect 3240 8823 3292 8832
rect 3240 8789 3249 8823
rect 3249 8789 3283 8823
rect 3283 8789 3292 8823
rect 3240 8780 3292 8789
rect 3976 8780 4028 8832
rect 8576 8848 8628 8900
rect 8760 8848 8812 8900
rect 10324 8848 10376 8900
rect 5540 8780 5592 8832
rect 7196 8780 7248 8832
rect 7288 8780 7340 8832
rect 2791 8678 2843 8730
rect 2855 8678 2907 8730
rect 2919 8678 2971 8730
rect 2983 8678 3035 8730
rect 6410 8678 6462 8730
rect 6474 8678 6526 8730
rect 6538 8678 6590 8730
rect 6602 8678 6654 8730
rect 10028 8678 10080 8730
rect 10092 8678 10144 8730
rect 10156 8678 10208 8730
rect 10220 8678 10272 8730
rect 3792 8576 3844 8628
rect 7196 8576 7248 8628
rect 8944 8576 8996 8628
rect 9036 8576 9088 8628
rect 10324 8619 10376 8628
rect 5448 8508 5500 8560
rect 4160 8440 4212 8492
rect 5632 8440 5684 8492
rect 9128 8508 9180 8560
rect 10324 8585 10333 8619
rect 10333 8585 10367 8619
rect 10367 8585 10376 8619
rect 10324 8576 10376 8585
rect 9956 8551 10008 8560
rect 9956 8517 9965 8551
rect 9965 8517 9999 8551
rect 9999 8517 10008 8551
rect 9956 8508 10008 8517
rect 3976 8415 4028 8424
rect 3424 8304 3476 8356
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 4436 8372 4488 8424
rect 5816 8372 5868 8424
rect 7104 8372 7156 8424
rect 7196 8372 7248 8424
rect 8852 8483 8904 8492
rect 8852 8449 8861 8483
rect 8861 8449 8895 8483
rect 8895 8449 8904 8483
rect 8852 8440 8904 8449
rect 7748 8415 7800 8424
rect 7748 8381 7757 8415
rect 7757 8381 7791 8415
rect 7791 8381 7800 8415
rect 7748 8372 7800 8381
rect 7840 8372 7892 8424
rect 4160 8304 4212 8356
rect 6184 8304 6236 8356
rect 4344 8236 4396 8288
rect 4896 8236 4948 8288
rect 6920 8304 6972 8356
rect 9128 8372 9180 8424
rect 10508 8415 10560 8424
rect 7932 8236 7984 8288
rect 8760 8236 8812 8288
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 9588 8304 9640 8356
rect 9496 8236 9548 8288
rect 9956 8236 10008 8288
rect 4600 8134 4652 8186
rect 4664 8134 4716 8186
rect 4728 8134 4780 8186
rect 4792 8134 4844 8186
rect 8219 8134 8271 8186
rect 8283 8134 8335 8186
rect 8347 8134 8399 8186
rect 8411 8134 8463 8186
rect 4252 8032 4304 8084
rect 2412 8007 2464 8016
rect 2412 7973 2421 8007
rect 2421 7973 2455 8007
rect 2455 7973 2464 8007
rect 2412 7964 2464 7973
rect 3700 7964 3752 8016
rect 4344 7964 4396 8016
rect 5080 8032 5132 8084
rect 8576 8075 8628 8084
rect 3608 7939 3660 7948
rect 3608 7905 3617 7939
rect 3617 7905 3651 7939
rect 3651 7905 3660 7939
rect 3608 7896 3660 7905
rect 5264 7939 5316 7948
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3516 7871 3568 7880
rect 3332 7828 3384 7837
rect 3516 7837 3525 7871
rect 3525 7837 3559 7871
rect 3559 7837 3568 7871
rect 3516 7828 3568 7837
rect 4160 7828 4212 7880
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 5540 7939 5592 7948
rect 5540 7905 5549 7939
rect 5549 7905 5583 7939
rect 5583 7905 5592 7939
rect 5540 7896 5592 7905
rect 5172 7828 5224 7880
rect 6368 7896 6420 7948
rect 7012 7896 7064 7948
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 7748 7896 7800 7948
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 8668 8032 8720 8084
rect 9864 8032 9916 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 8392 7964 8444 8016
rect 8944 7964 8996 8016
rect 8208 7896 8260 7948
rect 8576 7828 8628 7880
rect 9772 7896 9824 7948
rect 10692 7896 10744 7948
rect 11152 7939 11204 7948
rect 7656 7760 7708 7812
rect 11152 7905 11161 7939
rect 11161 7905 11195 7939
rect 11195 7905 11204 7939
rect 11152 7896 11204 7905
rect 4160 7692 4212 7744
rect 4344 7692 4396 7744
rect 7748 7692 7800 7744
rect 8024 7692 8076 7744
rect 8300 7692 8352 7744
rect 8668 7692 8720 7744
rect 9312 7692 9364 7744
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 2791 7590 2843 7642
rect 2855 7590 2907 7642
rect 2919 7590 2971 7642
rect 2983 7590 3035 7642
rect 6410 7590 6462 7642
rect 6474 7590 6526 7642
rect 6538 7590 6590 7642
rect 6602 7590 6654 7642
rect 10028 7590 10080 7642
rect 10092 7590 10144 7642
rect 10156 7590 10208 7642
rect 10220 7590 10272 7642
rect 2688 7488 2740 7540
rect 6736 7488 6788 7540
rect 9036 7488 9088 7540
rect 9680 7488 9732 7540
rect 3516 7352 3568 7404
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 3884 7420 3936 7472
rect 7196 7420 7248 7472
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 2320 7191 2372 7200
rect 2320 7157 2329 7191
rect 2329 7157 2363 7191
rect 2363 7157 2372 7191
rect 2320 7148 2372 7157
rect 2688 7327 2740 7336
rect 2688 7293 2697 7327
rect 2697 7293 2731 7327
rect 2731 7293 2740 7327
rect 2688 7284 2740 7293
rect 2780 7216 2832 7268
rect 3148 7216 3200 7268
rect 4068 7284 4120 7336
rect 4896 7327 4948 7336
rect 3516 7216 3568 7268
rect 4896 7293 4905 7327
rect 4905 7293 4939 7327
rect 4939 7293 4948 7327
rect 4896 7284 4948 7293
rect 5264 7352 5316 7404
rect 5540 7352 5592 7404
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5632 7327 5684 7336
rect 5172 7284 5224 7293
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 6000 7284 6052 7336
rect 6736 7284 6788 7336
rect 6184 7216 6236 7268
rect 7104 7284 7156 7336
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 7840 7420 7892 7472
rect 9220 7420 9272 7472
rect 9312 7420 9364 7472
rect 8024 7352 8076 7404
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 9036 7352 9088 7404
rect 10324 7352 10376 7404
rect 8760 7327 8812 7336
rect 6920 7216 6972 7268
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 9588 7284 9640 7336
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 10600 7327 10652 7336
rect 10600 7293 10609 7327
rect 10609 7293 10643 7327
rect 10643 7293 10652 7327
rect 10784 7327 10836 7336
rect 10600 7284 10652 7293
rect 10784 7293 10793 7327
rect 10793 7293 10827 7327
rect 10827 7293 10836 7327
rect 10784 7284 10836 7293
rect 11336 7327 11388 7336
rect 11336 7293 11345 7327
rect 11345 7293 11379 7327
rect 11379 7293 11388 7327
rect 11336 7284 11388 7293
rect 5724 7148 5776 7200
rect 8116 7148 8168 7200
rect 9220 7216 9272 7268
rect 11152 7216 11204 7268
rect 11428 7191 11480 7200
rect 11428 7157 11437 7191
rect 11437 7157 11471 7191
rect 11471 7157 11480 7191
rect 11428 7148 11480 7157
rect 4600 7046 4652 7098
rect 4664 7046 4716 7098
rect 4728 7046 4780 7098
rect 4792 7046 4844 7098
rect 8219 7046 8271 7098
rect 8283 7046 8335 7098
rect 8347 7046 8399 7098
rect 8411 7046 8463 7098
rect 1676 6876 1728 6928
rect 2780 6876 2832 6928
rect 3148 6851 3200 6860
rect 3148 6817 3157 6851
rect 3157 6817 3191 6851
rect 3191 6817 3200 6851
rect 3148 6808 3200 6817
rect 3884 6851 3936 6860
rect 3884 6817 3893 6851
rect 3893 6817 3927 6851
rect 3927 6817 3936 6851
rect 3884 6808 3936 6817
rect 6000 6944 6052 6996
rect 6828 6944 6880 6996
rect 10600 6944 10652 6996
rect 5448 6876 5500 6928
rect 6092 6876 6144 6928
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 6460 6808 6512 6860
rect 6736 6876 6788 6928
rect 6644 6851 6696 6860
rect 6644 6817 6653 6851
rect 6653 6817 6687 6851
rect 6687 6817 6696 6851
rect 6644 6808 6696 6817
rect 4896 6740 4948 6792
rect 4988 6740 5040 6792
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6092 6740 6144 6792
rect 3424 6672 3476 6724
rect 5816 6672 5868 6724
rect 7472 6808 7524 6860
rect 8116 6808 8168 6860
rect 8576 6808 8628 6860
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 7748 6740 7800 6792
rect 7656 6672 7708 6724
rect 5540 6604 5592 6656
rect 6276 6604 6328 6656
rect 9312 6876 9364 6928
rect 9588 6876 9640 6928
rect 9956 6876 10008 6928
rect 11428 6876 11480 6928
rect 9036 6740 9088 6792
rect 10600 6808 10652 6860
rect 10876 6808 10928 6860
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 10324 6604 10376 6656
rect 10784 6647 10836 6656
rect 10784 6613 10793 6647
rect 10793 6613 10827 6647
rect 10827 6613 10836 6647
rect 10784 6604 10836 6613
rect 2791 6502 2843 6554
rect 2855 6502 2907 6554
rect 2919 6502 2971 6554
rect 2983 6502 3035 6554
rect 6410 6502 6462 6554
rect 6474 6502 6526 6554
rect 6538 6502 6590 6554
rect 6602 6502 6654 6554
rect 10028 6502 10080 6554
rect 10092 6502 10144 6554
rect 10156 6502 10208 6554
rect 10220 6502 10272 6554
rect 4068 6400 4120 6452
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 10876 6400 10928 6452
rect 3240 6264 3292 6316
rect 6092 6264 6144 6316
rect 10968 6332 11020 6384
rect 3516 6196 3568 6248
rect 4988 6196 5040 6248
rect 5080 6239 5132 6248
rect 5080 6205 5089 6239
rect 5089 6205 5123 6239
rect 5123 6205 5132 6239
rect 5356 6239 5408 6248
rect 5080 6196 5132 6205
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 6184 6239 6236 6248
rect 3700 6171 3752 6180
rect 3700 6137 3709 6171
rect 3709 6137 3743 6171
rect 3743 6137 3752 6171
rect 3700 6128 3752 6137
rect 3884 6128 3936 6180
rect 6184 6205 6193 6239
rect 6193 6205 6227 6239
rect 6227 6205 6236 6239
rect 6184 6196 6236 6205
rect 6276 6196 6328 6248
rect 6644 6239 6696 6248
rect 6644 6205 6653 6239
rect 6653 6205 6687 6239
rect 6687 6205 6696 6239
rect 6644 6196 6696 6205
rect 6736 6196 6788 6248
rect 5816 6128 5868 6180
rect 7012 6196 7064 6248
rect 7656 6196 7708 6248
rect 8852 6264 8904 6316
rect 9220 6196 9272 6248
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 9680 6196 9732 6248
rect 10784 6264 10836 6316
rect 10416 6196 10468 6248
rect 7656 6060 7708 6112
rect 4600 5958 4652 6010
rect 4664 5958 4716 6010
rect 4728 5958 4780 6010
rect 4792 5958 4844 6010
rect 8219 5958 8271 6010
rect 8283 5958 8335 6010
rect 8347 5958 8399 6010
rect 8411 5958 8463 6010
rect 5356 5856 5408 5908
rect 5264 5788 5316 5840
rect 5448 5788 5500 5840
rect 3976 5720 4028 5772
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 5632 5695 5684 5704
rect 5632 5661 5641 5695
rect 5641 5661 5675 5695
rect 5675 5661 5684 5695
rect 5632 5652 5684 5661
rect 6276 5720 6328 5772
rect 6184 5652 6236 5704
rect 6552 5652 6604 5704
rect 7288 5788 7340 5840
rect 6736 5720 6788 5772
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 8116 5720 8168 5772
rect 9404 5720 9456 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 6920 5652 6972 5704
rect 7932 5652 7984 5704
rect 8852 5652 8904 5704
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 5816 5584 5868 5636
rect 6368 5584 6420 5636
rect 7196 5584 7248 5636
rect 7748 5584 7800 5636
rect 8116 5584 8168 5636
rect 10600 5584 10652 5636
rect 3700 5516 3752 5568
rect 8024 5516 8076 5568
rect 8576 5559 8628 5568
rect 8576 5525 8585 5559
rect 8585 5525 8619 5559
rect 8619 5525 8628 5559
rect 8576 5516 8628 5525
rect 2791 5414 2843 5466
rect 2855 5414 2907 5466
rect 2919 5414 2971 5466
rect 2983 5414 3035 5466
rect 6410 5414 6462 5466
rect 6474 5414 6526 5466
rect 6538 5414 6590 5466
rect 6602 5414 6654 5466
rect 10028 5414 10080 5466
rect 10092 5414 10144 5466
rect 10156 5414 10208 5466
rect 10220 5414 10272 5466
rect 6920 5312 6972 5364
rect 7104 5312 7156 5364
rect 5908 5244 5960 5296
rect 6552 5244 6604 5296
rect 7012 5176 7064 5228
rect 5724 5151 5776 5160
rect 3516 5040 3568 5092
rect 5724 5117 5733 5151
rect 5733 5117 5767 5151
rect 5767 5117 5776 5151
rect 5724 5108 5776 5117
rect 5816 5108 5868 5160
rect 5540 5040 5592 5092
rect 6368 5108 6420 5160
rect 6736 5108 6788 5160
rect 7196 5108 7248 5160
rect 7472 5108 7524 5160
rect 7748 5287 7800 5296
rect 7748 5253 7757 5287
rect 7757 5253 7791 5287
rect 7791 5253 7800 5287
rect 7748 5244 7800 5253
rect 9128 5176 9180 5228
rect 3332 4972 3384 5024
rect 3884 4972 3936 5024
rect 5448 4972 5500 5024
rect 6460 4972 6512 5024
rect 6920 5015 6972 5024
rect 6920 4981 6929 5015
rect 6929 4981 6963 5015
rect 6963 4981 6972 5015
rect 6920 4972 6972 4981
rect 8024 5040 8076 5092
rect 11336 5040 11388 5092
rect 9312 4972 9364 5024
rect 4600 4870 4652 4922
rect 4664 4870 4716 4922
rect 4728 4870 4780 4922
rect 4792 4870 4844 4922
rect 8219 4870 8271 4922
rect 8283 4870 8335 4922
rect 8347 4870 8399 4922
rect 8411 4870 8463 4922
rect 7288 4768 7340 4820
rect 7748 4768 7800 4820
rect 7564 4700 7616 4752
rect 3608 4564 3660 4616
rect 4068 4564 4120 4616
rect 6460 4675 6512 4684
rect 6460 4641 6469 4675
rect 6469 4641 6503 4675
rect 6503 4641 6512 4675
rect 6460 4632 6512 4641
rect 6552 4632 6604 4684
rect 7104 4675 7156 4684
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 7840 4632 7892 4684
rect 8392 4675 8444 4684
rect 8392 4641 8401 4675
rect 8401 4641 8435 4675
rect 8435 4641 8444 4675
rect 8392 4632 8444 4641
rect 9312 4700 9364 4752
rect 9496 4700 9548 4752
rect 8852 4632 8904 4684
rect 9128 4675 9180 4684
rect 9128 4641 9137 4675
rect 9137 4641 9171 4675
rect 9171 4641 9180 4675
rect 10508 4768 10560 4820
rect 9128 4632 9180 4641
rect 6644 4607 6696 4616
rect 5540 4428 5592 4480
rect 6092 4496 6144 4548
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7380 4564 7432 4616
rect 8760 4564 8812 4616
rect 7840 4496 7892 4548
rect 8392 4496 8444 4548
rect 8668 4496 8720 4548
rect 12256 4496 12308 4548
rect 8576 4428 8628 4480
rect 2791 4326 2843 4378
rect 2855 4326 2907 4378
rect 2919 4326 2971 4378
rect 2983 4326 3035 4378
rect 6410 4326 6462 4378
rect 6474 4326 6526 4378
rect 6538 4326 6590 4378
rect 6602 4326 6654 4378
rect 10028 4326 10080 4378
rect 10092 4326 10144 4378
rect 10156 4326 10208 4378
rect 10220 4326 10272 4378
rect 6276 4224 6328 4276
rect 7196 4224 7248 4276
rect 8944 4224 8996 4276
rect 5540 4156 5592 4208
rect 6828 4156 6880 4208
rect 4988 4088 5040 4140
rect 6000 4088 6052 4140
rect 9128 4131 9180 4140
rect 6184 4020 6236 4072
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 8852 4063 8904 4072
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 6092 3952 6144 4004
rect 7840 3952 7892 4004
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 10784 3952 10836 4004
rect 4600 3782 4652 3834
rect 4664 3782 4716 3834
rect 4728 3782 4780 3834
rect 4792 3782 4844 3834
rect 8219 3782 8271 3834
rect 8283 3782 8335 3834
rect 8347 3782 8399 3834
rect 8411 3782 8463 3834
rect 4436 3612 4488 3664
rect 4252 3544 4304 3596
rect 664 3340 716 3392
rect 2044 3340 2096 3392
rect 2791 3238 2843 3290
rect 2855 3238 2907 3290
rect 2919 3238 2971 3290
rect 2983 3238 3035 3290
rect 6410 3238 6462 3290
rect 6474 3238 6526 3290
rect 6538 3238 6590 3290
rect 6602 3238 6654 3290
rect 10028 3238 10080 3290
rect 10092 3238 10144 3290
rect 10156 3238 10208 3290
rect 10220 3238 10272 3290
rect 7840 2932 7892 2984
rect 7840 2839 7892 2848
rect 7840 2805 7849 2839
rect 7849 2805 7883 2839
rect 7883 2805 7892 2839
rect 7840 2796 7892 2805
rect 4600 2694 4652 2746
rect 4664 2694 4716 2746
rect 4728 2694 4780 2746
rect 4792 2694 4844 2746
rect 8219 2694 8271 2746
rect 8283 2694 8335 2746
rect 8347 2694 8399 2746
rect 8411 2694 8463 2746
rect 7656 2456 7708 2508
rect 6736 2252 6788 2304
rect 2791 2150 2843 2202
rect 2855 2150 2907 2202
rect 2919 2150 2971 2202
rect 2983 2150 3035 2202
rect 6410 2150 6462 2202
rect 6474 2150 6526 2202
rect 6538 2150 6590 2202
rect 6602 2150 6654 2202
rect 10028 2150 10080 2202
rect 10092 2150 10144 2202
rect 10156 2150 10208 2202
rect 10220 2150 10272 2202
<< metal2 >>
rect 662 14440 718 15240
rect 2042 14440 2098 15240
rect 3514 14440 3570 15240
rect 4986 14440 5042 15240
rect 6458 14440 6514 15240
rect 7838 14440 7894 15240
rect 9310 14440 9366 15240
rect 10782 14440 10838 15240
rect 12254 14440 12310 15240
rect 676 11082 704 14440
rect 2056 11762 2084 14440
rect 3422 13968 3478 13977
rect 3422 13903 3478 13912
rect 2765 13084 3061 13104
rect 2821 13082 2845 13084
rect 2901 13082 2925 13084
rect 2981 13082 3005 13084
rect 2843 13030 2845 13082
rect 2907 13030 2919 13082
rect 2981 13030 2983 13082
rect 2821 13028 2845 13030
rect 2901 13028 2925 13030
rect 2981 13028 3005 13030
rect 2765 13008 3061 13028
rect 2765 11996 3061 12016
rect 2821 11994 2845 11996
rect 2901 11994 2925 11996
rect 2981 11994 3005 11996
rect 2843 11942 2845 11994
rect 2907 11942 2919 11994
rect 2981 11942 2983 11994
rect 2821 11940 2845 11942
rect 2901 11940 2925 11942
rect 2981 11940 3005 11942
rect 2765 11920 3061 11940
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1950 11384 2006 11393
rect 1950 11319 2006 11328
rect 664 11076 716 11082
rect 664 11018 716 11024
rect 1964 9518 1992 11319
rect 2765 10908 3061 10928
rect 2821 10906 2845 10908
rect 2901 10906 2925 10908
rect 2981 10906 3005 10908
rect 2843 10854 2845 10906
rect 2907 10854 2919 10906
rect 2981 10854 2983 10906
rect 2821 10852 2845 10854
rect 2901 10852 2925 10854
rect 2981 10852 3005 10854
rect 2765 10832 3061 10852
rect 2765 9820 3061 9840
rect 2821 9818 2845 9820
rect 2901 9818 2925 9820
rect 2981 9818 3005 9820
rect 2843 9766 2845 9818
rect 2907 9766 2919 9818
rect 2981 9766 2983 9818
rect 2821 9764 2845 9766
rect 2901 9764 2925 9766
rect 2981 9764 3005 9766
rect 2765 9744 3061 9764
rect 3436 9586 3464 13903
rect 3528 11694 3556 14440
rect 4574 12540 4870 12560
rect 4630 12538 4654 12540
rect 4710 12538 4734 12540
rect 4790 12538 4814 12540
rect 4652 12486 4654 12538
rect 4716 12486 4728 12538
rect 4790 12486 4792 12538
rect 4630 12484 4654 12486
rect 4710 12484 4734 12486
rect 4790 12484 4814 12486
rect 4574 12464 4870 12484
rect 5000 11762 5028 14440
rect 6472 13274 6500 14440
rect 6472 13246 6776 13274
rect 6384 13084 6680 13104
rect 6440 13082 6464 13084
rect 6520 13082 6544 13084
rect 6600 13082 6624 13084
rect 6462 13030 6464 13082
rect 6526 13030 6538 13082
rect 6600 13030 6602 13082
rect 6440 13028 6464 13030
rect 6520 13028 6544 13030
rect 6600 13028 6624 13030
rect 6384 13008 6680 13028
rect 6384 11996 6680 12016
rect 6440 11994 6464 11996
rect 6520 11994 6544 11996
rect 6600 11994 6624 11996
rect 6462 11942 6464 11994
rect 6526 11942 6538 11994
rect 6600 11942 6602 11994
rect 6440 11940 6464 11942
rect 6520 11940 6544 11942
rect 6600 11940 6624 11942
rect 6384 11920 6680 11940
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3252 8838 3280 9454
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3528 8945 3556 8978
rect 3514 8936 3570 8945
rect 3514 8871 3570 8880
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 2765 8732 3061 8752
rect 2821 8730 2845 8732
rect 2901 8730 2925 8732
rect 2981 8730 3005 8732
rect 2843 8678 2845 8730
rect 2907 8678 2919 8730
rect 2981 8678 2983 8730
rect 2821 8676 2845 8678
rect 2901 8676 2925 8678
rect 2981 8676 3005 8678
rect 2765 8656 3061 8676
rect 2412 8016 2464 8022
rect 2410 7984 2412 7993
rect 2464 7984 2466 7993
rect 2410 7919 2466 7928
rect 2765 7644 3061 7664
rect 2821 7642 2845 7644
rect 2901 7642 2925 7644
rect 2981 7642 3005 7644
rect 2843 7590 2845 7642
rect 2907 7590 2919 7642
rect 2981 7590 2983 7642
rect 2821 7588 2845 7590
rect 2901 7588 2925 7590
rect 2981 7588 3005 7590
rect 2765 7568 3061 7588
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2318 7440 2374 7449
rect 2318 7375 2374 7384
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 6934 1716 7278
rect 2332 7206 2360 7375
rect 2700 7342 2728 7482
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 3146 7304 3202 7313
rect 2780 7268 2832 7274
rect 3146 7239 3148 7248
rect 2780 7210 2832 7216
rect 3200 7239 3202 7248
rect 3148 7210 3200 7216
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2792 6934 2820 7210
rect 1676 6928 1728 6934
rect 1676 6870 1728 6876
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3160 6769 3188 6802
rect 3146 6760 3202 6769
rect 3146 6695 3202 6704
rect 2765 6556 3061 6576
rect 2821 6554 2845 6556
rect 2901 6554 2925 6556
rect 2981 6554 3005 6556
rect 2843 6502 2845 6554
rect 2907 6502 2919 6554
rect 2981 6502 2983 6554
rect 2821 6500 2845 6502
rect 2901 6500 2925 6502
rect 2981 6500 3005 6502
rect 2765 6480 3061 6500
rect 3252 6322 3280 8774
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 2765 5468 3061 5488
rect 2821 5466 2845 5468
rect 2901 5466 2925 5468
rect 2981 5466 3005 5468
rect 2843 5414 2845 5466
rect 2907 5414 2919 5466
rect 2981 5414 2983 5466
rect 2821 5412 2845 5414
rect 2901 5412 2925 5414
rect 2981 5412 3005 5414
rect 2765 5392 3061 5412
rect 3344 5030 3372 7822
rect 3436 6730 3464 8298
rect 3528 7886 3556 8871
rect 3620 7954 3648 9318
rect 3712 8022 3740 9318
rect 4172 9042 4200 11494
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 3790 8936 3846 8945
rect 3790 8871 3846 8880
rect 4068 8900 4120 8906
rect 3804 8634 3832 8871
rect 4068 8842 4120 8848
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3988 8430 4016 8774
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3884 7472 3936 7478
rect 3804 7420 3884 7426
rect 3804 7414 3936 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3700 7404 3752 7410
rect 3804 7398 3924 7414
rect 3804 7392 3832 7398
rect 3752 7364 3832 7392
rect 3700 7346 3752 7352
rect 3528 7274 3556 7346
rect 4080 7342 4108 8842
rect 4172 8498 4200 8978
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4172 7886 4200 8298
rect 4264 8090 4292 9454
rect 4356 8412 4384 11698
rect 4574 11452 4870 11472
rect 4630 11450 4654 11452
rect 4710 11450 4734 11452
rect 4790 11450 4814 11452
rect 4652 11398 4654 11450
rect 4716 11398 4728 11450
rect 4790 11398 4792 11450
rect 4630 11396 4654 11398
rect 4710 11396 4734 11398
rect 4790 11396 4814 11398
rect 4574 11376 4870 11396
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 4574 10364 4870 10384
rect 4630 10362 4654 10364
rect 4710 10362 4734 10364
rect 4790 10362 4814 10364
rect 4652 10310 4654 10362
rect 4716 10310 4728 10362
rect 4790 10310 4792 10362
rect 4630 10308 4654 10310
rect 4710 10308 4734 10310
rect 4790 10308 4814 10310
rect 4574 10288 4870 10308
rect 5368 10130 5396 11018
rect 6384 10908 6680 10928
rect 6440 10906 6464 10908
rect 6520 10906 6544 10908
rect 6600 10906 6624 10908
rect 6462 10854 6464 10906
rect 6526 10854 6538 10906
rect 6600 10854 6602 10906
rect 6440 10852 6464 10854
rect 6520 10852 6544 10854
rect 6600 10852 6624 10854
rect 6384 10832 6680 10852
rect 6748 10674 6776 13246
rect 7852 12782 7880 14440
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6932 10606 6960 12582
rect 8193 12540 8489 12560
rect 8249 12538 8273 12540
rect 8329 12538 8353 12540
rect 8409 12538 8433 12540
rect 8271 12486 8273 12538
rect 8335 12486 8347 12538
rect 8409 12486 8411 12538
rect 8249 12484 8273 12486
rect 8329 12484 8353 12486
rect 8409 12484 8433 12486
rect 8193 12464 8489 12484
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5172 10056 5224 10062
rect 5172 9998 5224 10004
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4574 9276 4870 9296
rect 4630 9274 4654 9276
rect 4710 9274 4734 9276
rect 4790 9274 4814 9276
rect 4652 9222 4654 9274
rect 4716 9222 4728 9274
rect 4790 9222 4792 9274
rect 4630 9220 4654 9222
rect 4710 9220 4734 9222
rect 4790 9220 4814 9222
rect 4574 9200 4870 9220
rect 4436 8424 4488 8430
rect 4356 8384 4436 8412
rect 4436 8366 4488 8372
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4356 8022 4384 8230
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3436 6610 3464 6666
rect 3436 6582 3556 6610
rect 3528 6254 3556 6582
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3528 5098 3556 6190
rect 3896 6186 3924 6802
rect 4172 6458 4200 7686
rect 4356 7410 4384 7686
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4252 6792 4304 6798
rect 4448 6780 4476 8366
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4574 8188 4870 8208
rect 4630 8186 4654 8188
rect 4710 8186 4734 8188
rect 4790 8186 4814 8188
rect 4652 8134 4654 8186
rect 4716 8134 4728 8186
rect 4790 8134 4792 8186
rect 4630 8132 4654 8134
rect 4710 8132 4734 8134
rect 4790 8132 4814 8134
rect 4574 8112 4870 8132
rect 4908 7342 4936 8230
rect 5092 8090 5120 9590
rect 5184 9586 5212 9998
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5184 7886 5212 9522
rect 5276 8974 5304 9522
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5276 7954 5304 8910
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5170 7440 5226 7449
rect 5170 7375 5226 7384
rect 5264 7404 5316 7410
rect 5184 7342 5212 7375
rect 5264 7346 5316 7352
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 4574 7100 4870 7120
rect 4630 7098 4654 7100
rect 4710 7098 4734 7100
rect 4790 7098 4814 7100
rect 4652 7046 4654 7098
rect 4716 7046 4728 7098
rect 4790 7046 4792 7098
rect 4630 7044 4654 7046
rect 4710 7044 4734 7046
rect 4790 7044 4814 7046
rect 4574 7024 4870 7044
rect 4908 6798 4936 7278
rect 5276 7177 5304 7346
rect 5262 7168 5318 7177
rect 5262 7103 5318 7112
rect 4304 6752 4476 6780
rect 4896 6792 4948 6798
rect 4252 6734 4304 6740
rect 4896 6734 4948 6740
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3974 6352 4030 6361
rect 3974 6287 4030 6296
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 3712 5574 3740 6122
rect 3988 5778 4016 6287
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3516 5092 3568 5098
rect 3516 5034 3568 5040
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 2765 4380 3061 4400
rect 2821 4378 2845 4380
rect 2901 4378 2925 4380
rect 2981 4378 3005 4380
rect 2843 4326 2845 4378
rect 2907 4326 2919 4378
rect 2981 4326 2983 4378
rect 2821 4324 2845 4326
rect 2901 4324 2925 4326
rect 2981 4324 3005 4326
rect 2765 4304 3061 4324
rect 664 3392 716 3398
rect 664 3334 716 3340
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 676 800 704 3334
rect 2056 800 2084 3334
rect 2765 3292 3061 3312
rect 2821 3290 2845 3292
rect 2901 3290 2925 3292
rect 2981 3290 3005 3292
rect 2843 3238 2845 3290
rect 2907 3238 2919 3290
rect 2981 3238 2983 3290
rect 2821 3236 2845 3238
rect 2901 3236 2925 3238
rect 2981 3236 3005 3238
rect 2765 3216 3061 3236
rect 2765 2204 3061 2224
rect 2821 2202 2845 2204
rect 2901 2202 2925 2204
rect 2981 2202 3005 2204
rect 2843 2150 2845 2202
rect 2907 2150 2919 2202
rect 2981 2150 2983 2202
rect 2821 2148 2845 2150
rect 2901 2148 2925 2150
rect 2981 2148 3005 2150
rect 2765 2128 3061 2148
rect 3528 800 3556 5034
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3620 1329 3648 4558
rect 3896 3777 3924 4966
rect 4080 4622 4108 6394
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 3882 3768 3938 3777
rect 3882 3703 3938 3712
rect 4264 3602 4292 6734
rect 4574 6012 4870 6032
rect 4630 6010 4654 6012
rect 4710 6010 4734 6012
rect 4790 6010 4814 6012
rect 4652 5958 4654 6010
rect 4716 5958 4728 6010
rect 4790 5958 4792 6010
rect 4630 5956 4654 5958
rect 4710 5956 4734 5958
rect 4790 5956 4814 5958
rect 4574 5936 4870 5956
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4448 3670 4476 5714
rect 4908 4978 4936 6734
rect 5000 6254 5028 6734
rect 5368 6338 5396 10066
rect 6196 10062 6224 10406
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9042 5488 9454
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5460 8566 5488 8978
rect 5552 8838 5580 9590
rect 5644 9110 5672 9862
rect 5632 9104 5684 9110
rect 5632 9046 5684 9052
rect 5722 9072 5778 9081
rect 5722 9007 5724 9016
rect 5776 9007 5778 9016
rect 5724 8978 5776 8984
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5552 7954 5580 8774
rect 5644 8498 5672 8910
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5460 6474 5488 6870
rect 5552 6662 5580 7346
rect 5632 7336 5684 7342
rect 5630 7304 5632 7313
rect 5684 7304 5686 7313
rect 5630 7239 5686 7248
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5460 6446 5580 6474
rect 5276 6310 5396 6338
rect 4988 6248 5040 6254
rect 5080 6248 5132 6254
rect 4988 6190 5040 6196
rect 5078 6216 5080 6225
rect 5132 6216 5134 6225
rect 5078 6151 5134 6160
rect 5276 5846 5304 6310
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5368 5914 5396 6190
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5460 5030 5488 5782
rect 5552 5098 5580 6446
rect 5630 6216 5686 6225
rect 5630 6151 5686 6160
rect 5644 5710 5672 6151
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5736 5166 5764 7142
rect 5828 6730 5856 8366
rect 6104 7585 6132 9862
rect 6196 9586 6224 9998
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6196 7868 6224 8298
rect 6288 7970 6316 10406
rect 6380 10130 6408 10542
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6384 9820 6680 9840
rect 6440 9818 6464 9820
rect 6520 9818 6544 9820
rect 6600 9818 6624 9820
rect 6462 9766 6464 9818
rect 6526 9766 6538 9818
rect 6600 9766 6602 9818
rect 6440 9764 6464 9766
rect 6520 9764 6544 9766
rect 6600 9764 6624 9766
rect 6384 9744 6680 9764
rect 6460 9512 6512 9518
rect 6458 9480 6460 9489
rect 6512 9480 6514 9489
rect 6458 9415 6514 9424
rect 6460 9036 6512 9042
rect 6748 9024 6776 10406
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6512 8996 6776 9024
rect 6460 8978 6512 8984
rect 6472 8945 6500 8978
rect 6458 8936 6514 8945
rect 6458 8871 6514 8880
rect 6384 8732 6680 8752
rect 6440 8730 6464 8732
rect 6520 8730 6544 8732
rect 6600 8730 6624 8732
rect 6462 8678 6464 8730
rect 6526 8678 6538 8730
rect 6600 8678 6602 8730
rect 6440 8676 6464 8678
rect 6520 8676 6544 8678
rect 6600 8676 6624 8678
rect 6384 8656 6680 8676
rect 6840 8242 6868 9998
rect 6932 9382 6960 10066
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6932 8974 6960 9046
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8362 6960 8910
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6840 8214 6960 8242
rect 6288 7954 6408 7970
rect 6288 7948 6420 7954
rect 6288 7942 6368 7948
rect 6368 7890 6420 7896
rect 6196 7840 6316 7868
rect 6090 7576 6146 7585
rect 6090 7511 6146 7520
rect 6000 7336 6052 7342
rect 5906 7304 5962 7313
rect 6000 7278 6052 7284
rect 5906 7239 5962 7248
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5828 6186 5856 6666
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 5828 5166 5856 5578
rect 5920 5302 5948 7239
rect 6012 7002 6040 7278
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6104 6934 6132 7511
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 6196 7177 6224 7210
rect 6182 7168 6238 7177
rect 6182 7103 6238 7112
rect 6288 7018 6316 7840
rect 6384 7644 6680 7664
rect 6440 7642 6464 7644
rect 6520 7642 6544 7644
rect 6600 7642 6624 7644
rect 6462 7590 6464 7642
rect 6526 7590 6538 7642
rect 6600 7590 6602 7642
rect 6440 7588 6464 7590
rect 6520 7588 6544 7590
rect 6600 7588 6624 7590
rect 6384 7568 6680 7588
rect 6736 7540 6788 7546
rect 6196 6990 6316 7018
rect 6656 7500 6736 7528
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5448 5024 5500 5030
rect 4986 4992 5042 5001
rect 4908 4950 4986 4978
rect 4574 4924 4870 4944
rect 5448 4966 5500 4972
rect 4986 4927 5042 4936
rect 4630 4922 4654 4924
rect 4710 4922 4734 4924
rect 4790 4922 4814 4924
rect 4652 4870 4654 4922
rect 4716 4870 4728 4922
rect 4790 4870 4792 4922
rect 4630 4868 4654 4870
rect 4710 4868 4734 4870
rect 4790 4868 4814 4870
rect 4574 4848 4870 4868
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4214 5580 4422
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 6012 4146 6040 6734
rect 6104 6322 6132 6734
rect 6196 6361 6224 6990
rect 6656 6866 6684 7500
rect 6736 7482 6788 7488
rect 6932 7426 6960 8214
rect 7024 7954 7052 9930
rect 7116 8974 7144 11698
rect 8193 11452 8489 11472
rect 8249 11450 8273 11452
rect 8329 11450 8353 11452
rect 8409 11450 8433 11452
rect 8271 11398 8273 11450
rect 8335 11398 8347 11450
rect 8409 11398 8411 11450
rect 8249 11396 8273 11398
rect 8329 11396 8353 11398
rect 8409 11396 8433 11398
rect 8193 11376 8489 11396
rect 8574 11384 8630 11393
rect 8574 11319 8630 11328
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7208 9110 7236 10542
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7300 9518 7328 10134
rect 7392 10010 7420 10474
rect 8193 10364 8489 10384
rect 8249 10362 8273 10364
rect 8329 10362 8353 10364
rect 8409 10362 8433 10364
rect 8271 10310 8273 10362
rect 8335 10310 8347 10362
rect 8409 10310 8411 10362
rect 8249 10308 8273 10310
rect 8329 10308 8353 10310
rect 8409 10308 8433 10310
rect 8193 10288 8489 10308
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 7932 10192 7984 10198
rect 7932 10134 7984 10140
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7656 10056 7708 10062
rect 7392 9982 7512 10010
rect 7656 9998 7708 10004
rect 7760 10010 7788 10066
rect 7484 9926 7512 9982
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7208 8838 7236 8910
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7208 8430 7236 8570
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 7116 7834 7144 8366
rect 7300 7954 7328 8774
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7116 7806 7236 7834
rect 7208 7585 7236 7806
rect 7194 7576 7250 7585
rect 7194 7511 7250 7520
rect 7196 7472 7248 7478
rect 6932 7398 7052 7426
rect 7196 7414 7248 7420
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6748 6934 6776 7278
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6826 7032 6882 7041
rect 6826 6967 6828 6976
rect 6880 6967 6882 6976
rect 6828 6938 6880 6944
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6472 6769 6500 6802
rect 6458 6760 6514 6769
rect 6458 6695 6514 6704
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6182 6352 6238 6361
rect 6092 6316 6144 6322
rect 6182 6287 6238 6296
rect 6092 6258 6144 6264
rect 6288 6254 6316 6598
rect 6384 6556 6680 6576
rect 6440 6554 6464 6556
rect 6520 6554 6544 6556
rect 6600 6554 6624 6556
rect 6462 6502 6464 6554
rect 6526 6502 6538 6554
rect 6600 6502 6602 6554
rect 6440 6500 6464 6502
rect 6520 6500 6544 6502
rect 6600 6500 6624 6502
rect 6384 6480 6680 6500
rect 6550 6352 6606 6361
rect 6550 6287 6606 6296
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6196 6089 6224 6190
rect 6182 6080 6238 6089
rect 6182 6015 6238 6024
rect 6366 5808 6422 5817
rect 6276 5772 6328 5778
rect 6366 5743 6422 5752
rect 6276 5714 6328 5720
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 4574 3836 4870 3856
rect 4630 3834 4654 3836
rect 4710 3834 4734 3836
rect 4790 3834 4814 3836
rect 4652 3782 4654 3834
rect 4716 3782 4728 3834
rect 4790 3782 4792 3834
rect 4630 3780 4654 3782
rect 4710 3780 4734 3782
rect 4790 3780 4814 3782
rect 4574 3760 4870 3780
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4574 2748 4870 2768
rect 4630 2746 4654 2748
rect 4710 2746 4734 2748
rect 4790 2746 4814 2748
rect 4652 2694 4654 2746
rect 4716 2694 4728 2746
rect 4790 2694 4792 2746
rect 4630 2692 4654 2694
rect 4710 2692 4734 2694
rect 4790 2692 4814 2694
rect 4574 2672 4870 2692
rect 3606 1320 3662 1329
rect 3606 1255 3662 1264
rect 5000 800 5028 4082
rect 6104 4010 6132 4490
rect 6196 4078 6224 5646
rect 6288 5273 6316 5714
rect 6380 5642 6408 5743
rect 6564 5710 6592 6287
rect 6748 6254 6776 6870
rect 6932 6746 6960 7210
rect 6840 6718 6960 6746
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6656 6089 6684 6190
rect 6642 6080 6698 6089
rect 6642 6015 6698 6024
rect 6840 5930 6868 6718
rect 7024 6338 7052 7398
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 6748 5902 6868 5930
rect 6932 6310 7052 6338
rect 6748 5778 6776 5902
rect 6932 5794 6960 6310
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6840 5766 6960 5794
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6734 5672 6790 5681
rect 6368 5636 6420 5642
rect 6734 5607 6790 5616
rect 6368 5578 6420 5584
rect 6384 5468 6680 5488
rect 6440 5466 6464 5468
rect 6520 5466 6544 5468
rect 6600 5466 6624 5468
rect 6462 5414 6464 5466
rect 6526 5414 6538 5466
rect 6600 5414 6602 5466
rect 6440 5412 6464 5414
rect 6520 5412 6544 5414
rect 6600 5412 6624 5414
rect 6384 5392 6680 5412
rect 6552 5296 6604 5302
rect 6274 5264 6330 5273
rect 6552 5238 6604 5244
rect 6274 5199 6330 5208
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4570 6408 5102
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4690 6500 4966
rect 6564 4690 6592 5238
rect 6748 5166 6776 5607
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6642 4720 6698 4729
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6552 4684 6604 4690
rect 6642 4655 6698 4664
rect 6552 4626 6604 4632
rect 6656 4622 6684 4655
rect 6288 4542 6408 4570
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6288 4282 6316 4542
rect 6384 4380 6680 4400
rect 6440 4378 6464 4380
rect 6520 4378 6544 4380
rect 6600 4378 6624 4380
rect 6462 4326 6464 4378
rect 6526 4326 6538 4378
rect 6600 4326 6602 4378
rect 6440 4324 6464 4326
rect 6520 4324 6544 4326
rect 6600 4324 6624 4326
rect 6384 4304 6680 4324
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6840 4214 6868 5766
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6932 5370 6960 5646
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6918 5264 6974 5273
rect 7024 5234 7052 6190
rect 7116 5370 7144 7278
rect 7208 5778 7236 7414
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7300 5846 7328 7278
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7196 5636 7248 5642
rect 7196 5578 7248 5584
rect 7104 5364 7156 5370
rect 7104 5306 7156 5312
rect 6918 5199 6974 5208
rect 7012 5228 7064 5234
rect 6932 5030 6960 5199
rect 7012 5170 7064 5176
rect 7208 5166 7236 5578
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 7102 4992 7158 5001
rect 7102 4927 7158 4936
rect 7116 4690 7144 4927
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7208 4282 7236 5102
rect 7300 4826 7328 5782
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7392 4622 7420 9658
rect 7484 9625 7512 9862
rect 7470 9616 7526 9625
rect 7470 9551 7526 9560
rect 7576 9042 7604 9862
rect 7668 9722 7696 9998
rect 7760 9982 7880 10010
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7654 9616 7710 9625
rect 7654 9551 7710 9560
rect 7668 9518 7696 9551
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7562 8936 7618 8945
rect 7562 8871 7618 8880
rect 7470 8256 7526 8265
rect 7470 8191 7526 8200
rect 7484 7562 7512 8191
rect 7576 7698 7604 8871
rect 7668 7818 7696 9454
rect 7760 8430 7788 9658
rect 7852 9081 7880 9982
rect 7944 9722 7972 10134
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 8036 9518 8064 10202
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8116 9512 8168 9518
rect 8220 9489 8248 9522
rect 8116 9454 8168 9460
rect 8206 9480 8262 9489
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 7838 9072 7894 9081
rect 7838 9007 7894 9016
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7852 8430 7880 8910
rect 7944 8809 7972 9386
rect 7930 8800 7986 8809
rect 7930 8735 7986 8744
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7930 8392 7986 8401
rect 7760 7954 7788 8366
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7748 7744 7800 7750
rect 7654 7712 7710 7721
rect 7576 7670 7654 7698
rect 7748 7686 7800 7692
rect 7654 7647 7710 7656
rect 7484 7534 7604 7562
rect 7576 6905 7604 7534
rect 7562 6896 7618 6905
rect 7472 6860 7524 6866
rect 7562 6831 7618 6840
rect 7472 6802 7524 6808
rect 7484 5817 7512 6802
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7470 5808 7526 5817
rect 7470 5743 7526 5752
rect 7484 5166 7512 5743
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7576 4758 7604 6734
rect 7668 6730 7696 7647
rect 7760 7290 7788 7686
rect 7852 7478 7880 8366
rect 7930 8327 7986 8336
rect 7944 8294 7972 8327
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 7857 7972 8230
rect 7930 7848 7986 7857
rect 7930 7783 7986 7792
rect 8036 7750 8064 9454
rect 8128 9110 8156 9454
rect 8206 9415 8262 9424
rect 8193 9276 8489 9296
rect 8249 9274 8273 9276
rect 8329 9274 8353 9276
rect 8409 9274 8433 9276
rect 8271 9222 8273 9274
rect 8335 9222 8347 9274
rect 8409 9222 8411 9274
rect 8249 9220 8273 9222
rect 8329 9220 8353 9222
rect 8409 9220 8433 9222
rect 8193 9200 8489 9220
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7840 7472 7892 7478
rect 7838 7440 7840 7449
rect 7892 7440 7894 7449
rect 8128 7426 8156 9046
rect 8588 9024 8616 11319
rect 9324 10810 9352 14440
rect 9586 13968 9642 13977
rect 9586 13903 9642 13912
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8496 8996 8616 9024
rect 8496 8401 8524 8996
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8482 8392 8538 8401
rect 8482 8327 8538 8336
rect 8193 8188 8489 8208
rect 8249 8186 8273 8188
rect 8329 8186 8353 8188
rect 8409 8186 8433 8188
rect 8271 8134 8273 8186
rect 8335 8134 8347 8186
rect 8409 8134 8411 8186
rect 8249 8132 8273 8134
rect 8329 8132 8353 8134
rect 8409 8132 8433 8134
rect 8193 8112 8489 8132
rect 8588 8090 8616 8842
rect 8680 8090 8708 10678
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8772 8906 8800 9998
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 8864 8498 8892 9318
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8956 8634 8984 8910
rect 9048 8634 9076 9454
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8392 8016 8444 8022
rect 8390 7984 8392 7993
rect 8444 7984 8446 7993
rect 8208 7948 8260 7954
rect 8390 7919 8446 7928
rect 8208 7890 8260 7896
rect 8220 7562 8248 7890
rect 8576 7880 8628 7886
rect 8312 7828 8576 7834
rect 8312 7822 8628 7828
rect 8312 7806 8616 7822
rect 8312 7750 8340 7806
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8574 7576 8630 7585
rect 8220 7534 8340 7562
rect 8128 7410 8248 7426
rect 8024 7404 8076 7410
rect 7838 7375 7894 7384
rect 7852 7349 7880 7375
rect 7944 7364 8024 7392
rect 7838 7304 7894 7313
rect 7760 7262 7838 7290
rect 7838 7239 7894 7248
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7654 6624 7710 6633
rect 7654 6559 7710 6568
rect 7668 6254 7696 6559
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 4808 7696 6054
rect 7760 5778 7788 6734
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7760 5642 7788 5714
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 7760 5001 7788 5238
rect 7746 4992 7802 5001
rect 7746 4927 7802 4936
rect 7748 4820 7800 4826
rect 7668 4780 7748 4808
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7196 4276 7248 4282
rect 7196 4218 7248 4224
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6840 4078 6868 4150
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6384 3292 6680 3312
rect 6440 3290 6464 3292
rect 6520 3290 6544 3292
rect 6600 3290 6624 3292
rect 6462 3238 6464 3290
rect 6526 3238 6538 3290
rect 6600 3238 6602 3290
rect 6440 3236 6464 3238
rect 6520 3236 6544 3238
rect 6600 3236 6624 3238
rect 6384 3216 6680 3236
rect 7668 2514 7696 4780
rect 7748 4762 7800 4768
rect 7852 4690 7880 7239
rect 7944 5710 7972 7364
rect 8128 7404 8260 7410
rect 8128 7398 8208 7404
rect 8024 7346 8076 7352
rect 8208 7346 8260 7352
rect 8312 7290 8340 7534
rect 8574 7511 8630 7520
rect 8036 7262 8340 7290
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8036 5574 8064 7262
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8128 6866 8156 7142
rect 8193 7100 8489 7120
rect 8249 7098 8273 7100
rect 8329 7098 8353 7100
rect 8409 7098 8433 7100
rect 8271 7046 8273 7098
rect 8335 7046 8347 7098
rect 8409 7046 8411 7098
rect 8249 7044 8273 7046
rect 8329 7044 8353 7046
rect 8409 7044 8433 7046
rect 8193 7024 8489 7044
rect 8588 6866 8616 7511
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8128 5778 8156 6802
rect 8193 6012 8489 6032
rect 8249 6010 8273 6012
rect 8329 6010 8353 6012
rect 8409 6010 8433 6012
rect 8271 5958 8273 6010
rect 8335 5958 8347 6010
rect 8409 5958 8411 6010
rect 8249 5956 8273 5958
rect 8329 5956 8353 5958
rect 8409 5956 8433 5958
rect 8193 5936 8489 5956
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8114 5672 8170 5681
rect 8114 5607 8116 5616
rect 8168 5607 8170 5616
rect 8116 5578 8168 5584
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8036 4729 8064 5034
rect 8193 4924 8489 4944
rect 8249 4922 8273 4924
rect 8329 4922 8353 4924
rect 8409 4922 8433 4924
rect 8271 4870 8273 4922
rect 8335 4870 8347 4922
rect 8409 4870 8411 4922
rect 8249 4868 8273 4870
rect 8329 4868 8353 4870
rect 8409 4868 8433 4870
rect 8193 4848 8489 4868
rect 8022 4720 8078 4729
rect 7840 4684 7892 4690
rect 8022 4655 8078 4664
rect 8392 4684 8444 4690
rect 7840 4626 7892 4632
rect 8392 4626 8444 4632
rect 8404 4554 8432 4626
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 7852 4010 7880 4490
rect 8588 4486 8616 5510
rect 8680 4554 8708 7686
rect 8772 7342 8800 8230
rect 8864 7410 8892 8434
rect 8956 8022 8984 8570
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 9048 7868 9076 8570
rect 9140 8566 9168 8978
rect 9128 8560 9180 8566
rect 9128 8502 9180 8508
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8956 7840 9076 7868
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8772 4622 8800 7278
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8864 5710 8892 6258
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8668 4548 8720 4554
rect 8668 4490 8720 4496
rect 8576 4480 8628 4486
rect 8576 4422 8628 4428
rect 8864 4078 8892 4626
rect 8956 4282 8984 7840
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9048 7410 9076 7482
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9140 7342 9168 8366
rect 9324 7750 9352 10746
rect 9600 9178 9628 13903
rect 10002 13084 10298 13104
rect 10058 13082 10082 13084
rect 10138 13082 10162 13084
rect 10218 13082 10242 13084
rect 10080 13030 10082 13082
rect 10144 13030 10156 13082
rect 10218 13030 10220 13082
rect 10058 13028 10082 13030
rect 10138 13028 10162 13030
rect 10218 13028 10242 13030
rect 10002 13008 10298 13028
rect 10002 11996 10298 12016
rect 10058 11994 10082 11996
rect 10138 11994 10162 11996
rect 10218 11994 10242 11996
rect 10080 11942 10082 11994
rect 10144 11942 10156 11994
rect 10218 11942 10220 11994
rect 10058 11940 10082 11942
rect 10138 11940 10162 11942
rect 10218 11940 10242 11942
rect 10002 11920 10298 11940
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10002 10908 10298 10928
rect 10058 10906 10082 10908
rect 10138 10906 10162 10908
rect 10218 10906 10242 10908
rect 10080 10854 10082 10906
rect 10144 10854 10156 10906
rect 10218 10854 10220 10906
rect 10058 10852 10082 10854
rect 10138 10852 10162 10854
rect 10218 10852 10242 10854
rect 10002 10832 10298 10852
rect 10002 9820 10298 9840
rect 10058 9818 10082 9820
rect 10138 9818 10162 9820
rect 10218 9818 10242 9820
rect 10080 9766 10082 9818
rect 10144 9766 10156 9818
rect 10218 9766 10220 9818
rect 10058 9764 10082 9766
rect 10138 9764 10162 9766
rect 10218 9764 10242 9766
rect 10002 9744 10298 9764
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9402 7848 9458 7857
rect 9402 7783 9458 7792
rect 9312 7744 9364 7750
rect 9218 7712 9274 7721
rect 9312 7686 9364 7692
rect 9218 7647 9274 7656
rect 9232 7562 9260 7647
rect 9232 7534 9352 7562
rect 9324 7478 9352 7534
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9048 6361 9076 6734
rect 9034 6352 9090 6361
rect 9034 6287 9090 6296
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 7852 2990 7880 3946
rect 8193 3836 8489 3856
rect 8249 3834 8273 3836
rect 8329 3834 8353 3836
rect 8409 3834 8433 3836
rect 8271 3782 8273 3834
rect 8335 3782 8347 3834
rect 8409 3782 8411 3834
rect 8249 3780 8273 3782
rect 8329 3780 8353 3782
rect 8409 3780 8433 3782
rect 8193 3760 8489 3780
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6384 2204 6680 2224
rect 6440 2202 6464 2204
rect 6520 2202 6544 2204
rect 6600 2202 6624 2204
rect 6462 2150 6464 2202
rect 6526 2150 6538 2202
rect 6600 2150 6602 2202
rect 6440 2148 6464 2150
rect 6520 2148 6544 2150
rect 6600 2148 6624 2150
rect 6384 2128 6680 2148
rect 6748 1170 6776 2246
rect 6472 1142 6776 1170
rect 6472 800 6500 1142
rect 7852 800 7880 2790
rect 8193 2748 8489 2768
rect 8249 2746 8273 2748
rect 8329 2746 8353 2748
rect 8409 2746 8433 2748
rect 8271 2694 8273 2746
rect 8335 2694 8347 2746
rect 8409 2694 8411 2746
rect 8249 2692 8273 2694
rect 8329 2692 8353 2694
rect 8409 2692 8433 2694
rect 8193 2672 8489 2692
rect 9048 1329 9076 5646
rect 9140 5234 9168 7278
rect 9232 7274 9260 7414
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9324 6662 9352 6870
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 5710 9260 6190
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9324 5030 9352 6598
rect 9416 5778 9444 7783
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9508 4758 9536 8230
rect 9600 7342 9628 8298
rect 9692 7834 9720 9590
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 7954 9812 8978
rect 9876 8090 9904 9522
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10002 8732 10298 8752
rect 10058 8730 10082 8732
rect 10138 8730 10162 8732
rect 10218 8730 10242 8732
rect 10080 8678 10082 8730
rect 10144 8678 10156 8730
rect 10218 8678 10220 8730
rect 10058 8676 10082 8678
rect 10138 8676 10162 8678
rect 10218 8676 10242 8678
rect 10002 8656 10298 8676
rect 10336 8634 10364 8842
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9968 8294 9996 8502
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9692 7806 9812 7834
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9692 7188 9720 7482
rect 9784 7324 9812 7806
rect 10002 7644 10298 7664
rect 10058 7642 10082 7644
rect 10138 7642 10162 7644
rect 10218 7642 10242 7644
rect 10080 7590 10082 7642
rect 10144 7590 10156 7642
rect 10218 7590 10220 7642
rect 10058 7588 10082 7590
rect 10138 7588 10162 7590
rect 10218 7588 10242 7590
rect 10002 7568 10298 7588
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 9956 7336 10008 7342
rect 9784 7296 9956 7324
rect 9956 7278 10008 7284
rect 9600 7160 9720 7188
rect 9600 6934 9628 7160
rect 9968 6934 9996 7278
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 10046 6896 10102 6905
rect 9968 6746 9996 6870
rect 10046 6831 10102 6840
rect 10060 6798 10088 6831
rect 9876 6718 9996 6746
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9680 6248 9732 6254
rect 9876 6225 9904 6718
rect 10336 6662 10364 7346
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10002 6556 10298 6576
rect 10058 6554 10082 6556
rect 10138 6554 10162 6556
rect 10218 6554 10242 6556
rect 10080 6502 10082 6554
rect 10144 6502 10156 6554
rect 10218 6502 10220 6554
rect 10058 6500 10082 6502
rect 10138 6500 10162 6502
rect 10218 6500 10242 6502
rect 10002 6480 10298 6500
rect 10428 6254 10456 9114
rect 10520 8430 10548 11018
rect 10796 9518 10824 14440
rect 12268 11082 12296 14440
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10690 8936 10746 8945
rect 10690 8871 10746 8880
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10416 6248 10468 6254
rect 9680 6190 9732 6196
rect 9862 6216 9918 6225
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9140 4146 9168 4626
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9034 1320 9090 1329
rect 9034 1255 9090 1264
rect 9324 800 9352 4694
rect 9600 3777 9628 6190
rect 9692 5778 9720 6190
rect 10416 6190 10468 6196
rect 9862 6151 9918 6160
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 10002 5468 10298 5488
rect 10058 5466 10082 5468
rect 10138 5466 10162 5468
rect 10218 5466 10242 5468
rect 10080 5414 10082 5466
rect 10144 5414 10156 5466
rect 10218 5414 10220 5466
rect 10058 5412 10082 5414
rect 10138 5412 10162 5414
rect 10218 5412 10242 5414
rect 10002 5392 10298 5412
rect 10520 4826 10548 8366
rect 10704 8090 10732 8871
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10612 7002 10640 7278
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10704 6882 10732 7890
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10784 7336 10836 7342
rect 10782 7304 10784 7313
rect 10836 7304 10838 7313
rect 10782 7239 10838 7248
rect 10612 6866 10732 6882
rect 10600 6860 10732 6866
rect 10652 6854 10732 6860
rect 10876 6860 10928 6866
rect 10600 6802 10652 6808
rect 10876 6802 10928 6808
rect 10612 5642 10640 6802
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6322 10824 6598
rect 10888 6458 10916 6802
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10888 6361 10916 6394
rect 10980 6390 11008 7686
rect 11164 7274 11192 7890
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 10968 6384 11020 6390
rect 10874 6352 10930 6361
rect 10784 6316 10836 6322
rect 10968 6326 11020 6332
rect 10874 6287 10930 6296
rect 10784 6258 10836 6264
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 11348 5098 11376 7278
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6934 11468 7142
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11336 5092 11388 5098
rect 11336 5034 11388 5040
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 10002 4380 10298 4400
rect 10058 4378 10082 4380
rect 10138 4378 10162 4380
rect 10218 4378 10242 4380
rect 10080 4326 10082 4378
rect 10144 4326 10156 4378
rect 10218 4326 10220 4378
rect 10058 4324 10082 4326
rect 10138 4324 10162 4326
rect 10218 4324 10242 4326
rect 10002 4304 10298 4324
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 9586 3768 9642 3777
rect 9586 3703 9642 3712
rect 10002 3292 10298 3312
rect 10058 3290 10082 3292
rect 10138 3290 10162 3292
rect 10218 3290 10242 3292
rect 10080 3238 10082 3290
rect 10144 3238 10156 3290
rect 10218 3238 10220 3290
rect 10058 3236 10082 3238
rect 10138 3236 10162 3238
rect 10218 3236 10242 3238
rect 10002 3216 10298 3236
rect 10002 2204 10298 2224
rect 10058 2202 10082 2204
rect 10138 2202 10162 2204
rect 10218 2202 10242 2204
rect 10080 2150 10082 2202
rect 10144 2150 10156 2202
rect 10218 2150 10220 2202
rect 10058 2148 10082 2150
rect 10138 2148 10162 2150
rect 10218 2148 10242 2150
rect 10002 2128 10298 2148
rect 10796 800 10824 3946
rect 12268 800 12296 4490
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4986 0 5042 800
rect 6458 0 6514 800
rect 7838 0 7894 800
rect 9310 0 9366 800
rect 10782 0 10838 800
rect 12254 0 12310 800
<< via2 >>
rect 3422 13912 3478 13968
rect 2765 13082 2821 13084
rect 2845 13082 2901 13084
rect 2925 13082 2981 13084
rect 3005 13082 3061 13084
rect 2765 13030 2791 13082
rect 2791 13030 2821 13082
rect 2845 13030 2855 13082
rect 2855 13030 2901 13082
rect 2925 13030 2971 13082
rect 2971 13030 2981 13082
rect 3005 13030 3035 13082
rect 3035 13030 3061 13082
rect 2765 13028 2821 13030
rect 2845 13028 2901 13030
rect 2925 13028 2981 13030
rect 3005 13028 3061 13030
rect 2765 11994 2821 11996
rect 2845 11994 2901 11996
rect 2925 11994 2981 11996
rect 3005 11994 3061 11996
rect 2765 11942 2791 11994
rect 2791 11942 2821 11994
rect 2845 11942 2855 11994
rect 2855 11942 2901 11994
rect 2925 11942 2971 11994
rect 2971 11942 2981 11994
rect 3005 11942 3035 11994
rect 3035 11942 3061 11994
rect 2765 11940 2821 11942
rect 2845 11940 2901 11942
rect 2925 11940 2981 11942
rect 3005 11940 3061 11942
rect 1950 11328 2006 11384
rect 2765 10906 2821 10908
rect 2845 10906 2901 10908
rect 2925 10906 2981 10908
rect 3005 10906 3061 10908
rect 2765 10854 2791 10906
rect 2791 10854 2821 10906
rect 2845 10854 2855 10906
rect 2855 10854 2901 10906
rect 2925 10854 2971 10906
rect 2971 10854 2981 10906
rect 3005 10854 3035 10906
rect 3035 10854 3061 10906
rect 2765 10852 2821 10854
rect 2845 10852 2901 10854
rect 2925 10852 2981 10854
rect 3005 10852 3061 10854
rect 2765 9818 2821 9820
rect 2845 9818 2901 9820
rect 2925 9818 2981 9820
rect 3005 9818 3061 9820
rect 2765 9766 2791 9818
rect 2791 9766 2821 9818
rect 2845 9766 2855 9818
rect 2855 9766 2901 9818
rect 2925 9766 2971 9818
rect 2971 9766 2981 9818
rect 3005 9766 3035 9818
rect 3035 9766 3061 9818
rect 2765 9764 2821 9766
rect 2845 9764 2901 9766
rect 2925 9764 2981 9766
rect 3005 9764 3061 9766
rect 4574 12538 4630 12540
rect 4654 12538 4710 12540
rect 4734 12538 4790 12540
rect 4814 12538 4870 12540
rect 4574 12486 4600 12538
rect 4600 12486 4630 12538
rect 4654 12486 4664 12538
rect 4664 12486 4710 12538
rect 4734 12486 4780 12538
rect 4780 12486 4790 12538
rect 4814 12486 4844 12538
rect 4844 12486 4870 12538
rect 4574 12484 4630 12486
rect 4654 12484 4710 12486
rect 4734 12484 4790 12486
rect 4814 12484 4870 12486
rect 6384 13082 6440 13084
rect 6464 13082 6520 13084
rect 6544 13082 6600 13084
rect 6624 13082 6680 13084
rect 6384 13030 6410 13082
rect 6410 13030 6440 13082
rect 6464 13030 6474 13082
rect 6474 13030 6520 13082
rect 6544 13030 6590 13082
rect 6590 13030 6600 13082
rect 6624 13030 6654 13082
rect 6654 13030 6680 13082
rect 6384 13028 6440 13030
rect 6464 13028 6520 13030
rect 6544 13028 6600 13030
rect 6624 13028 6680 13030
rect 6384 11994 6440 11996
rect 6464 11994 6520 11996
rect 6544 11994 6600 11996
rect 6624 11994 6680 11996
rect 6384 11942 6410 11994
rect 6410 11942 6440 11994
rect 6464 11942 6474 11994
rect 6474 11942 6520 11994
rect 6544 11942 6590 11994
rect 6590 11942 6600 11994
rect 6624 11942 6654 11994
rect 6654 11942 6680 11994
rect 6384 11940 6440 11942
rect 6464 11940 6520 11942
rect 6544 11940 6600 11942
rect 6624 11940 6680 11942
rect 3514 8880 3570 8936
rect 2765 8730 2821 8732
rect 2845 8730 2901 8732
rect 2925 8730 2981 8732
rect 3005 8730 3061 8732
rect 2765 8678 2791 8730
rect 2791 8678 2821 8730
rect 2845 8678 2855 8730
rect 2855 8678 2901 8730
rect 2925 8678 2971 8730
rect 2971 8678 2981 8730
rect 3005 8678 3035 8730
rect 3035 8678 3061 8730
rect 2765 8676 2821 8678
rect 2845 8676 2901 8678
rect 2925 8676 2981 8678
rect 3005 8676 3061 8678
rect 2410 7964 2412 7984
rect 2412 7964 2464 7984
rect 2464 7964 2466 7984
rect 2410 7928 2466 7964
rect 2765 7642 2821 7644
rect 2845 7642 2901 7644
rect 2925 7642 2981 7644
rect 3005 7642 3061 7644
rect 2765 7590 2791 7642
rect 2791 7590 2821 7642
rect 2845 7590 2855 7642
rect 2855 7590 2901 7642
rect 2925 7590 2971 7642
rect 2971 7590 2981 7642
rect 3005 7590 3035 7642
rect 3035 7590 3061 7642
rect 2765 7588 2821 7590
rect 2845 7588 2901 7590
rect 2925 7588 2981 7590
rect 3005 7588 3061 7590
rect 2318 7384 2374 7440
rect 3146 7268 3202 7304
rect 3146 7248 3148 7268
rect 3148 7248 3200 7268
rect 3200 7248 3202 7268
rect 3146 6704 3202 6760
rect 2765 6554 2821 6556
rect 2845 6554 2901 6556
rect 2925 6554 2981 6556
rect 3005 6554 3061 6556
rect 2765 6502 2791 6554
rect 2791 6502 2821 6554
rect 2845 6502 2855 6554
rect 2855 6502 2901 6554
rect 2925 6502 2971 6554
rect 2971 6502 2981 6554
rect 3005 6502 3035 6554
rect 3035 6502 3061 6554
rect 2765 6500 2821 6502
rect 2845 6500 2901 6502
rect 2925 6500 2981 6502
rect 3005 6500 3061 6502
rect 2765 5466 2821 5468
rect 2845 5466 2901 5468
rect 2925 5466 2981 5468
rect 3005 5466 3061 5468
rect 2765 5414 2791 5466
rect 2791 5414 2821 5466
rect 2845 5414 2855 5466
rect 2855 5414 2901 5466
rect 2925 5414 2971 5466
rect 2971 5414 2981 5466
rect 3005 5414 3035 5466
rect 3035 5414 3061 5466
rect 2765 5412 2821 5414
rect 2845 5412 2901 5414
rect 2925 5412 2981 5414
rect 3005 5412 3061 5414
rect 3790 8880 3846 8936
rect 4574 11450 4630 11452
rect 4654 11450 4710 11452
rect 4734 11450 4790 11452
rect 4814 11450 4870 11452
rect 4574 11398 4600 11450
rect 4600 11398 4630 11450
rect 4654 11398 4664 11450
rect 4664 11398 4710 11450
rect 4734 11398 4780 11450
rect 4780 11398 4790 11450
rect 4814 11398 4844 11450
rect 4844 11398 4870 11450
rect 4574 11396 4630 11398
rect 4654 11396 4710 11398
rect 4734 11396 4790 11398
rect 4814 11396 4870 11398
rect 4574 10362 4630 10364
rect 4654 10362 4710 10364
rect 4734 10362 4790 10364
rect 4814 10362 4870 10364
rect 4574 10310 4600 10362
rect 4600 10310 4630 10362
rect 4654 10310 4664 10362
rect 4664 10310 4710 10362
rect 4734 10310 4780 10362
rect 4780 10310 4790 10362
rect 4814 10310 4844 10362
rect 4844 10310 4870 10362
rect 4574 10308 4630 10310
rect 4654 10308 4710 10310
rect 4734 10308 4790 10310
rect 4814 10308 4870 10310
rect 6384 10906 6440 10908
rect 6464 10906 6520 10908
rect 6544 10906 6600 10908
rect 6624 10906 6680 10908
rect 6384 10854 6410 10906
rect 6410 10854 6440 10906
rect 6464 10854 6474 10906
rect 6474 10854 6520 10906
rect 6544 10854 6590 10906
rect 6590 10854 6600 10906
rect 6624 10854 6654 10906
rect 6654 10854 6680 10906
rect 6384 10852 6440 10854
rect 6464 10852 6520 10854
rect 6544 10852 6600 10854
rect 6624 10852 6680 10854
rect 8193 12538 8249 12540
rect 8273 12538 8329 12540
rect 8353 12538 8409 12540
rect 8433 12538 8489 12540
rect 8193 12486 8219 12538
rect 8219 12486 8249 12538
rect 8273 12486 8283 12538
rect 8283 12486 8329 12538
rect 8353 12486 8399 12538
rect 8399 12486 8409 12538
rect 8433 12486 8463 12538
rect 8463 12486 8489 12538
rect 8193 12484 8249 12486
rect 8273 12484 8329 12486
rect 8353 12484 8409 12486
rect 8433 12484 8489 12486
rect 4574 9274 4630 9276
rect 4654 9274 4710 9276
rect 4734 9274 4790 9276
rect 4814 9274 4870 9276
rect 4574 9222 4600 9274
rect 4600 9222 4630 9274
rect 4654 9222 4664 9274
rect 4664 9222 4710 9274
rect 4734 9222 4780 9274
rect 4780 9222 4790 9274
rect 4814 9222 4844 9274
rect 4844 9222 4870 9274
rect 4574 9220 4630 9222
rect 4654 9220 4710 9222
rect 4734 9220 4790 9222
rect 4814 9220 4870 9222
rect 4574 8186 4630 8188
rect 4654 8186 4710 8188
rect 4734 8186 4790 8188
rect 4814 8186 4870 8188
rect 4574 8134 4600 8186
rect 4600 8134 4630 8186
rect 4654 8134 4664 8186
rect 4664 8134 4710 8186
rect 4734 8134 4780 8186
rect 4780 8134 4790 8186
rect 4814 8134 4844 8186
rect 4844 8134 4870 8186
rect 4574 8132 4630 8134
rect 4654 8132 4710 8134
rect 4734 8132 4790 8134
rect 4814 8132 4870 8134
rect 5170 7384 5226 7440
rect 4574 7098 4630 7100
rect 4654 7098 4710 7100
rect 4734 7098 4790 7100
rect 4814 7098 4870 7100
rect 4574 7046 4600 7098
rect 4600 7046 4630 7098
rect 4654 7046 4664 7098
rect 4664 7046 4710 7098
rect 4734 7046 4780 7098
rect 4780 7046 4790 7098
rect 4814 7046 4844 7098
rect 4844 7046 4870 7098
rect 4574 7044 4630 7046
rect 4654 7044 4710 7046
rect 4734 7044 4790 7046
rect 4814 7044 4870 7046
rect 5262 7112 5318 7168
rect 3974 6296 4030 6352
rect 2765 4378 2821 4380
rect 2845 4378 2901 4380
rect 2925 4378 2981 4380
rect 3005 4378 3061 4380
rect 2765 4326 2791 4378
rect 2791 4326 2821 4378
rect 2845 4326 2855 4378
rect 2855 4326 2901 4378
rect 2925 4326 2971 4378
rect 2971 4326 2981 4378
rect 3005 4326 3035 4378
rect 3035 4326 3061 4378
rect 2765 4324 2821 4326
rect 2845 4324 2901 4326
rect 2925 4324 2981 4326
rect 3005 4324 3061 4326
rect 2765 3290 2821 3292
rect 2845 3290 2901 3292
rect 2925 3290 2981 3292
rect 3005 3290 3061 3292
rect 2765 3238 2791 3290
rect 2791 3238 2821 3290
rect 2845 3238 2855 3290
rect 2855 3238 2901 3290
rect 2925 3238 2971 3290
rect 2971 3238 2981 3290
rect 3005 3238 3035 3290
rect 3035 3238 3061 3290
rect 2765 3236 2821 3238
rect 2845 3236 2901 3238
rect 2925 3236 2981 3238
rect 3005 3236 3061 3238
rect 2765 2202 2821 2204
rect 2845 2202 2901 2204
rect 2925 2202 2981 2204
rect 3005 2202 3061 2204
rect 2765 2150 2791 2202
rect 2791 2150 2821 2202
rect 2845 2150 2855 2202
rect 2855 2150 2901 2202
rect 2925 2150 2971 2202
rect 2971 2150 2981 2202
rect 3005 2150 3035 2202
rect 3035 2150 3061 2202
rect 2765 2148 2821 2150
rect 2845 2148 2901 2150
rect 2925 2148 2981 2150
rect 3005 2148 3061 2150
rect 3882 3712 3938 3768
rect 4574 6010 4630 6012
rect 4654 6010 4710 6012
rect 4734 6010 4790 6012
rect 4814 6010 4870 6012
rect 4574 5958 4600 6010
rect 4600 5958 4630 6010
rect 4654 5958 4664 6010
rect 4664 5958 4710 6010
rect 4734 5958 4780 6010
rect 4780 5958 4790 6010
rect 4814 5958 4844 6010
rect 4844 5958 4870 6010
rect 4574 5956 4630 5958
rect 4654 5956 4710 5958
rect 4734 5956 4790 5958
rect 4814 5956 4870 5958
rect 5722 9036 5778 9072
rect 5722 9016 5724 9036
rect 5724 9016 5776 9036
rect 5776 9016 5778 9036
rect 5630 7284 5632 7304
rect 5632 7284 5684 7304
rect 5684 7284 5686 7304
rect 5630 7248 5686 7284
rect 5078 6196 5080 6216
rect 5080 6196 5132 6216
rect 5132 6196 5134 6216
rect 5078 6160 5134 6196
rect 5630 6160 5686 6216
rect 6384 9818 6440 9820
rect 6464 9818 6520 9820
rect 6544 9818 6600 9820
rect 6624 9818 6680 9820
rect 6384 9766 6410 9818
rect 6410 9766 6440 9818
rect 6464 9766 6474 9818
rect 6474 9766 6520 9818
rect 6544 9766 6590 9818
rect 6590 9766 6600 9818
rect 6624 9766 6654 9818
rect 6654 9766 6680 9818
rect 6384 9764 6440 9766
rect 6464 9764 6520 9766
rect 6544 9764 6600 9766
rect 6624 9764 6680 9766
rect 6458 9460 6460 9480
rect 6460 9460 6512 9480
rect 6512 9460 6514 9480
rect 6458 9424 6514 9460
rect 6458 8880 6514 8936
rect 6384 8730 6440 8732
rect 6464 8730 6520 8732
rect 6544 8730 6600 8732
rect 6624 8730 6680 8732
rect 6384 8678 6410 8730
rect 6410 8678 6440 8730
rect 6464 8678 6474 8730
rect 6474 8678 6520 8730
rect 6544 8678 6590 8730
rect 6590 8678 6600 8730
rect 6624 8678 6654 8730
rect 6654 8678 6680 8730
rect 6384 8676 6440 8678
rect 6464 8676 6520 8678
rect 6544 8676 6600 8678
rect 6624 8676 6680 8678
rect 6090 7520 6146 7576
rect 5906 7248 5962 7304
rect 6182 7112 6238 7168
rect 6384 7642 6440 7644
rect 6464 7642 6520 7644
rect 6544 7642 6600 7644
rect 6624 7642 6680 7644
rect 6384 7590 6410 7642
rect 6410 7590 6440 7642
rect 6464 7590 6474 7642
rect 6474 7590 6520 7642
rect 6544 7590 6590 7642
rect 6590 7590 6600 7642
rect 6624 7590 6654 7642
rect 6654 7590 6680 7642
rect 6384 7588 6440 7590
rect 6464 7588 6520 7590
rect 6544 7588 6600 7590
rect 6624 7588 6680 7590
rect 4986 4936 5042 4992
rect 4574 4922 4630 4924
rect 4654 4922 4710 4924
rect 4734 4922 4790 4924
rect 4814 4922 4870 4924
rect 4574 4870 4600 4922
rect 4600 4870 4630 4922
rect 4654 4870 4664 4922
rect 4664 4870 4710 4922
rect 4734 4870 4780 4922
rect 4780 4870 4790 4922
rect 4814 4870 4844 4922
rect 4844 4870 4870 4922
rect 4574 4868 4630 4870
rect 4654 4868 4710 4870
rect 4734 4868 4790 4870
rect 4814 4868 4870 4870
rect 8193 11450 8249 11452
rect 8273 11450 8329 11452
rect 8353 11450 8409 11452
rect 8433 11450 8489 11452
rect 8193 11398 8219 11450
rect 8219 11398 8249 11450
rect 8273 11398 8283 11450
rect 8283 11398 8329 11450
rect 8353 11398 8399 11450
rect 8399 11398 8409 11450
rect 8433 11398 8463 11450
rect 8463 11398 8489 11450
rect 8193 11396 8249 11398
rect 8273 11396 8329 11398
rect 8353 11396 8409 11398
rect 8433 11396 8489 11398
rect 8574 11328 8630 11384
rect 8193 10362 8249 10364
rect 8273 10362 8329 10364
rect 8353 10362 8409 10364
rect 8433 10362 8489 10364
rect 8193 10310 8219 10362
rect 8219 10310 8249 10362
rect 8273 10310 8283 10362
rect 8283 10310 8329 10362
rect 8353 10310 8399 10362
rect 8399 10310 8409 10362
rect 8433 10310 8463 10362
rect 8463 10310 8489 10362
rect 8193 10308 8249 10310
rect 8273 10308 8329 10310
rect 8353 10308 8409 10310
rect 8433 10308 8489 10310
rect 7194 7520 7250 7576
rect 6826 6996 6882 7032
rect 6826 6976 6828 6996
rect 6828 6976 6880 6996
rect 6880 6976 6882 6996
rect 6458 6704 6514 6760
rect 6182 6296 6238 6352
rect 6384 6554 6440 6556
rect 6464 6554 6520 6556
rect 6544 6554 6600 6556
rect 6624 6554 6680 6556
rect 6384 6502 6410 6554
rect 6410 6502 6440 6554
rect 6464 6502 6474 6554
rect 6474 6502 6520 6554
rect 6544 6502 6590 6554
rect 6590 6502 6600 6554
rect 6624 6502 6654 6554
rect 6654 6502 6680 6554
rect 6384 6500 6440 6502
rect 6464 6500 6520 6502
rect 6544 6500 6600 6502
rect 6624 6500 6680 6502
rect 6550 6296 6606 6352
rect 6182 6024 6238 6080
rect 6366 5752 6422 5808
rect 4574 3834 4630 3836
rect 4654 3834 4710 3836
rect 4734 3834 4790 3836
rect 4814 3834 4870 3836
rect 4574 3782 4600 3834
rect 4600 3782 4630 3834
rect 4654 3782 4664 3834
rect 4664 3782 4710 3834
rect 4734 3782 4780 3834
rect 4780 3782 4790 3834
rect 4814 3782 4844 3834
rect 4844 3782 4870 3834
rect 4574 3780 4630 3782
rect 4654 3780 4710 3782
rect 4734 3780 4790 3782
rect 4814 3780 4870 3782
rect 4574 2746 4630 2748
rect 4654 2746 4710 2748
rect 4734 2746 4790 2748
rect 4814 2746 4870 2748
rect 4574 2694 4600 2746
rect 4600 2694 4630 2746
rect 4654 2694 4664 2746
rect 4664 2694 4710 2746
rect 4734 2694 4780 2746
rect 4780 2694 4790 2746
rect 4814 2694 4844 2746
rect 4844 2694 4870 2746
rect 4574 2692 4630 2694
rect 4654 2692 4710 2694
rect 4734 2692 4790 2694
rect 4814 2692 4870 2694
rect 3606 1264 3662 1320
rect 6642 6024 6698 6080
rect 6734 5616 6790 5672
rect 6384 5466 6440 5468
rect 6464 5466 6520 5468
rect 6544 5466 6600 5468
rect 6624 5466 6680 5468
rect 6384 5414 6410 5466
rect 6410 5414 6440 5466
rect 6464 5414 6474 5466
rect 6474 5414 6520 5466
rect 6544 5414 6590 5466
rect 6590 5414 6600 5466
rect 6624 5414 6654 5466
rect 6654 5414 6680 5466
rect 6384 5412 6440 5414
rect 6464 5412 6520 5414
rect 6544 5412 6600 5414
rect 6624 5412 6680 5414
rect 6274 5208 6330 5264
rect 6642 4664 6698 4720
rect 6384 4378 6440 4380
rect 6464 4378 6520 4380
rect 6544 4378 6600 4380
rect 6624 4378 6680 4380
rect 6384 4326 6410 4378
rect 6410 4326 6440 4378
rect 6464 4326 6474 4378
rect 6474 4326 6520 4378
rect 6544 4326 6590 4378
rect 6590 4326 6600 4378
rect 6624 4326 6654 4378
rect 6654 4326 6680 4378
rect 6384 4324 6440 4326
rect 6464 4324 6520 4326
rect 6544 4324 6600 4326
rect 6624 4324 6680 4326
rect 6918 5208 6974 5264
rect 7102 4936 7158 4992
rect 7470 9560 7526 9616
rect 7654 9560 7710 9616
rect 7562 8880 7618 8936
rect 7470 8200 7526 8256
rect 7838 9016 7894 9072
rect 7930 8744 7986 8800
rect 7654 7656 7710 7712
rect 7562 6840 7618 6896
rect 7470 5752 7526 5808
rect 7930 8336 7986 8392
rect 7930 7792 7986 7848
rect 8206 9424 8262 9480
rect 8193 9274 8249 9276
rect 8273 9274 8329 9276
rect 8353 9274 8409 9276
rect 8433 9274 8489 9276
rect 8193 9222 8219 9274
rect 8219 9222 8249 9274
rect 8273 9222 8283 9274
rect 8283 9222 8329 9274
rect 8353 9222 8399 9274
rect 8399 9222 8409 9274
rect 8433 9222 8463 9274
rect 8463 9222 8489 9274
rect 8193 9220 8249 9222
rect 8273 9220 8329 9222
rect 8353 9220 8409 9222
rect 8433 9220 8489 9222
rect 7838 7420 7840 7440
rect 7840 7420 7892 7440
rect 7892 7420 7894 7440
rect 7838 7384 7894 7420
rect 9586 13912 9642 13968
rect 8482 8336 8538 8392
rect 8193 8186 8249 8188
rect 8273 8186 8329 8188
rect 8353 8186 8409 8188
rect 8433 8186 8489 8188
rect 8193 8134 8219 8186
rect 8219 8134 8249 8186
rect 8273 8134 8283 8186
rect 8283 8134 8329 8186
rect 8353 8134 8399 8186
rect 8399 8134 8409 8186
rect 8433 8134 8463 8186
rect 8463 8134 8489 8186
rect 8193 8132 8249 8134
rect 8273 8132 8329 8134
rect 8353 8132 8409 8134
rect 8433 8132 8489 8134
rect 8390 7964 8392 7984
rect 8392 7964 8444 7984
rect 8444 7964 8446 7984
rect 8390 7928 8446 7964
rect 7838 7248 7894 7304
rect 7654 6568 7710 6624
rect 7746 4936 7802 4992
rect 6384 3290 6440 3292
rect 6464 3290 6520 3292
rect 6544 3290 6600 3292
rect 6624 3290 6680 3292
rect 6384 3238 6410 3290
rect 6410 3238 6440 3290
rect 6464 3238 6474 3290
rect 6474 3238 6520 3290
rect 6544 3238 6590 3290
rect 6590 3238 6600 3290
rect 6624 3238 6654 3290
rect 6654 3238 6680 3290
rect 6384 3236 6440 3238
rect 6464 3236 6520 3238
rect 6544 3236 6600 3238
rect 6624 3236 6680 3238
rect 8574 7520 8630 7576
rect 8193 7098 8249 7100
rect 8273 7098 8329 7100
rect 8353 7098 8409 7100
rect 8433 7098 8489 7100
rect 8193 7046 8219 7098
rect 8219 7046 8249 7098
rect 8273 7046 8283 7098
rect 8283 7046 8329 7098
rect 8353 7046 8399 7098
rect 8399 7046 8409 7098
rect 8433 7046 8463 7098
rect 8463 7046 8489 7098
rect 8193 7044 8249 7046
rect 8273 7044 8329 7046
rect 8353 7044 8409 7046
rect 8433 7044 8489 7046
rect 8193 6010 8249 6012
rect 8273 6010 8329 6012
rect 8353 6010 8409 6012
rect 8433 6010 8489 6012
rect 8193 5958 8219 6010
rect 8219 5958 8249 6010
rect 8273 5958 8283 6010
rect 8283 5958 8329 6010
rect 8353 5958 8399 6010
rect 8399 5958 8409 6010
rect 8433 5958 8463 6010
rect 8463 5958 8489 6010
rect 8193 5956 8249 5958
rect 8273 5956 8329 5958
rect 8353 5956 8409 5958
rect 8433 5956 8489 5958
rect 8114 5636 8170 5672
rect 8114 5616 8116 5636
rect 8116 5616 8168 5636
rect 8168 5616 8170 5636
rect 8193 4922 8249 4924
rect 8273 4922 8329 4924
rect 8353 4922 8409 4924
rect 8433 4922 8489 4924
rect 8193 4870 8219 4922
rect 8219 4870 8249 4922
rect 8273 4870 8283 4922
rect 8283 4870 8329 4922
rect 8353 4870 8399 4922
rect 8399 4870 8409 4922
rect 8433 4870 8463 4922
rect 8463 4870 8489 4922
rect 8193 4868 8249 4870
rect 8273 4868 8329 4870
rect 8353 4868 8409 4870
rect 8433 4868 8489 4870
rect 8022 4664 8078 4720
rect 10002 13082 10058 13084
rect 10082 13082 10138 13084
rect 10162 13082 10218 13084
rect 10242 13082 10298 13084
rect 10002 13030 10028 13082
rect 10028 13030 10058 13082
rect 10082 13030 10092 13082
rect 10092 13030 10138 13082
rect 10162 13030 10208 13082
rect 10208 13030 10218 13082
rect 10242 13030 10272 13082
rect 10272 13030 10298 13082
rect 10002 13028 10058 13030
rect 10082 13028 10138 13030
rect 10162 13028 10218 13030
rect 10242 13028 10298 13030
rect 10002 11994 10058 11996
rect 10082 11994 10138 11996
rect 10162 11994 10218 11996
rect 10242 11994 10298 11996
rect 10002 11942 10028 11994
rect 10028 11942 10058 11994
rect 10082 11942 10092 11994
rect 10092 11942 10138 11994
rect 10162 11942 10208 11994
rect 10208 11942 10218 11994
rect 10242 11942 10272 11994
rect 10272 11942 10298 11994
rect 10002 11940 10058 11942
rect 10082 11940 10138 11942
rect 10162 11940 10218 11942
rect 10242 11940 10298 11942
rect 10002 10906 10058 10908
rect 10082 10906 10138 10908
rect 10162 10906 10218 10908
rect 10242 10906 10298 10908
rect 10002 10854 10028 10906
rect 10028 10854 10058 10906
rect 10082 10854 10092 10906
rect 10092 10854 10138 10906
rect 10162 10854 10208 10906
rect 10208 10854 10218 10906
rect 10242 10854 10272 10906
rect 10272 10854 10298 10906
rect 10002 10852 10058 10854
rect 10082 10852 10138 10854
rect 10162 10852 10218 10854
rect 10242 10852 10298 10854
rect 10002 9818 10058 9820
rect 10082 9818 10138 9820
rect 10162 9818 10218 9820
rect 10242 9818 10298 9820
rect 10002 9766 10028 9818
rect 10028 9766 10058 9818
rect 10082 9766 10092 9818
rect 10092 9766 10138 9818
rect 10162 9766 10208 9818
rect 10208 9766 10218 9818
rect 10242 9766 10272 9818
rect 10272 9766 10298 9818
rect 10002 9764 10058 9766
rect 10082 9764 10138 9766
rect 10162 9764 10218 9766
rect 10242 9764 10298 9766
rect 9402 7792 9458 7848
rect 9218 7656 9274 7712
rect 9034 6296 9090 6352
rect 8193 3834 8249 3836
rect 8273 3834 8329 3836
rect 8353 3834 8409 3836
rect 8433 3834 8489 3836
rect 8193 3782 8219 3834
rect 8219 3782 8249 3834
rect 8273 3782 8283 3834
rect 8283 3782 8329 3834
rect 8353 3782 8399 3834
rect 8399 3782 8409 3834
rect 8433 3782 8463 3834
rect 8463 3782 8489 3834
rect 8193 3780 8249 3782
rect 8273 3780 8329 3782
rect 8353 3780 8409 3782
rect 8433 3780 8489 3782
rect 6384 2202 6440 2204
rect 6464 2202 6520 2204
rect 6544 2202 6600 2204
rect 6624 2202 6680 2204
rect 6384 2150 6410 2202
rect 6410 2150 6440 2202
rect 6464 2150 6474 2202
rect 6474 2150 6520 2202
rect 6544 2150 6590 2202
rect 6590 2150 6600 2202
rect 6624 2150 6654 2202
rect 6654 2150 6680 2202
rect 6384 2148 6440 2150
rect 6464 2148 6520 2150
rect 6544 2148 6600 2150
rect 6624 2148 6680 2150
rect 8193 2746 8249 2748
rect 8273 2746 8329 2748
rect 8353 2746 8409 2748
rect 8433 2746 8489 2748
rect 8193 2694 8219 2746
rect 8219 2694 8249 2746
rect 8273 2694 8283 2746
rect 8283 2694 8329 2746
rect 8353 2694 8399 2746
rect 8399 2694 8409 2746
rect 8433 2694 8463 2746
rect 8463 2694 8489 2746
rect 8193 2692 8249 2694
rect 8273 2692 8329 2694
rect 8353 2692 8409 2694
rect 8433 2692 8489 2694
rect 10002 8730 10058 8732
rect 10082 8730 10138 8732
rect 10162 8730 10218 8732
rect 10242 8730 10298 8732
rect 10002 8678 10028 8730
rect 10028 8678 10058 8730
rect 10082 8678 10092 8730
rect 10092 8678 10138 8730
rect 10162 8678 10208 8730
rect 10208 8678 10218 8730
rect 10242 8678 10272 8730
rect 10272 8678 10298 8730
rect 10002 8676 10058 8678
rect 10082 8676 10138 8678
rect 10162 8676 10218 8678
rect 10242 8676 10298 8678
rect 10002 7642 10058 7644
rect 10082 7642 10138 7644
rect 10162 7642 10218 7644
rect 10242 7642 10298 7644
rect 10002 7590 10028 7642
rect 10028 7590 10058 7642
rect 10082 7590 10092 7642
rect 10092 7590 10138 7642
rect 10162 7590 10208 7642
rect 10208 7590 10218 7642
rect 10242 7590 10272 7642
rect 10272 7590 10298 7642
rect 10002 7588 10058 7590
rect 10082 7588 10138 7590
rect 10162 7588 10218 7590
rect 10242 7588 10298 7590
rect 10046 6840 10102 6896
rect 10002 6554 10058 6556
rect 10082 6554 10138 6556
rect 10162 6554 10218 6556
rect 10242 6554 10298 6556
rect 10002 6502 10028 6554
rect 10028 6502 10058 6554
rect 10082 6502 10092 6554
rect 10092 6502 10138 6554
rect 10162 6502 10208 6554
rect 10208 6502 10218 6554
rect 10242 6502 10272 6554
rect 10272 6502 10298 6554
rect 10002 6500 10058 6502
rect 10082 6500 10138 6502
rect 10162 6500 10218 6502
rect 10242 6500 10298 6502
rect 10690 8880 10746 8936
rect 9034 1264 9090 1320
rect 9862 6160 9918 6216
rect 10002 5466 10058 5468
rect 10082 5466 10138 5468
rect 10162 5466 10218 5468
rect 10242 5466 10298 5468
rect 10002 5414 10028 5466
rect 10028 5414 10058 5466
rect 10082 5414 10092 5466
rect 10092 5414 10138 5466
rect 10162 5414 10208 5466
rect 10208 5414 10218 5466
rect 10242 5414 10272 5466
rect 10272 5414 10298 5466
rect 10002 5412 10058 5414
rect 10082 5412 10138 5414
rect 10162 5412 10218 5414
rect 10242 5412 10298 5414
rect 10782 7284 10784 7304
rect 10784 7284 10836 7304
rect 10836 7284 10838 7304
rect 10782 7248 10838 7284
rect 10874 6296 10930 6352
rect 10002 4378 10058 4380
rect 10082 4378 10138 4380
rect 10162 4378 10218 4380
rect 10242 4378 10298 4380
rect 10002 4326 10028 4378
rect 10028 4326 10058 4378
rect 10082 4326 10092 4378
rect 10092 4326 10138 4378
rect 10162 4326 10208 4378
rect 10208 4326 10218 4378
rect 10242 4326 10272 4378
rect 10272 4326 10298 4378
rect 10002 4324 10058 4326
rect 10082 4324 10138 4326
rect 10162 4324 10218 4326
rect 10242 4324 10298 4326
rect 9586 3712 9642 3768
rect 10002 3290 10058 3292
rect 10082 3290 10138 3292
rect 10162 3290 10218 3292
rect 10242 3290 10298 3292
rect 10002 3238 10028 3290
rect 10028 3238 10058 3290
rect 10082 3238 10092 3290
rect 10092 3238 10138 3290
rect 10162 3238 10208 3290
rect 10208 3238 10218 3290
rect 10242 3238 10272 3290
rect 10272 3238 10298 3290
rect 10002 3236 10058 3238
rect 10082 3236 10138 3238
rect 10162 3236 10218 3238
rect 10242 3236 10298 3238
rect 10002 2202 10058 2204
rect 10082 2202 10138 2204
rect 10162 2202 10218 2204
rect 10242 2202 10298 2204
rect 10002 2150 10028 2202
rect 10028 2150 10058 2202
rect 10082 2150 10092 2202
rect 10092 2150 10138 2202
rect 10162 2150 10208 2202
rect 10208 2150 10218 2202
rect 10242 2150 10272 2202
rect 10272 2150 10298 2202
rect 10002 2148 10058 2150
rect 10082 2148 10138 2150
rect 10162 2148 10218 2150
rect 10242 2148 10298 2150
<< metal3 >>
rect 0 13970 800 14000
rect 3417 13970 3483 13973
rect 0 13968 3483 13970
rect 0 13912 3422 13968
rect 3478 13912 3483 13968
rect 0 13910 3483 13912
rect 0 13880 800 13910
rect 3417 13907 3483 13910
rect 9581 13970 9647 13973
rect 12296 13970 13096 14000
rect 9581 13968 13096 13970
rect 9581 13912 9586 13968
rect 9642 13912 13096 13968
rect 9581 13910 13096 13912
rect 9581 13907 9647 13910
rect 12296 13880 13096 13910
rect 2753 13088 3073 13089
rect 2753 13024 2761 13088
rect 2825 13024 2841 13088
rect 2905 13024 2921 13088
rect 2985 13024 3001 13088
rect 3065 13024 3073 13088
rect 2753 13023 3073 13024
rect 6372 13088 6692 13089
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 13023 6692 13024
rect 9990 13088 10310 13089
rect 9990 13024 9998 13088
rect 10062 13024 10078 13088
rect 10142 13024 10158 13088
rect 10222 13024 10238 13088
rect 10302 13024 10310 13088
rect 9990 13023 10310 13024
rect 4562 12544 4882 12545
rect 4562 12480 4570 12544
rect 4634 12480 4650 12544
rect 4714 12480 4730 12544
rect 4794 12480 4810 12544
rect 4874 12480 4882 12544
rect 4562 12479 4882 12480
rect 8181 12544 8501 12545
rect 8181 12480 8189 12544
rect 8253 12480 8269 12544
rect 8333 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8501 12544
rect 8181 12479 8501 12480
rect 2753 12000 3073 12001
rect 2753 11936 2761 12000
rect 2825 11936 2841 12000
rect 2905 11936 2921 12000
rect 2985 11936 3001 12000
rect 3065 11936 3073 12000
rect 2753 11935 3073 11936
rect 6372 12000 6692 12001
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 11935 6692 11936
rect 9990 12000 10310 12001
rect 9990 11936 9998 12000
rect 10062 11936 10078 12000
rect 10142 11936 10158 12000
rect 10222 11936 10238 12000
rect 10302 11936 10310 12000
rect 9990 11935 10310 11936
rect 4562 11456 4882 11457
rect 0 11386 800 11416
rect 4562 11392 4570 11456
rect 4634 11392 4650 11456
rect 4714 11392 4730 11456
rect 4794 11392 4810 11456
rect 4874 11392 4882 11456
rect 4562 11391 4882 11392
rect 8181 11456 8501 11457
rect 8181 11392 8189 11456
rect 8253 11392 8269 11456
rect 8333 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8501 11456
rect 8181 11391 8501 11392
rect 1945 11386 2011 11389
rect 0 11384 2011 11386
rect 0 11328 1950 11384
rect 2006 11328 2011 11384
rect 0 11326 2011 11328
rect 0 11296 800 11326
rect 1945 11323 2011 11326
rect 8569 11386 8635 11389
rect 12296 11386 13096 11416
rect 8569 11384 13096 11386
rect 8569 11328 8574 11384
rect 8630 11328 13096 11384
rect 8569 11326 13096 11328
rect 8569 11323 8635 11326
rect 12296 11296 13096 11326
rect 2753 10912 3073 10913
rect 2753 10848 2761 10912
rect 2825 10848 2841 10912
rect 2905 10848 2921 10912
rect 2985 10848 3001 10912
rect 3065 10848 3073 10912
rect 2753 10847 3073 10848
rect 6372 10912 6692 10913
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 10847 6692 10848
rect 9990 10912 10310 10913
rect 9990 10848 9998 10912
rect 10062 10848 10078 10912
rect 10142 10848 10158 10912
rect 10222 10848 10238 10912
rect 10302 10848 10310 10912
rect 9990 10847 10310 10848
rect 4562 10368 4882 10369
rect 4562 10304 4570 10368
rect 4634 10304 4650 10368
rect 4714 10304 4730 10368
rect 4794 10304 4810 10368
rect 4874 10304 4882 10368
rect 4562 10303 4882 10304
rect 8181 10368 8501 10369
rect 8181 10304 8189 10368
rect 8253 10304 8269 10368
rect 8333 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8501 10368
rect 8181 10303 8501 10304
rect 2753 9824 3073 9825
rect 2753 9760 2761 9824
rect 2825 9760 2841 9824
rect 2905 9760 2921 9824
rect 2985 9760 3001 9824
rect 3065 9760 3073 9824
rect 2753 9759 3073 9760
rect 6372 9824 6692 9825
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6372 9759 6692 9760
rect 9990 9824 10310 9825
rect 9990 9760 9998 9824
rect 10062 9760 10078 9824
rect 10142 9760 10158 9824
rect 10222 9760 10238 9824
rect 10302 9760 10310 9824
rect 9990 9759 10310 9760
rect 7465 9618 7531 9621
rect 7649 9618 7715 9621
rect 7465 9616 7715 9618
rect 7465 9560 7470 9616
rect 7526 9560 7654 9616
rect 7710 9560 7715 9616
rect 7465 9558 7715 9560
rect 7465 9555 7531 9558
rect 7649 9555 7715 9558
rect 6453 9482 6519 9485
rect 8201 9482 8267 9485
rect 6453 9480 8267 9482
rect 6453 9424 6458 9480
rect 6514 9424 8206 9480
rect 8262 9424 8267 9480
rect 6453 9422 8267 9424
rect 6453 9419 6519 9422
rect 8201 9419 8267 9422
rect 4562 9280 4882 9281
rect 4562 9216 4570 9280
rect 4634 9216 4650 9280
rect 4714 9216 4730 9280
rect 4794 9216 4810 9280
rect 4874 9216 4882 9280
rect 4562 9215 4882 9216
rect 8181 9280 8501 9281
rect 8181 9216 8189 9280
rect 8253 9216 8269 9280
rect 8333 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8501 9280
rect 8181 9215 8501 9216
rect 5717 9074 5783 9077
rect 7833 9074 7899 9077
rect 5717 9072 7899 9074
rect 5717 9016 5722 9072
rect 5778 9016 7838 9072
rect 7894 9016 7899 9072
rect 5717 9014 7899 9016
rect 5717 9011 5783 9014
rect 0 8938 800 8968
rect 7560 8941 7620 9014
rect 7833 9011 7899 9014
rect 3509 8938 3575 8941
rect 0 8936 3575 8938
rect 0 8880 3514 8936
rect 3570 8880 3575 8936
rect 0 8878 3575 8880
rect 0 8848 800 8878
rect 3509 8875 3575 8878
rect 3785 8938 3851 8941
rect 6126 8938 6132 8940
rect 3785 8936 6132 8938
rect 3785 8880 3790 8936
rect 3846 8880 6132 8936
rect 3785 8878 6132 8880
rect 3785 8875 3851 8878
rect 6126 8876 6132 8878
rect 6196 8938 6202 8940
rect 6453 8938 6519 8941
rect 6196 8936 6519 8938
rect 6196 8880 6458 8936
rect 6514 8880 6519 8936
rect 6196 8878 6519 8880
rect 6196 8876 6202 8878
rect 6453 8875 6519 8878
rect 7557 8936 7623 8941
rect 7557 8880 7562 8936
rect 7618 8880 7623 8936
rect 7557 8875 7623 8880
rect 10685 8938 10751 8941
rect 12296 8938 13096 8968
rect 10685 8936 13096 8938
rect 10685 8880 10690 8936
rect 10746 8880 13096 8936
rect 10685 8878 13096 8880
rect 10685 8875 10751 8878
rect 12296 8848 13096 8878
rect 7925 8802 7991 8805
rect 7606 8800 7991 8802
rect 7606 8744 7930 8800
rect 7986 8744 7991 8800
rect 7606 8742 7991 8744
rect 2753 8736 3073 8737
rect 2753 8672 2761 8736
rect 2825 8672 2841 8736
rect 2905 8672 2921 8736
rect 2985 8672 3001 8736
rect 3065 8672 3073 8736
rect 2753 8671 3073 8672
rect 6372 8736 6692 8737
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 8671 6692 8672
rect 7465 8258 7531 8261
rect 7606 8258 7666 8742
rect 7925 8739 7991 8742
rect 9990 8736 10310 8737
rect 9990 8672 9998 8736
rect 10062 8672 10078 8736
rect 10142 8672 10158 8736
rect 10222 8672 10238 8736
rect 10302 8672 10310 8736
rect 9990 8671 10310 8672
rect 7925 8394 7991 8397
rect 8477 8394 8543 8397
rect 7925 8392 8543 8394
rect 7925 8336 7930 8392
rect 7986 8336 8482 8392
rect 8538 8336 8543 8392
rect 7925 8334 8543 8336
rect 7925 8331 7991 8334
rect 8477 8331 8543 8334
rect 7465 8256 7666 8258
rect 7465 8200 7470 8256
rect 7526 8200 7666 8256
rect 7465 8198 7666 8200
rect 7465 8195 7531 8198
rect 4562 8192 4882 8193
rect 4562 8128 4570 8192
rect 4634 8128 4650 8192
rect 4714 8128 4730 8192
rect 4794 8128 4810 8192
rect 4874 8128 4882 8192
rect 4562 8127 4882 8128
rect 8181 8192 8501 8193
rect 8181 8128 8189 8192
rect 8253 8128 8269 8192
rect 8333 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8501 8192
rect 8181 8127 8501 8128
rect 2405 7986 2471 7989
rect 8385 7986 8451 7989
rect 2405 7984 8451 7986
rect 2405 7928 2410 7984
rect 2466 7928 8390 7984
rect 8446 7928 8451 7984
rect 2405 7926 8451 7928
rect 2405 7923 2471 7926
rect 8385 7923 8451 7926
rect 7925 7850 7991 7853
rect 9397 7850 9463 7853
rect 7925 7848 9463 7850
rect 7925 7792 7930 7848
rect 7986 7792 9402 7848
rect 9458 7792 9463 7848
rect 7925 7790 9463 7792
rect 7925 7787 7991 7790
rect 9397 7787 9463 7790
rect 7649 7714 7715 7717
rect 9213 7714 9279 7717
rect 7649 7712 9279 7714
rect 7649 7656 7654 7712
rect 7710 7656 9218 7712
rect 9274 7656 9279 7712
rect 7649 7654 9279 7656
rect 7649 7651 7715 7654
rect 9213 7651 9279 7654
rect 2753 7648 3073 7649
rect 2753 7584 2761 7648
rect 2825 7584 2841 7648
rect 2905 7584 2921 7648
rect 2985 7584 3001 7648
rect 3065 7584 3073 7648
rect 2753 7583 3073 7584
rect 6372 7648 6692 7649
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 7583 6692 7584
rect 9990 7648 10310 7649
rect 9990 7584 9998 7648
rect 10062 7584 10078 7648
rect 10142 7584 10158 7648
rect 10222 7584 10238 7648
rect 10302 7584 10310 7648
rect 9990 7583 10310 7584
rect 6085 7578 6151 7581
rect 5030 7576 6151 7578
rect 5030 7520 6090 7576
rect 6146 7520 6151 7576
rect 5030 7518 6151 7520
rect 2313 7442 2379 7445
rect 5030 7442 5090 7518
rect 6085 7515 6151 7518
rect 7189 7578 7255 7581
rect 8569 7578 8635 7581
rect 7189 7576 8635 7578
rect 7189 7520 7194 7576
rect 7250 7520 8574 7576
rect 8630 7520 8635 7576
rect 7189 7518 8635 7520
rect 7189 7515 7255 7518
rect 8569 7515 8635 7518
rect 2313 7440 5090 7442
rect 2313 7384 2318 7440
rect 2374 7384 5090 7440
rect 2313 7382 5090 7384
rect 5165 7442 5231 7445
rect 7833 7442 7899 7445
rect 5165 7440 7899 7442
rect 5165 7384 5170 7440
rect 5226 7384 7838 7440
rect 7894 7384 7899 7440
rect 5165 7382 7899 7384
rect 2313 7379 2379 7382
rect 5165 7379 5231 7382
rect 7833 7379 7899 7382
rect 3141 7306 3207 7309
rect 5625 7306 5691 7309
rect 5901 7306 5967 7309
rect 3141 7304 5967 7306
rect 3141 7248 3146 7304
rect 3202 7248 5630 7304
rect 5686 7248 5906 7304
rect 5962 7248 5967 7304
rect 3141 7246 5967 7248
rect 3141 7243 3207 7246
rect 5625 7243 5691 7246
rect 5901 7243 5967 7246
rect 7833 7306 7899 7309
rect 10777 7306 10843 7309
rect 7833 7304 10843 7306
rect 7833 7248 7838 7304
rect 7894 7248 10782 7304
rect 10838 7248 10843 7304
rect 7833 7246 10843 7248
rect 7833 7243 7899 7246
rect 10777 7243 10843 7246
rect 5257 7170 5323 7173
rect 6177 7170 6243 7173
rect 5257 7168 6243 7170
rect 5257 7112 5262 7168
rect 5318 7112 6182 7168
rect 6238 7112 6243 7168
rect 5257 7110 6243 7112
rect 5257 7107 5323 7110
rect 6177 7107 6243 7110
rect 4562 7104 4882 7105
rect 4562 7040 4570 7104
rect 4634 7040 4650 7104
rect 4714 7040 4730 7104
rect 4794 7040 4810 7104
rect 4874 7040 4882 7104
rect 4562 7039 4882 7040
rect 8181 7104 8501 7105
rect 8181 7040 8189 7104
rect 8253 7040 8269 7104
rect 8333 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8501 7104
rect 8181 7039 8501 7040
rect 6821 7036 6887 7037
rect 6821 7032 6868 7036
rect 6932 7034 6938 7036
rect 6821 6976 6826 7032
rect 6821 6972 6868 6976
rect 6932 6974 6978 7034
rect 6932 6972 6938 6974
rect 6821 6971 6887 6972
rect 7557 6898 7623 6901
rect 10041 6898 10107 6901
rect 5214 6896 10107 6898
rect 5214 6840 7562 6896
rect 7618 6840 10046 6896
rect 10102 6840 10107 6896
rect 5214 6838 10107 6840
rect 3141 6762 3207 6765
rect 5214 6762 5274 6838
rect 7557 6835 7623 6838
rect 10041 6835 10107 6838
rect 3141 6760 5274 6762
rect 3141 6704 3146 6760
rect 3202 6704 5274 6760
rect 3141 6702 5274 6704
rect 6453 6762 6519 6765
rect 6453 6760 6930 6762
rect 6453 6704 6458 6760
rect 6514 6704 6930 6760
rect 6453 6702 6930 6704
rect 3141 6699 3207 6702
rect 6453 6699 6519 6702
rect 6870 6626 6930 6702
rect 7649 6626 7715 6629
rect 6870 6624 7715 6626
rect 6870 6568 7654 6624
rect 7710 6568 7715 6624
rect 6870 6566 7715 6568
rect 7649 6563 7715 6566
rect 2753 6560 3073 6561
rect 2753 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2921 6560
rect 2985 6496 3001 6560
rect 3065 6496 3073 6560
rect 2753 6495 3073 6496
rect 6372 6560 6692 6561
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6372 6495 6692 6496
rect 9990 6560 10310 6561
rect 9990 6496 9998 6560
rect 10062 6496 10078 6560
rect 10142 6496 10158 6560
rect 10222 6496 10238 6560
rect 10302 6496 10310 6560
rect 9990 6495 10310 6496
rect 0 6354 800 6384
rect 3969 6354 4035 6357
rect 0 6352 4035 6354
rect 0 6296 3974 6352
rect 4030 6296 4035 6352
rect 0 6294 4035 6296
rect 0 6264 800 6294
rect 3969 6291 4035 6294
rect 6177 6354 6243 6357
rect 6545 6354 6611 6357
rect 9029 6354 9095 6357
rect 6177 6352 9095 6354
rect 6177 6296 6182 6352
rect 6238 6296 6550 6352
rect 6606 6296 9034 6352
rect 9090 6296 9095 6352
rect 6177 6294 9095 6296
rect 6177 6291 6243 6294
rect 6545 6291 6611 6294
rect 9029 6291 9095 6294
rect 10869 6354 10935 6357
rect 12296 6354 13096 6384
rect 10869 6352 13096 6354
rect 10869 6296 10874 6352
rect 10930 6296 13096 6352
rect 10869 6294 13096 6296
rect 10869 6291 10935 6294
rect 12296 6264 13096 6294
rect 5073 6218 5139 6221
rect 5625 6218 5691 6221
rect 9857 6218 9923 6221
rect 5073 6216 9923 6218
rect 5073 6160 5078 6216
rect 5134 6160 5630 6216
rect 5686 6160 9862 6216
rect 9918 6160 9923 6216
rect 5073 6158 9923 6160
rect 5073 6155 5139 6158
rect 5625 6155 5691 6158
rect 9857 6155 9923 6158
rect 6177 6084 6243 6085
rect 6126 6020 6132 6084
rect 6196 6082 6243 6084
rect 6637 6082 6703 6085
rect 6862 6082 6868 6084
rect 6196 6080 6288 6082
rect 6238 6024 6288 6080
rect 6196 6022 6288 6024
rect 6637 6080 6868 6082
rect 6637 6024 6642 6080
rect 6698 6024 6868 6080
rect 6637 6022 6868 6024
rect 6196 6020 6243 6022
rect 6177 6019 6243 6020
rect 6637 6019 6703 6022
rect 6862 6020 6868 6022
rect 6932 6020 6938 6084
rect 4562 6016 4882 6017
rect 4562 5952 4570 6016
rect 4634 5952 4650 6016
rect 4714 5952 4730 6016
rect 4794 5952 4810 6016
rect 4874 5952 4882 6016
rect 4562 5951 4882 5952
rect 8181 6016 8501 6017
rect 8181 5952 8189 6016
rect 8253 5952 8269 6016
rect 8333 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8501 6016
rect 8181 5951 8501 5952
rect 6361 5810 6427 5813
rect 7465 5810 7531 5813
rect 6361 5808 7531 5810
rect 6361 5752 6366 5808
rect 6422 5752 7470 5808
rect 7526 5752 7531 5808
rect 6361 5750 7531 5752
rect 6361 5747 6427 5750
rect 7465 5747 7531 5750
rect 6729 5674 6795 5677
rect 8109 5674 8175 5677
rect 6729 5672 8175 5674
rect 6729 5616 6734 5672
rect 6790 5616 8114 5672
rect 8170 5616 8175 5672
rect 6729 5614 8175 5616
rect 6729 5611 6795 5614
rect 8109 5611 8175 5614
rect 2753 5472 3073 5473
rect 2753 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2921 5472
rect 2985 5408 3001 5472
rect 3065 5408 3073 5472
rect 2753 5407 3073 5408
rect 6372 5472 6692 5473
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 5407 6692 5408
rect 9990 5472 10310 5473
rect 9990 5408 9998 5472
rect 10062 5408 10078 5472
rect 10142 5408 10158 5472
rect 10222 5408 10238 5472
rect 10302 5408 10310 5472
rect 9990 5407 10310 5408
rect 6269 5266 6335 5269
rect 6913 5266 6979 5269
rect 6269 5264 6979 5266
rect 6269 5208 6274 5264
rect 6330 5208 6918 5264
rect 6974 5208 6979 5264
rect 6269 5206 6979 5208
rect 6269 5203 6335 5206
rect 6913 5203 6979 5206
rect 4981 4994 5047 4997
rect 7097 4994 7163 4997
rect 7741 4994 7807 4997
rect 4981 4992 7807 4994
rect 4981 4936 4986 4992
rect 5042 4936 7102 4992
rect 7158 4936 7746 4992
rect 7802 4936 7807 4992
rect 4981 4934 7807 4936
rect 4981 4931 5047 4934
rect 7097 4931 7163 4934
rect 7741 4931 7807 4934
rect 4562 4928 4882 4929
rect 4562 4864 4570 4928
rect 4634 4864 4650 4928
rect 4714 4864 4730 4928
rect 4794 4864 4810 4928
rect 4874 4864 4882 4928
rect 4562 4863 4882 4864
rect 8181 4928 8501 4929
rect 8181 4864 8189 4928
rect 8253 4864 8269 4928
rect 8333 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8501 4928
rect 8181 4863 8501 4864
rect 6637 4722 6703 4725
rect 8017 4722 8083 4725
rect 6637 4720 8083 4722
rect 6637 4664 6642 4720
rect 6698 4664 8022 4720
rect 8078 4664 8083 4720
rect 6637 4662 8083 4664
rect 6637 4659 6703 4662
rect 8017 4659 8083 4662
rect 2753 4384 3073 4385
rect 2753 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2921 4384
rect 2985 4320 3001 4384
rect 3065 4320 3073 4384
rect 2753 4319 3073 4320
rect 6372 4384 6692 4385
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 4319 6692 4320
rect 9990 4384 10310 4385
rect 9990 4320 9998 4384
rect 10062 4320 10078 4384
rect 10142 4320 10158 4384
rect 10222 4320 10238 4384
rect 10302 4320 10310 4384
rect 9990 4319 10310 4320
rect 4562 3840 4882 3841
rect 0 3770 800 3800
rect 4562 3776 4570 3840
rect 4634 3776 4650 3840
rect 4714 3776 4730 3840
rect 4794 3776 4810 3840
rect 4874 3776 4882 3840
rect 4562 3775 4882 3776
rect 8181 3840 8501 3841
rect 8181 3776 8189 3840
rect 8253 3776 8269 3840
rect 8333 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8501 3840
rect 8181 3775 8501 3776
rect 3877 3770 3943 3773
rect 0 3768 3943 3770
rect 0 3712 3882 3768
rect 3938 3712 3943 3768
rect 0 3710 3943 3712
rect 0 3680 800 3710
rect 3877 3707 3943 3710
rect 9581 3770 9647 3773
rect 12296 3770 13096 3800
rect 9581 3768 13096 3770
rect 9581 3712 9586 3768
rect 9642 3712 13096 3768
rect 9581 3710 13096 3712
rect 9581 3707 9647 3710
rect 12296 3680 13096 3710
rect 2753 3296 3073 3297
rect 2753 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2921 3296
rect 2985 3232 3001 3296
rect 3065 3232 3073 3296
rect 2753 3231 3073 3232
rect 6372 3296 6692 3297
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 3231 6692 3232
rect 9990 3296 10310 3297
rect 9990 3232 9998 3296
rect 10062 3232 10078 3296
rect 10142 3232 10158 3296
rect 10222 3232 10238 3296
rect 10302 3232 10310 3296
rect 9990 3231 10310 3232
rect 4562 2752 4882 2753
rect 4562 2688 4570 2752
rect 4634 2688 4650 2752
rect 4714 2688 4730 2752
rect 4794 2688 4810 2752
rect 4874 2688 4882 2752
rect 4562 2687 4882 2688
rect 8181 2752 8501 2753
rect 8181 2688 8189 2752
rect 8253 2688 8269 2752
rect 8333 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8501 2752
rect 8181 2687 8501 2688
rect 2753 2208 3073 2209
rect 2753 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2921 2208
rect 2985 2144 3001 2208
rect 3065 2144 3073 2208
rect 2753 2143 3073 2144
rect 6372 2208 6692 2209
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2143 6692 2144
rect 9990 2208 10310 2209
rect 9990 2144 9998 2208
rect 10062 2144 10078 2208
rect 10142 2144 10158 2208
rect 10222 2144 10238 2208
rect 10302 2144 10310 2208
rect 9990 2143 10310 2144
rect 0 1322 800 1352
rect 3601 1322 3667 1325
rect 0 1320 3667 1322
rect 0 1264 3606 1320
rect 3662 1264 3667 1320
rect 0 1262 3667 1264
rect 0 1232 800 1262
rect 3601 1259 3667 1262
rect 9029 1322 9095 1325
rect 12296 1322 13096 1352
rect 9029 1320 13096 1322
rect 9029 1264 9034 1320
rect 9090 1264 13096 1320
rect 9029 1262 13096 1264
rect 9029 1259 9095 1262
rect 12296 1232 13096 1262
<< via3 >>
rect 2761 13084 2825 13088
rect 2761 13028 2765 13084
rect 2765 13028 2821 13084
rect 2821 13028 2825 13084
rect 2761 13024 2825 13028
rect 2841 13084 2905 13088
rect 2841 13028 2845 13084
rect 2845 13028 2901 13084
rect 2901 13028 2905 13084
rect 2841 13024 2905 13028
rect 2921 13084 2985 13088
rect 2921 13028 2925 13084
rect 2925 13028 2981 13084
rect 2981 13028 2985 13084
rect 2921 13024 2985 13028
rect 3001 13084 3065 13088
rect 3001 13028 3005 13084
rect 3005 13028 3061 13084
rect 3061 13028 3065 13084
rect 3001 13024 3065 13028
rect 6380 13084 6444 13088
rect 6380 13028 6384 13084
rect 6384 13028 6440 13084
rect 6440 13028 6444 13084
rect 6380 13024 6444 13028
rect 6460 13084 6524 13088
rect 6460 13028 6464 13084
rect 6464 13028 6520 13084
rect 6520 13028 6524 13084
rect 6460 13024 6524 13028
rect 6540 13084 6604 13088
rect 6540 13028 6544 13084
rect 6544 13028 6600 13084
rect 6600 13028 6604 13084
rect 6540 13024 6604 13028
rect 6620 13084 6684 13088
rect 6620 13028 6624 13084
rect 6624 13028 6680 13084
rect 6680 13028 6684 13084
rect 6620 13024 6684 13028
rect 9998 13084 10062 13088
rect 9998 13028 10002 13084
rect 10002 13028 10058 13084
rect 10058 13028 10062 13084
rect 9998 13024 10062 13028
rect 10078 13084 10142 13088
rect 10078 13028 10082 13084
rect 10082 13028 10138 13084
rect 10138 13028 10142 13084
rect 10078 13024 10142 13028
rect 10158 13084 10222 13088
rect 10158 13028 10162 13084
rect 10162 13028 10218 13084
rect 10218 13028 10222 13084
rect 10158 13024 10222 13028
rect 10238 13084 10302 13088
rect 10238 13028 10242 13084
rect 10242 13028 10298 13084
rect 10298 13028 10302 13084
rect 10238 13024 10302 13028
rect 4570 12540 4634 12544
rect 4570 12484 4574 12540
rect 4574 12484 4630 12540
rect 4630 12484 4634 12540
rect 4570 12480 4634 12484
rect 4650 12540 4714 12544
rect 4650 12484 4654 12540
rect 4654 12484 4710 12540
rect 4710 12484 4714 12540
rect 4650 12480 4714 12484
rect 4730 12540 4794 12544
rect 4730 12484 4734 12540
rect 4734 12484 4790 12540
rect 4790 12484 4794 12540
rect 4730 12480 4794 12484
rect 4810 12540 4874 12544
rect 4810 12484 4814 12540
rect 4814 12484 4870 12540
rect 4870 12484 4874 12540
rect 4810 12480 4874 12484
rect 8189 12540 8253 12544
rect 8189 12484 8193 12540
rect 8193 12484 8249 12540
rect 8249 12484 8253 12540
rect 8189 12480 8253 12484
rect 8269 12540 8333 12544
rect 8269 12484 8273 12540
rect 8273 12484 8329 12540
rect 8329 12484 8333 12540
rect 8269 12480 8333 12484
rect 8349 12540 8413 12544
rect 8349 12484 8353 12540
rect 8353 12484 8409 12540
rect 8409 12484 8413 12540
rect 8349 12480 8413 12484
rect 8429 12540 8493 12544
rect 8429 12484 8433 12540
rect 8433 12484 8489 12540
rect 8489 12484 8493 12540
rect 8429 12480 8493 12484
rect 2761 11996 2825 12000
rect 2761 11940 2765 11996
rect 2765 11940 2821 11996
rect 2821 11940 2825 11996
rect 2761 11936 2825 11940
rect 2841 11996 2905 12000
rect 2841 11940 2845 11996
rect 2845 11940 2901 11996
rect 2901 11940 2905 11996
rect 2841 11936 2905 11940
rect 2921 11996 2985 12000
rect 2921 11940 2925 11996
rect 2925 11940 2981 11996
rect 2981 11940 2985 11996
rect 2921 11936 2985 11940
rect 3001 11996 3065 12000
rect 3001 11940 3005 11996
rect 3005 11940 3061 11996
rect 3061 11940 3065 11996
rect 3001 11936 3065 11940
rect 6380 11996 6444 12000
rect 6380 11940 6384 11996
rect 6384 11940 6440 11996
rect 6440 11940 6444 11996
rect 6380 11936 6444 11940
rect 6460 11996 6524 12000
rect 6460 11940 6464 11996
rect 6464 11940 6520 11996
rect 6520 11940 6524 11996
rect 6460 11936 6524 11940
rect 6540 11996 6604 12000
rect 6540 11940 6544 11996
rect 6544 11940 6600 11996
rect 6600 11940 6604 11996
rect 6540 11936 6604 11940
rect 6620 11996 6684 12000
rect 6620 11940 6624 11996
rect 6624 11940 6680 11996
rect 6680 11940 6684 11996
rect 6620 11936 6684 11940
rect 9998 11996 10062 12000
rect 9998 11940 10002 11996
rect 10002 11940 10058 11996
rect 10058 11940 10062 11996
rect 9998 11936 10062 11940
rect 10078 11996 10142 12000
rect 10078 11940 10082 11996
rect 10082 11940 10138 11996
rect 10138 11940 10142 11996
rect 10078 11936 10142 11940
rect 10158 11996 10222 12000
rect 10158 11940 10162 11996
rect 10162 11940 10218 11996
rect 10218 11940 10222 11996
rect 10158 11936 10222 11940
rect 10238 11996 10302 12000
rect 10238 11940 10242 11996
rect 10242 11940 10298 11996
rect 10298 11940 10302 11996
rect 10238 11936 10302 11940
rect 4570 11452 4634 11456
rect 4570 11396 4574 11452
rect 4574 11396 4630 11452
rect 4630 11396 4634 11452
rect 4570 11392 4634 11396
rect 4650 11452 4714 11456
rect 4650 11396 4654 11452
rect 4654 11396 4710 11452
rect 4710 11396 4714 11452
rect 4650 11392 4714 11396
rect 4730 11452 4794 11456
rect 4730 11396 4734 11452
rect 4734 11396 4790 11452
rect 4790 11396 4794 11452
rect 4730 11392 4794 11396
rect 4810 11452 4874 11456
rect 4810 11396 4814 11452
rect 4814 11396 4870 11452
rect 4870 11396 4874 11452
rect 4810 11392 4874 11396
rect 8189 11452 8253 11456
rect 8189 11396 8193 11452
rect 8193 11396 8249 11452
rect 8249 11396 8253 11452
rect 8189 11392 8253 11396
rect 8269 11452 8333 11456
rect 8269 11396 8273 11452
rect 8273 11396 8329 11452
rect 8329 11396 8333 11452
rect 8269 11392 8333 11396
rect 8349 11452 8413 11456
rect 8349 11396 8353 11452
rect 8353 11396 8409 11452
rect 8409 11396 8413 11452
rect 8349 11392 8413 11396
rect 8429 11452 8493 11456
rect 8429 11396 8433 11452
rect 8433 11396 8489 11452
rect 8489 11396 8493 11452
rect 8429 11392 8493 11396
rect 2761 10908 2825 10912
rect 2761 10852 2765 10908
rect 2765 10852 2821 10908
rect 2821 10852 2825 10908
rect 2761 10848 2825 10852
rect 2841 10908 2905 10912
rect 2841 10852 2845 10908
rect 2845 10852 2901 10908
rect 2901 10852 2905 10908
rect 2841 10848 2905 10852
rect 2921 10908 2985 10912
rect 2921 10852 2925 10908
rect 2925 10852 2981 10908
rect 2981 10852 2985 10908
rect 2921 10848 2985 10852
rect 3001 10908 3065 10912
rect 3001 10852 3005 10908
rect 3005 10852 3061 10908
rect 3061 10852 3065 10908
rect 3001 10848 3065 10852
rect 6380 10908 6444 10912
rect 6380 10852 6384 10908
rect 6384 10852 6440 10908
rect 6440 10852 6444 10908
rect 6380 10848 6444 10852
rect 6460 10908 6524 10912
rect 6460 10852 6464 10908
rect 6464 10852 6520 10908
rect 6520 10852 6524 10908
rect 6460 10848 6524 10852
rect 6540 10908 6604 10912
rect 6540 10852 6544 10908
rect 6544 10852 6600 10908
rect 6600 10852 6604 10908
rect 6540 10848 6604 10852
rect 6620 10908 6684 10912
rect 6620 10852 6624 10908
rect 6624 10852 6680 10908
rect 6680 10852 6684 10908
rect 6620 10848 6684 10852
rect 9998 10908 10062 10912
rect 9998 10852 10002 10908
rect 10002 10852 10058 10908
rect 10058 10852 10062 10908
rect 9998 10848 10062 10852
rect 10078 10908 10142 10912
rect 10078 10852 10082 10908
rect 10082 10852 10138 10908
rect 10138 10852 10142 10908
rect 10078 10848 10142 10852
rect 10158 10908 10222 10912
rect 10158 10852 10162 10908
rect 10162 10852 10218 10908
rect 10218 10852 10222 10908
rect 10158 10848 10222 10852
rect 10238 10908 10302 10912
rect 10238 10852 10242 10908
rect 10242 10852 10298 10908
rect 10298 10852 10302 10908
rect 10238 10848 10302 10852
rect 4570 10364 4634 10368
rect 4570 10308 4574 10364
rect 4574 10308 4630 10364
rect 4630 10308 4634 10364
rect 4570 10304 4634 10308
rect 4650 10364 4714 10368
rect 4650 10308 4654 10364
rect 4654 10308 4710 10364
rect 4710 10308 4714 10364
rect 4650 10304 4714 10308
rect 4730 10364 4794 10368
rect 4730 10308 4734 10364
rect 4734 10308 4790 10364
rect 4790 10308 4794 10364
rect 4730 10304 4794 10308
rect 4810 10364 4874 10368
rect 4810 10308 4814 10364
rect 4814 10308 4870 10364
rect 4870 10308 4874 10364
rect 4810 10304 4874 10308
rect 8189 10364 8253 10368
rect 8189 10308 8193 10364
rect 8193 10308 8249 10364
rect 8249 10308 8253 10364
rect 8189 10304 8253 10308
rect 8269 10364 8333 10368
rect 8269 10308 8273 10364
rect 8273 10308 8329 10364
rect 8329 10308 8333 10364
rect 8269 10304 8333 10308
rect 8349 10364 8413 10368
rect 8349 10308 8353 10364
rect 8353 10308 8409 10364
rect 8409 10308 8413 10364
rect 8349 10304 8413 10308
rect 8429 10364 8493 10368
rect 8429 10308 8433 10364
rect 8433 10308 8489 10364
rect 8489 10308 8493 10364
rect 8429 10304 8493 10308
rect 2761 9820 2825 9824
rect 2761 9764 2765 9820
rect 2765 9764 2821 9820
rect 2821 9764 2825 9820
rect 2761 9760 2825 9764
rect 2841 9820 2905 9824
rect 2841 9764 2845 9820
rect 2845 9764 2901 9820
rect 2901 9764 2905 9820
rect 2841 9760 2905 9764
rect 2921 9820 2985 9824
rect 2921 9764 2925 9820
rect 2925 9764 2981 9820
rect 2981 9764 2985 9820
rect 2921 9760 2985 9764
rect 3001 9820 3065 9824
rect 3001 9764 3005 9820
rect 3005 9764 3061 9820
rect 3061 9764 3065 9820
rect 3001 9760 3065 9764
rect 6380 9820 6444 9824
rect 6380 9764 6384 9820
rect 6384 9764 6440 9820
rect 6440 9764 6444 9820
rect 6380 9760 6444 9764
rect 6460 9820 6524 9824
rect 6460 9764 6464 9820
rect 6464 9764 6520 9820
rect 6520 9764 6524 9820
rect 6460 9760 6524 9764
rect 6540 9820 6604 9824
rect 6540 9764 6544 9820
rect 6544 9764 6600 9820
rect 6600 9764 6604 9820
rect 6540 9760 6604 9764
rect 6620 9820 6684 9824
rect 6620 9764 6624 9820
rect 6624 9764 6680 9820
rect 6680 9764 6684 9820
rect 6620 9760 6684 9764
rect 9998 9820 10062 9824
rect 9998 9764 10002 9820
rect 10002 9764 10058 9820
rect 10058 9764 10062 9820
rect 9998 9760 10062 9764
rect 10078 9820 10142 9824
rect 10078 9764 10082 9820
rect 10082 9764 10138 9820
rect 10138 9764 10142 9820
rect 10078 9760 10142 9764
rect 10158 9820 10222 9824
rect 10158 9764 10162 9820
rect 10162 9764 10218 9820
rect 10218 9764 10222 9820
rect 10158 9760 10222 9764
rect 10238 9820 10302 9824
rect 10238 9764 10242 9820
rect 10242 9764 10298 9820
rect 10298 9764 10302 9820
rect 10238 9760 10302 9764
rect 4570 9276 4634 9280
rect 4570 9220 4574 9276
rect 4574 9220 4630 9276
rect 4630 9220 4634 9276
rect 4570 9216 4634 9220
rect 4650 9276 4714 9280
rect 4650 9220 4654 9276
rect 4654 9220 4710 9276
rect 4710 9220 4714 9276
rect 4650 9216 4714 9220
rect 4730 9276 4794 9280
rect 4730 9220 4734 9276
rect 4734 9220 4790 9276
rect 4790 9220 4794 9276
rect 4730 9216 4794 9220
rect 4810 9276 4874 9280
rect 4810 9220 4814 9276
rect 4814 9220 4870 9276
rect 4870 9220 4874 9276
rect 4810 9216 4874 9220
rect 8189 9276 8253 9280
rect 8189 9220 8193 9276
rect 8193 9220 8249 9276
rect 8249 9220 8253 9276
rect 8189 9216 8253 9220
rect 8269 9276 8333 9280
rect 8269 9220 8273 9276
rect 8273 9220 8329 9276
rect 8329 9220 8333 9276
rect 8269 9216 8333 9220
rect 8349 9276 8413 9280
rect 8349 9220 8353 9276
rect 8353 9220 8409 9276
rect 8409 9220 8413 9276
rect 8349 9216 8413 9220
rect 8429 9276 8493 9280
rect 8429 9220 8433 9276
rect 8433 9220 8489 9276
rect 8489 9220 8493 9276
rect 8429 9216 8493 9220
rect 6132 8876 6196 8940
rect 2761 8732 2825 8736
rect 2761 8676 2765 8732
rect 2765 8676 2821 8732
rect 2821 8676 2825 8732
rect 2761 8672 2825 8676
rect 2841 8732 2905 8736
rect 2841 8676 2845 8732
rect 2845 8676 2901 8732
rect 2901 8676 2905 8732
rect 2841 8672 2905 8676
rect 2921 8732 2985 8736
rect 2921 8676 2925 8732
rect 2925 8676 2981 8732
rect 2981 8676 2985 8732
rect 2921 8672 2985 8676
rect 3001 8732 3065 8736
rect 3001 8676 3005 8732
rect 3005 8676 3061 8732
rect 3061 8676 3065 8732
rect 3001 8672 3065 8676
rect 6380 8732 6444 8736
rect 6380 8676 6384 8732
rect 6384 8676 6440 8732
rect 6440 8676 6444 8732
rect 6380 8672 6444 8676
rect 6460 8732 6524 8736
rect 6460 8676 6464 8732
rect 6464 8676 6520 8732
rect 6520 8676 6524 8732
rect 6460 8672 6524 8676
rect 6540 8732 6604 8736
rect 6540 8676 6544 8732
rect 6544 8676 6600 8732
rect 6600 8676 6604 8732
rect 6540 8672 6604 8676
rect 6620 8732 6684 8736
rect 6620 8676 6624 8732
rect 6624 8676 6680 8732
rect 6680 8676 6684 8732
rect 6620 8672 6684 8676
rect 9998 8732 10062 8736
rect 9998 8676 10002 8732
rect 10002 8676 10058 8732
rect 10058 8676 10062 8732
rect 9998 8672 10062 8676
rect 10078 8732 10142 8736
rect 10078 8676 10082 8732
rect 10082 8676 10138 8732
rect 10138 8676 10142 8732
rect 10078 8672 10142 8676
rect 10158 8732 10222 8736
rect 10158 8676 10162 8732
rect 10162 8676 10218 8732
rect 10218 8676 10222 8732
rect 10158 8672 10222 8676
rect 10238 8732 10302 8736
rect 10238 8676 10242 8732
rect 10242 8676 10298 8732
rect 10298 8676 10302 8732
rect 10238 8672 10302 8676
rect 4570 8188 4634 8192
rect 4570 8132 4574 8188
rect 4574 8132 4630 8188
rect 4630 8132 4634 8188
rect 4570 8128 4634 8132
rect 4650 8188 4714 8192
rect 4650 8132 4654 8188
rect 4654 8132 4710 8188
rect 4710 8132 4714 8188
rect 4650 8128 4714 8132
rect 4730 8188 4794 8192
rect 4730 8132 4734 8188
rect 4734 8132 4790 8188
rect 4790 8132 4794 8188
rect 4730 8128 4794 8132
rect 4810 8188 4874 8192
rect 4810 8132 4814 8188
rect 4814 8132 4870 8188
rect 4870 8132 4874 8188
rect 4810 8128 4874 8132
rect 8189 8188 8253 8192
rect 8189 8132 8193 8188
rect 8193 8132 8249 8188
rect 8249 8132 8253 8188
rect 8189 8128 8253 8132
rect 8269 8188 8333 8192
rect 8269 8132 8273 8188
rect 8273 8132 8329 8188
rect 8329 8132 8333 8188
rect 8269 8128 8333 8132
rect 8349 8188 8413 8192
rect 8349 8132 8353 8188
rect 8353 8132 8409 8188
rect 8409 8132 8413 8188
rect 8349 8128 8413 8132
rect 8429 8188 8493 8192
rect 8429 8132 8433 8188
rect 8433 8132 8489 8188
rect 8489 8132 8493 8188
rect 8429 8128 8493 8132
rect 2761 7644 2825 7648
rect 2761 7588 2765 7644
rect 2765 7588 2821 7644
rect 2821 7588 2825 7644
rect 2761 7584 2825 7588
rect 2841 7644 2905 7648
rect 2841 7588 2845 7644
rect 2845 7588 2901 7644
rect 2901 7588 2905 7644
rect 2841 7584 2905 7588
rect 2921 7644 2985 7648
rect 2921 7588 2925 7644
rect 2925 7588 2981 7644
rect 2981 7588 2985 7644
rect 2921 7584 2985 7588
rect 3001 7644 3065 7648
rect 3001 7588 3005 7644
rect 3005 7588 3061 7644
rect 3061 7588 3065 7644
rect 3001 7584 3065 7588
rect 6380 7644 6444 7648
rect 6380 7588 6384 7644
rect 6384 7588 6440 7644
rect 6440 7588 6444 7644
rect 6380 7584 6444 7588
rect 6460 7644 6524 7648
rect 6460 7588 6464 7644
rect 6464 7588 6520 7644
rect 6520 7588 6524 7644
rect 6460 7584 6524 7588
rect 6540 7644 6604 7648
rect 6540 7588 6544 7644
rect 6544 7588 6600 7644
rect 6600 7588 6604 7644
rect 6540 7584 6604 7588
rect 6620 7644 6684 7648
rect 6620 7588 6624 7644
rect 6624 7588 6680 7644
rect 6680 7588 6684 7644
rect 6620 7584 6684 7588
rect 9998 7644 10062 7648
rect 9998 7588 10002 7644
rect 10002 7588 10058 7644
rect 10058 7588 10062 7644
rect 9998 7584 10062 7588
rect 10078 7644 10142 7648
rect 10078 7588 10082 7644
rect 10082 7588 10138 7644
rect 10138 7588 10142 7644
rect 10078 7584 10142 7588
rect 10158 7644 10222 7648
rect 10158 7588 10162 7644
rect 10162 7588 10218 7644
rect 10218 7588 10222 7644
rect 10158 7584 10222 7588
rect 10238 7644 10302 7648
rect 10238 7588 10242 7644
rect 10242 7588 10298 7644
rect 10298 7588 10302 7644
rect 10238 7584 10302 7588
rect 4570 7100 4634 7104
rect 4570 7044 4574 7100
rect 4574 7044 4630 7100
rect 4630 7044 4634 7100
rect 4570 7040 4634 7044
rect 4650 7100 4714 7104
rect 4650 7044 4654 7100
rect 4654 7044 4710 7100
rect 4710 7044 4714 7100
rect 4650 7040 4714 7044
rect 4730 7100 4794 7104
rect 4730 7044 4734 7100
rect 4734 7044 4790 7100
rect 4790 7044 4794 7100
rect 4730 7040 4794 7044
rect 4810 7100 4874 7104
rect 4810 7044 4814 7100
rect 4814 7044 4870 7100
rect 4870 7044 4874 7100
rect 4810 7040 4874 7044
rect 8189 7100 8253 7104
rect 8189 7044 8193 7100
rect 8193 7044 8249 7100
rect 8249 7044 8253 7100
rect 8189 7040 8253 7044
rect 8269 7100 8333 7104
rect 8269 7044 8273 7100
rect 8273 7044 8329 7100
rect 8329 7044 8333 7100
rect 8269 7040 8333 7044
rect 8349 7100 8413 7104
rect 8349 7044 8353 7100
rect 8353 7044 8409 7100
rect 8409 7044 8413 7100
rect 8349 7040 8413 7044
rect 8429 7100 8493 7104
rect 8429 7044 8433 7100
rect 8433 7044 8489 7100
rect 8489 7044 8493 7100
rect 8429 7040 8493 7044
rect 6868 7032 6932 7036
rect 6868 6976 6882 7032
rect 6882 6976 6932 7032
rect 6868 6972 6932 6976
rect 2761 6556 2825 6560
rect 2761 6500 2765 6556
rect 2765 6500 2821 6556
rect 2821 6500 2825 6556
rect 2761 6496 2825 6500
rect 2841 6556 2905 6560
rect 2841 6500 2845 6556
rect 2845 6500 2901 6556
rect 2901 6500 2905 6556
rect 2841 6496 2905 6500
rect 2921 6556 2985 6560
rect 2921 6500 2925 6556
rect 2925 6500 2981 6556
rect 2981 6500 2985 6556
rect 2921 6496 2985 6500
rect 3001 6556 3065 6560
rect 3001 6500 3005 6556
rect 3005 6500 3061 6556
rect 3061 6500 3065 6556
rect 3001 6496 3065 6500
rect 6380 6556 6444 6560
rect 6380 6500 6384 6556
rect 6384 6500 6440 6556
rect 6440 6500 6444 6556
rect 6380 6496 6444 6500
rect 6460 6556 6524 6560
rect 6460 6500 6464 6556
rect 6464 6500 6520 6556
rect 6520 6500 6524 6556
rect 6460 6496 6524 6500
rect 6540 6556 6604 6560
rect 6540 6500 6544 6556
rect 6544 6500 6600 6556
rect 6600 6500 6604 6556
rect 6540 6496 6604 6500
rect 6620 6556 6684 6560
rect 6620 6500 6624 6556
rect 6624 6500 6680 6556
rect 6680 6500 6684 6556
rect 6620 6496 6684 6500
rect 9998 6556 10062 6560
rect 9998 6500 10002 6556
rect 10002 6500 10058 6556
rect 10058 6500 10062 6556
rect 9998 6496 10062 6500
rect 10078 6556 10142 6560
rect 10078 6500 10082 6556
rect 10082 6500 10138 6556
rect 10138 6500 10142 6556
rect 10078 6496 10142 6500
rect 10158 6556 10222 6560
rect 10158 6500 10162 6556
rect 10162 6500 10218 6556
rect 10218 6500 10222 6556
rect 10158 6496 10222 6500
rect 10238 6556 10302 6560
rect 10238 6500 10242 6556
rect 10242 6500 10298 6556
rect 10298 6500 10302 6556
rect 10238 6496 10302 6500
rect 6132 6080 6196 6084
rect 6132 6024 6182 6080
rect 6182 6024 6196 6080
rect 6132 6020 6196 6024
rect 6868 6020 6932 6084
rect 4570 6012 4634 6016
rect 4570 5956 4574 6012
rect 4574 5956 4630 6012
rect 4630 5956 4634 6012
rect 4570 5952 4634 5956
rect 4650 6012 4714 6016
rect 4650 5956 4654 6012
rect 4654 5956 4710 6012
rect 4710 5956 4714 6012
rect 4650 5952 4714 5956
rect 4730 6012 4794 6016
rect 4730 5956 4734 6012
rect 4734 5956 4790 6012
rect 4790 5956 4794 6012
rect 4730 5952 4794 5956
rect 4810 6012 4874 6016
rect 4810 5956 4814 6012
rect 4814 5956 4870 6012
rect 4870 5956 4874 6012
rect 4810 5952 4874 5956
rect 8189 6012 8253 6016
rect 8189 5956 8193 6012
rect 8193 5956 8249 6012
rect 8249 5956 8253 6012
rect 8189 5952 8253 5956
rect 8269 6012 8333 6016
rect 8269 5956 8273 6012
rect 8273 5956 8329 6012
rect 8329 5956 8333 6012
rect 8269 5952 8333 5956
rect 8349 6012 8413 6016
rect 8349 5956 8353 6012
rect 8353 5956 8409 6012
rect 8409 5956 8413 6012
rect 8349 5952 8413 5956
rect 8429 6012 8493 6016
rect 8429 5956 8433 6012
rect 8433 5956 8489 6012
rect 8489 5956 8493 6012
rect 8429 5952 8493 5956
rect 2761 5468 2825 5472
rect 2761 5412 2765 5468
rect 2765 5412 2821 5468
rect 2821 5412 2825 5468
rect 2761 5408 2825 5412
rect 2841 5468 2905 5472
rect 2841 5412 2845 5468
rect 2845 5412 2901 5468
rect 2901 5412 2905 5468
rect 2841 5408 2905 5412
rect 2921 5468 2985 5472
rect 2921 5412 2925 5468
rect 2925 5412 2981 5468
rect 2981 5412 2985 5468
rect 2921 5408 2985 5412
rect 3001 5468 3065 5472
rect 3001 5412 3005 5468
rect 3005 5412 3061 5468
rect 3061 5412 3065 5468
rect 3001 5408 3065 5412
rect 6380 5468 6444 5472
rect 6380 5412 6384 5468
rect 6384 5412 6440 5468
rect 6440 5412 6444 5468
rect 6380 5408 6444 5412
rect 6460 5468 6524 5472
rect 6460 5412 6464 5468
rect 6464 5412 6520 5468
rect 6520 5412 6524 5468
rect 6460 5408 6524 5412
rect 6540 5468 6604 5472
rect 6540 5412 6544 5468
rect 6544 5412 6600 5468
rect 6600 5412 6604 5468
rect 6540 5408 6604 5412
rect 6620 5468 6684 5472
rect 6620 5412 6624 5468
rect 6624 5412 6680 5468
rect 6680 5412 6684 5468
rect 6620 5408 6684 5412
rect 9998 5468 10062 5472
rect 9998 5412 10002 5468
rect 10002 5412 10058 5468
rect 10058 5412 10062 5468
rect 9998 5408 10062 5412
rect 10078 5468 10142 5472
rect 10078 5412 10082 5468
rect 10082 5412 10138 5468
rect 10138 5412 10142 5468
rect 10078 5408 10142 5412
rect 10158 5468 10222 5472
rect 10158 5412 10162 5468
rect 10162 5412 10218 5468
rect 10218 5412 10222 5468
rect 10158 5408 10222 5412
rect 10238 5468 10302 5472
rect 10238 5412 10242 5468
rect 10242 5412 10298 5468
rect 10298 5412 10302 5468
rect 10238 5408 10302 5412
rect 4570 4924 4634 4928
rect 4570 4868 4574 4924
rect 4574 4868 4630 4924
rect 4630 4868 4634 4924
rect 4570 4864 4634 4868
rect 4650 4924 4714 4928
rect 4650 4868 4654 4924
rect 4654 4868 4710 4924
rect 4710 4868 4714 4924
rect 4650 4864 4714 4868
rect 4730 4924 4794 4928
rect 4730 4868 4734 4924
rect 4734 4868 4790 4924
rect 4790 4868 4794 4924
rect 4730 4864 4794 4868
rect 4810 4924 4874 4928
rect 4810 4868 4814 4924
rect 4814 4868 4870 4924
rect 4870 4868 4874 4924
rect 4810 4864 4874 4868
rect 8189 4924 8253 4928
rect 8189 4868 8193 4924
rect 8193 4868 8249 4924
rect 8249 4868 8253 4924
rect 8189 4864 8253 4868
rect 8269 4924 8333 4928
rect 8269 4868 8273 4924
rect 8273 4868 8329 4924
rect 8329 4868 8333 4924
rect 8269 4864 8333 4868
rect 8349 4924 8413 4928
rect 8349 4868 8353 4924
rect 8353 4868 8409 4924
rect 8409 4868 8413 4924
rect 8349 4864 8413 4868
rect 8429 4924 8493 4928
rect 8429 4868 8433 4924
rect 8433 4868 8489 4924
rect 8489 4868 8493 4924
rect 8429 4864 8493 4868
rect 2761 4380 2825 4384
rect 2761 4324 2765 4380
rect 2765 4324 2821 4380
rect 2821 4324 2825 4380
rect 2761 4320 2825 4324
rect 2841 4380 2905 4384
rect 2841 4324 2845 4380
rect 2845 4324 2901 4380
rect 2901 4324 2905 4380
rect 2841 4320 2905 4324
rect 2921 4380 2985 4384
rect 2921 4324 2925 4380
rect 2925 4324 2981 4380
rect 2981 4324 2985 4380
rect 2921 4320 2985 4324
rect 3001 4380 3065 4384
rect 3001 4324 3005 4380
rect 3005 4324 3061 4380
rect 3061 4324 3065 4380
rect 3001 4320 3065 4324
rect 6380 4380 6444 4384
rect 6380 4324 6384 4380
rect 6384 4324 6440 4380
rect 6440 4324 6444 4380
rect 6380 4320 6444 4324
rect 6460 4380 6524 4384
rect 6460 4324 6464 4380
rect 6464 4324 6520 4380
rect 6520 4324 6524 4380
rect 6460 4320 6524 4324
rect 6540 4380 6604 4384
rect 6540 4324 6544 4380
rect 6544 4324 6600 4380
rect 6600 4324 6604 4380
rect 6540 4320 6604 4324
rect 6620 4380 6684 4384
rect 6620 4324 6624 4380
rect 6624 4324 6680 4380
rect 6680 4324 6684 4380
rect 6620 4320 6684 4324
rect 9998 4380 10062 4384
rect 9998 4324 10002 4380
rect 10002 4324 10058 4380
rect 10058 4324 10062 4380
rect 9998 4320 10062 4324
rect 10078 4380 10142 4384
rect 10078 4324 10082 4380
rect 10082 4324 10138 4380
rect 10138 4324 10142 4380
rect 10078 4320 10142 4324
rect 10158 4380 10222 4384
rect 10158 4324 10162 4380
rect 10162 4324 10218 4380
rect 10218 4324 10222 4380
rect 10158 4320 10222 4324
rect 10238 4380 10302 4384
rect 10238 4324 10242 4380
rect 10242 4324 10298 4380
rect 10298 4324 10302 4380
rect 10238 4320 10302 4324
rect 4570 3836 4634 3840
rect 4570 3780 4574 3836
rect 4574 3780 4630 3836
rect 4630 3780 4634 3836
rect 4570 3776 4634 3780
rect 4650 3836 4714 3840
rect 4650 3780 4654 3836
rect 4654 3780 4710 3836
rect 4710 3780 4714 3836
rect 4650 3776 4714 3780
rect 4730 3836 4794 3840
rect 4730 3780 4734 3836
rect 4734 3780 4790 3836
rect 4790 3780 4794 3836
rect 4730 3776 4794 3780
rect 4810 3836 4874 3840
rect 4810 3780 4814 3836
rect 4814 3780 4870 3836
rect 4870 3780 4874 3836
rect 4810 3776 4874 3780
rect 8189 3836 8253 3840
rect 8189 3780 8193 3836
rect 8193 3780 8249 3836
rect 8249 3780 8253 3836
rect 8189 3776 8253 3780
rect 8269 3836 8333 3840
rect 8269 3780 8273 3836
rect 8273 3780 8329 3836
rect 8329 3780 8333 3836
rect 8269 3776 8333 3780
rect 8349 3836 8413 3840
rect 8349 3780 8353 3836
rect 8353 3780 8409 3836
rect 8409 3780 8413 3836
rect 8349 3776 8413 3780
rect 8429 3836 8493 3840
rect 8429 3780 8433 3836
rect 8433 3780 8489 3836
rect 8489 3780 8493 3836
rect 8429 3776 8493 3780
rect 2761 3292 2825 3296
rect 2761 3236 2765 3292
rect 2765 3236 2821 3292
rect 2821 3236 2825 3292
rect 2761 3232 2825 3236
rect 2841 3292 2905 3296
rect 2841 3236 2845 3292
rect 2845 3236 2901 3292
rect 2901 3236 2905 3292
rect 2841 3232 2905 3236
rect 2921 3292 2985 3296
rect 2921 3236 2925 3292
rect 2925 3236 2981 3292
rect 2981 3236 2985 3292
rect 2921 3232 2985 3236
rect 3001 3292 3065 3296
rect 3001 3236 3005 3292
rect 3005 3236 3061 3292
rect 3061 3236 3065 3292
rect 3001 3232 3065 3236
rect 6380 3292 6444 3296
rect 6380 3236 6384 3292
rect 6384 3236 6440 3292
rect 6440 3236 6444 3292
rect 6380 3232 6444 3236
rect 6460 3292 6524 3296
rect 6460 3236 6464 3292
rect 6464 3236 6520 3292
rect 6520 3236 6524 3292
rect 6460 3232 6524 3236
rect 6540 3292 6604 3296
rect 6540 3236 6544 3292
rect 6544 3236 6600 3292
rect 6600 3236 6604 3292
rect 6540 3232 6604 3236
rect 6620 3292 6684 3296
rect 6620 3236 6624 3292
rect 6624 3236 6680 3292
rect 6680 3236 6684 3292
rect 6620 3232 6684 3236
rect 9998 3292 10062 3296
rect 9998 3236 10002 3292
rect 10002 3236 10058 3292
rect 10058 3236 10062 3292
rect 9998 3232 10062 3236
rect 10078 3292 10142 3296
rect 10078 3236 10082 3292
rect 10082 3236 10138 3292
rect 10138 3236 10142 3292
rect 10078 3232 10142 3236
rect 10158 3292 10222 3296
rect 10158 3236 10162 3292
rect 10162 3236 10218 3292
rect 10218 3236 10222 3292
rect 10158 3232 10222 3236
rect 10238 3292 10302 3296
rect 10238 3236 10242 3292
rect 10242 3236 10298 3292
rect 10298 3236 10302 3292
rect 10238 3232 10302 3236
rect 4570 2748 4634 2752
rect 4570 2692 4574 2748
rect 4574 2692 4630 2748
rect 4630 2692 4634 2748
rect 4570 2688 4634 2692
rect 4650 2748 4714 2752
rect 4650 2692 4654 2748
rect 4654 2692 4710 2748
rect 4710 2692 4714 2748
rect 4650 2688 4714 2692
rect 4730 2748 4794 2752
rect 4730 2692 4734 2748
rect 4734 2692 4790 2748
rect 4790 2692 4794 2748
rect 4730 2688 4794 2692
rect 4810 2748 4874 2752
rect 4810 2692 4814 2748
rect 4814 2692 4870 2748
rect 4870 2692 4874 2748
rect 4810 2688 4874 2692
rect 8189 2748 8253 2752
rect 8189 2692 8193 2748
rect 8193 2692 8249 2748
rect 8249 2692 8253 2748
rect 8189 2688 8253 2692
rect 8269 2748 8333 2752
rect 8269 2692 8273 2748
rect 8273 2692 8329 2748
rect 8329 2692 8333 2748
rect 8269 2688 8333 2692
rect 8349 2748 8413 2752
rect 8349 2692 8353 2748
rect 8353 2692 8409 2748
rect 8409 2692 8413 2748
rect 8349 2688 8413 2692
rect 8429 2748 8493 2752
rect 8429 2692 8433 2748
rect 8433 2692 8489 2748
rect 8489 2692 8493 2748
rect 8429 2688 8493 2692
rect 2761 2204 2825 2208
rect 2761 2148 2765 2204
rect 2765 2148 2821 2204
rect 2821 2148 2825 2204
rect 2761 2144 2825 2148
rect 2841 2204 2905 2208
rect 2841 2148 2845 2204
rect 2845 2148 2901 2204
rect 2901 2148 2905 2204
rect 2841 2144 2905 2148
rect 2921 2204 2985 2208
rect 2921 2148 2925 2204
rect 2925 2148 2981 2204
rect 2981 2148 2985 2204
rect 2921 2144 2985 2148
rect 3001 2204 3065 2208
rect 3001 2148 3005 2204
rect 3005 2148 3061 2204
rect 3061 2148 3065 2204
rect 3001 2144 3065 2148
rect 6380 2204 6444 2208
rect 6380 2148 6384 2204
rect 6384 2148 6440 2204
rect 6440 2148 6444 2204
rect 6380 2144 6444 2148
rect 6460 2204 6524 2208
rect 6460 2148 6464 2204
rect 6464 2148 6520 2204
rect 6520 2148 6524 2204
rect 6460 2144 6524 2148
rect 6540 2204 6604 2208
rect 6540 2148 6544 2204
rect 6544 2148 6600 2204
rect 6600 2148 6604 2204
rect 6540 2144 6604 2148
rect 6620 2204 6684 2208
rect 6620 2148 6624 2204
rect 6624 2148 6680 2204
rect 6680 2148 6684 2204
rect 6620 2144 6684 2148
rect 9998 2204 10062 2208
rect 9998 2148 10002 2204
rect 10002 2148 10058 2204
rect 10058 2148 10062 2204
rect 9998 2144 10062 2148
rect 10078 2204 10142 2208
rect 10078 2148 10082 2204
rect 10082 2148 10138 2204
rect 10138 2148 10142 2204
rect 10078 2144 10142 2148
rect 10158 2204 10222 2208
rect 10158 2148 10162 2204
rect 10162 2148 10218 2204
rect 10218 2148 10222 2204
rect 10158 2144 10222 2148
rect 10238 2204 10302 2208
rect 10238 2148 10242 2204
rect 10242 2148 10298 2204
rect 10298 2148 10302 2204
rect 10238 2144 10302 2148
<< metal4 >>
rect 2753 13088 3073 13104
rect 2753 13024 2761 13088
rect 2825 13024 2841 13088
rect 2905 13024 2921 13088
rect 2985 13024 3001 13088
rect 3065 13024 3073 13088
rect 2753 12000 3073 13024
rect 2753 11936 2761 12000
rect 2825 11936 2841 12000
rect 2905 11936 2921 12000
rect 2985 11936 3001 12000
rect 3065 11936 3073 12000
rect 2753 10912 3073 11936
rect 2753 10848 2761 10912
rect 2825 10848 2841 10912
rect 2905 10848 2921 10912
rect 2985 10848 3001 10912
rect 3065 10848 3073 10912
rect 2753 9824 3073 10848
rect 2753 9760 2761 9824
rect 2825 9760 2841 9824
rect 2905 9760 2921 9824
rect 2985 9760 3001 9824
rect 3065 9760 3073 9824
rect 2753 8736 3073 9760
rect 2753 8672 2761 8736
rect 2825 8672 2841 8736
rect 2905 8672 2921 8736
rect 2985 8672 3001 8736
rect 3065 8672 3073 8736
rect 2753 7648 3073 8672
rect 2753 7584 2761 7648
rect 2825 7584 2841 7648
rect 2905 7584 2921 7648
rect 2985 7584 3001 7648
rect 3065 7584 3073 7648
rect 2753 6560 3073 7584
rect 2753 6496 2761 6560
rect 2825 6496 2841 6560
rect 2905 6496 2921 6560
rect 2985 6496 3001 6560
rect 3065 6496 3073 6560
rect 2753 5472 3073 6496
rect 2753 5408 2761 5472
rect 2825 5408 2841 5472
rect 2905 5408 2921 5472
rect 2985 5408 3001 5472
rect 3065 5408 3073 5472
rect 2753 4384 3073 5408
rect 2753 4320 2761 4384
rect 2825 4320 2841 4384
rect 2905 4320 2921 4384
rect 2985 4320 3001 4384
rect 3065 4320 3073 4384
rect 2753 3296 3073 4320
rect 2753 3232 2761 3296
rect 2825 3232 2841 3296
rect 2905 3232 2921 3296
rect 2985 3232 3001 3296
rect 3065 3232 3073 3296
rect 2753 2208 3073 3232
rect 2753 2144 2761 2208
rect 2825 2144 2841 2208
rect 2905 2144 2921 2208
rect 2985 2144 3001 2208
rect 3065 2144 3073 2208
rect 2753 2128 3073 2144
rect 4562 12544 4883 13104
rect 4562 12480 4570 12544
rect 4634 12480 4650 12544
rect 4714 12480 4730 12544
rect 4794 12480 4810 12544
rect 4874 12480 4883 12544
rect 4562 11456 4883 12480
rect 4562 11392 4570 11456
rect 4634 11392 4650 11456
rect 4714 11392 4730 11456
rect 4794 11392 4810 11456
rect 4874 11392 4883 11456
rect 4562 10368 4883 11392
rect 4562 10304 4570 10368
rect 4634 10304 4650 10368
rect 4714 10304 4730 10368
rect 4794 10304 4810 10368
rect 4874 10304 4883 10368
rect 4562 9280 4883 10304
rect 4562 9216 4570 9280
rect 4634 9216 4650 9280
rect 4714 9216 4730 9280
rect 4794 9216 4810 9280
rect 4874 9216 4883 9280
rect 4562 8192 4883 9216
rect 6372 13088 6692 13104
rect 6372 13024 6380 13088
rect 6444 13024 6460 13088
rect 6524 13024 6540 13088
rect 6604 13024 6620 13088
rect 6684 13024 6692 13088
rect 6372 12000 6692 13024
rect 6372 11936 6380 12000
rect 6444 11936 6460 12000
rect 6524 11936 6540 12000
rect 6604 11936 6620 12000
rect 6684 11936 6692 12000
rect 6372 10912 6692 11936
rect 6372 10848 6380 10912
rect 6444 10848 6460 10912
rect 6524 10848 6540 10912
rect 6604 10848 6620 10912
rect 6684 10848 6692 10912
rect 6372 9824 6692 10848
rect 6372 9760 6380 9824
rect 6444 9760 6460 9824
rect 6524 9760 6540 9824
rect 6604 9760 6620 9824
rect 6684 9760 6692 9824
rect 6131 8940 6197 8941
rect 6131 8876 6132 8940
rect 6196 8876 6197 8940
rect 6131 8875 6197 8876
rect 4562 8128 4570 8192
rect 4634 8128 4650 8192
rect 4714 8128 4730 8192
rect 4794 8128 4810 8192
rect 4874 8128 4883 8192
rect 4562 7104 4883 8128
rect 4562 7040 4570 7104
rect 4634 7040 4650 7104
rect 4714 7040 4730 7104
rect 4794 7040 4810 7104
rect 4874 7040 4883 7104
rect 4562 6016 4883 7040
rect 6134 6085 6194 8875
rect 6372 8736 6692 9760
rect 6372 8672 6380 8736
rect 6444 8672 6460 8736
rect 6524 8672 6540 8736
rect 6604 8672 6620 8736
rect 6684 8672 6692 8736
rect 6372 7648 6692 8672
rect 6372 7584 6380 7648
rect 6444 7584 6460 7648
rect 6524 7584 6540 7648
rect 6604 7584 6620 7648
rect 6684 7584 6692 7648
rect 6372 6560 6692 7584
rect 8181 12544 8501 13104
rect 8181 12480 8189 12544
rect 8253 12480 8269 12544
rect 8333 12480 8349 12544
rect 8413 12480 8429 12544
rect 8493 12480 8501 12544
rect 8181 11456 8501 12480
rect 8181 11392 8189 11456
rect 8253 11392 8269 11456
rect 8333 11392 8349 11456
rect 8413 11392 8429 11456
rect 8493 11392 8501 11456
rect 8181 10368 8501 11392
rect 8181 10304 8189 10368
rect 8253 10304 8269 10368
rect 8333 10304 8349 10368
rect 8413 10304 8429 10368
rect 8493 10304 8501 10368
rect 8181 9280 8501 10304
rect 8181 9216 8189 9280
rect 8253 9216 8269 9280
rect 8333 9216 8349 9280
rect 8413 9216 8429 9280
rect 8493 9216 8501 9280
rect 8181 8192 8501 9216
rect 8181 8128 8189 8192
rect 8253 8128 8269 8192
rect 8333 8128 8349 8192
rect 8413 8128 8429 8192
rect 8493 8128 8501 8192
rect 8181 7104 8501 8128
rect 8181 7040 8189 7104
rect 8253 7040 8269 7104
rect 8333 7040 8349 7104
rect 8413 7040 8429 7104
rect 8493 7040 8501 7104
rect 6867 7036 6933 7037
rect 6867 6972 6868 7036
rect 6932 6972 6933 7036
rect 6867 6971 6933 6972
rect 6372 6496 6380 6560
rect 6444 6496 6460 6560
rect 6524 6496 6540 6560
rect 6604 6496 6620 6560
rect 6684 6496 6692 6560
rect 6131 6084 6197 6085
rect 6131 6020 6132 6084
rect 6196 6020 6197 6084
rect 6131 6019 6197 6020
rect 4562 5952 4570 6016
rect 4634 5952 4650 6016
rect 4714 5952 4730 6016
rect 4794 5952 4810 6016
rect 4874 5952 4883 6016
rect 4562 4928 4883 5952
rect 4562 4864 4570 4928
rect 4634 4864 4650 4928
rect 4714 4864 4730 4928
rect 4794 4864 4810 4928
rect 4874 4864 4883 4928
rect 4562 3840 4883 4864
rect 4562 3776 4570 3840
rect 4634 3776 4650 3840
rect 4714 3776 4730 3840
rect 4794 3776 4810 3840
rect 4874 3776 4883 3840
rect 4562 2752 4883 3776
rect 4562 2688 4570 2752
rect 4634 2688 4650 2752
rect 4714 2688 4730 2752
rect 4794 2688 4810 2752
rect 4874 2688 4883 2752
rect 4562 2128 4883 2688
rect 6372 5472 6692 6496
rect 6870 6085 6930 6971
rect 6867 6084 6933 6085
rect 6867 6020 6868 6084
rect 6932 6020 6933 6084
rect 6867 6019 6933 6020
rect 6372 5408 6380 5472
rect 6444 5408 6460 5472
rect 6524 5408 6540 5472
rect 6604 5408 6620 5472
rect 6684 5408 6692 5472
rect 6372 4384 6692 5408
rect 6372 4320 6380 4384
rect 6444 4320 6460 4384
rect 6524 4320 6540 4384
rect 6604 4320 6620 4384
rect 6684 4320 6692 4384
rect 6372 3296 6692 4320
rect 6372 3232 6380 3296
rect 6444 3232 6460 3296
rect 6524 3232 6540 3296
rect 6604 3232 6620 3296
rect 6684 3232 6692 3296
rect 6372 2208 6692 3232
rect 6372 2144 6380 2208
rect 6444 2144 6460 2208
rect 6524 2144 6540 2208
rect 6604 2144 6620 2208
rect 6684 2144 6692 2208
rect 6372 2128 6692 2144
rect 8181 6016 8501 7040
rect 8181 5952 8189 6016
rect 8253 5952 8269 6016
rect 8333 5952 8349 6016
rect 8413 5952 8429 6016
rect 8493 5952 8501 6016
rect 8181 4928 8501 5952
rect 8181 4864 8189 4928
rect 8253 4864 8269 4928
rect 8333 4864 8349 4928
rect 8413 4864 8429 4928
rect 8493 4864 8501 4928
rect 8181 3840 8501 4864
rect 8181 3776 8189 3840
rect 8253 3776 8269 3840
rect 8333 3776 8349 3840
rect 8413 3776 8429 3840
rect 8493 3776 8501 3840
rect 8181 2752 8501 3776
rect 8181 2688 8189 2752
rect 8253 2688 8269 2752
rect 8333 2688 8349 2752
rect 8413 2688 8429 2752
rect 8493 2688 8501 2752
rect 8181 2128 8501 2688
rect 9990 13088 10311 13104
rect 9990 13024 9998 13088
rect 10062 13024 10078 13088
rect 10142 13024 10158 13088
rect 10222 13024 10238 13088
rect 10302 13024 10311 13088
rect 9990 12000 10311 13024
rect 9990 11936 9998 12000
rect 10062 11936 10078 12000
rect 10142 11936 10158 12000
rect 10222 11936 10238 12000
rect 10302 11936 10311 12000
rect 9990 10912 10311 11936
rect 9990 10848 9998 10912
rect 10062 10848 10078 10912
rect 10142 10848 10158 10912
rect 10222 10848 10238 10912
rect 10302 10848 10311 10912
rect 9990 9824 10311 10848
rect 9990 9760 9998 9824
rect 10062 9760 10078 9824
rect 10142 9760 10158 9824
rect 10222 9760 10238 9824
rect 10302 9760 10311 9824
rect 9990 8736 10311 9760
rect 9990 8672 9998 8736
rect 10062 8672 10078 8736
rect 10142 8672 10158 8736
rect 10222 8672 10238 8736
rect 10302 8672 10311 8736
rect 9990 7648 10311 8672
rect 9990 7584 9998 7648
rect 10062 7584 10078 7648
rect 10142 7584 10158 7648
rect 10222 7584 10238 7648
rect 10302 7584 10311 7648
rect 9990 6560 10311 7584
rect 9990 6496 9998 6560
rect 10062 6496 10078 6560
rect 10142 6496 10158 6560
rect 10222 6496 10238 6560
rect 10302 6496 10311 6560
rect 9990 5472 10311 6496
rect 9990 5408 9998 5472
rect 10062 5408 10078 5472
rect 10142 5408 10158 5472
rect 10222 5408 10238 5472
rect 10302 5408 10311 5472
rect 9990 4384 10311 5408
rect 9990 4320 9998 4384
rect 10062 4320 10078 4384
rect 10142 4320 10158 4384
rect 10222 4320 10238 4384
rect 10302 4320 10311 4384
rect 9990 3296 10311 4320
rect 9990 3232 9998 3296
rect 10062 3232 10078 3296
rect 10142 3232 10158 3296
rect 10222 3232 10238 3296
rect 10302 3232 10311 3296
rect 9990 2208 10311 3232
rect 9990 2144 9998 2208
rect 10062 2144 10078 2208
rect 10142 2144 10158 2208
rect 10222 2144 10238 2208
rect 10302 2144 10311 2208
rect 9990 2128 10311 2144
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1608164981
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608164981
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608164981
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608164981
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608164981
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608164981
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608164981
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608164981
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_62
timestamp 1608164981
transform 1 0 6808 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1608164981
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1608164981
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6992 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp 1608164981
transform 1 0 7544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_75
timestamp 1608164981
transform 1 0 8004 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_79
timestamp 1608164981
transform 1 0 8372 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_67
timestamp 1608164981
transform 1 0 7268 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_99
timestamp 1608164981
transform 1 0 10212 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_87
timestamp 1608164981
transform 1 0 9108 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1608164981
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1608164981
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1608164981
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_111
timestamp 1608164981
transform 1 0 11316 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_114
timestamp 1608164981
transform 1 0 11592 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106
timestamp 1608164981
transform 1 0 10856 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608164981
transform -1 0 11960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608164981
transform -1 0 11960 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_18
timestamp 1608164981
transform 1 0 2760 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_13
timestamp 1608164981
transform 1 0 2300 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_7
timestamp 1608164981
transform 1 0 1748 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608164981
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _160_
timestamp 1608164981
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _158_
timestamp 1608164981
transform 1 0 2392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1608164981
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1608164981
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1608164981
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1608164981
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1608164981
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1608164981
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1608164981
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1608164981
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1608164981
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1608164981
transform 1 0 11500 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_105
timestamp 1608164981
transform 1 0 10764 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608164981
transform -1 0 11960 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1608164981
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608164981
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608164981
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1608164981
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1608164981
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1608164981
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1608164981
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1608164981
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_65
timestamp 1608164981
transform 1 0 7084 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1608164981
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1608164981
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8188 0 1 3808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_3_91
timestamp 1608164981
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_103
timestamp 1608164981
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608164981
transform -1 0 11960 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608164981
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608164981
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608164981
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608164981
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608164981
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608164981
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_44
timestamp 1608164981
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1608164981
transform 1 0 5336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1608164981
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6164 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1608164981
transform 1 0 5888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_73
timestamp 1608164981
transform 1 0 7820 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8372 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _077_
timestamp 1608164981
transform 1 0 6992 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1608164981
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608164981
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 1608164981
transform 1 0 9016 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_109
timestamp 1608164981
transform 1 0 11132 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608164981
transform -1 0 11960 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608164981
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608164981
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608164981
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608164981
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_4  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 4692 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_5_44
timestamp 1608164981
transform 1 0 5152 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 5244 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _101_
timestamp 1608164981
transform 1 0 6072 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608164981
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _147_
timestamp 1608164981
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _079_
timestamp 1608164981
transform 1 0 7636 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_92
timestamp 1608164981
transform 1 0 9568 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1608164981
transform 1 0 8464 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_112
timestamp 1608164981
transform 1 0 11408 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1608164981
transform 1 0 10672 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608164981
transform -1 0 11960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1608164981
transform 1 0 2484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608164981
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608164981
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608164981
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608164981
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608164981
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1608164981
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1608164981
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608164981
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608164981
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 4508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 3680 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _127_
timestamp 1608164981
transform 1 0 4232 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1608164981
transform 1 0 3404 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1608164981
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _149_
timestamp 1608164981
transform 1 0 5060 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _142_
timestamp 1608164981
transform 1 0 6164 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_4  _089_
timestamp 1608164981
transform 1 0 5612 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608164981
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _150_
timestamp 1608164981
transform 1 0 7452 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _132_
timestamp 1608164981
transform 1 0 8280 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__a32o_4  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 6808 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_4  _090_
timestamp 1608164981
transform 1 0 8372 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_6_96
timestamp 1608164981
transform 1 0 9936 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608164981
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__a22oi_4  _125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 8832 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1608164981
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1608164981
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_101
timestamp 1608164981
transform 1 0 10396 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_114
timestamp 1608164981
transform 1 0 11592 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_108
timestamp 1608164981
transform 1 0 11040 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608164981
transform -1 0 11960 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608164981
transform -1 0 11960 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608164981
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608164981
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _119_
timestamp 1608164981
transform 1 0 2484 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1608164981
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608164981
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 4232 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 3128 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_4  _096_
timestamp 1608164981
transform 1 0 5980 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__a32o_4  _145_
timestamp 1608164981
transform 1 0 7544 0 -1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1608164981
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608164981
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _144_
timestamp 1608164981
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1608164981
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_109
timestamp 1608164981
transform 1 0 11132 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608164981
transform -1 0 11960 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _117_
timestamp 1608164981
transform 1 0 10488 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1608164981
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608164981
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _100_
timestamp 1608164981
transform 1 0 2208 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1608164981
transform 1 0 1656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1608164981
transform 1 0 1932 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _140_
timestamp 1608164981
transform 1 0 3036 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _115_
timestamp 1608164981
transform 1 0 3864 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__a32o_4  _120_
timestamp 1608164981
transform 1 0 5152 0 1 7072
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608164981
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _141_
timestamp 1608164981
transform 1 0 6808 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__o22a_4  _081_
timestamp 1608164981
transform 1 0 8096 0 1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_4  _153_
timestamp 1608164981
transform 1 0 9384 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_114
timestamp 1608164981
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608164981
transform -1 0 11960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1608164981
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _138_
timestamp 1608164981
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1608164981
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1608164981
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608164981
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1608164981
transform 1 0 2300 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _129_
timestamp 1608164981
transform 1 0 2576 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1608164981
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608164981
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _114_
timestamp 1608164981
transform 1 0 4692 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _071_
timestamp 1608164981
transform 1 0 4048 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_4  _083_
timestamp 1608164981
transform 1 0 5796 0 -1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__a2bb2o_4  _123_
timestamp 1608164981
transform 1 0 7360 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1608164981
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608164981
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _157_
timestamp 1608164981
transform 1 0 8832 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _110_
timestamp 1608164981
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_112
timestamp 1608164981
transform 1 0 11408 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608164981
transform -1 0 11960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _159_
timestamp 1608164981
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 1608164981
transform 1 0 11132 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1608164981
transform 1 0 10856 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1608164981
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608164981
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608164981
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _084_
timestamp 1608164981
transform 1 0 2852 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _163_
timestamp 1608164981
transform 1 0 4324 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__nor2_4  _070_
timestamp 1608164981
transform 1 0 3496 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _137_
timestamp 1608164981
transform 1 0 6072 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608164981
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _131_
timestamp 1608164981
transform 1 0 6808 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_4  _080_
timestamp 1608164981
transform 1 0 8372 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__or4_4  _093_
timestamp 1608164981
transform 1 0 9660 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1608164981
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_105
timestamp 1608164981
transform 1 0 10764 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608164981
transform -1 0 11960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp 1608164981
transform 1 0 10488 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_15
timestamp 1608164981
transform 1 0 2484 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608164981
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608164981
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_25
timestamp 1608164981
transform 1 0 3404 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_21
timestamp 1608164981
transform 1 0 3036 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608164981
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _133_
timestamp 1608164981
transform 1 0 4600 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1608164981
transform 1 0 3128 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_4  _095_
timestamp 1608164981
transform 1 0 5704 0 -1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__o22a_4  _124_
timestamp 1608164981
transform 1 0 7268 0 -1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1608164981
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1608164981
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608164981
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _082_
timestamp 1608164981
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_113
timestamp 1608164981
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_105
timestamp 1608164981
transform 1 0 10764 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608164981
transform -1 0 11960 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608164981
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608164981
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_12
timestamp 1608164981
transform 1 0 2208 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 1608164981
transform 1 0 1380 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608164981
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608164981
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1608164981
transform 1 0 1932 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608164981
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608164981
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_39
timestamp 1608164981
transform 1 0 4692 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_32
timestamp 1608164981
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_24
timestamp 1608164981
transform 1 0 3312 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608164981
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _130_
timestamp 1608164981
transform 1 0 4232 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_4  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608164981
transform 1 0 3404 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_14_44
timestamp 1608164981
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _155_
timestamp 1608164981
transform 1 0 4784 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _111_
timestamp 1608164981
transform 1 0 5612 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _109_
timestamp 1608164981
transform 1 0 5888 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1608164981
transform 1 0 5612 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1608164981
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_79
timestamp 1608164981
transform 1 0 8372 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608164981
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _152_
timestamp 1608164981
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _134_
timestamp 1608164981
transform 1 0 6992 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _107_
timestamp 1608164981
transform 1 0 7912 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1608164981
transform 1 0 7820 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1608164981
transform 1 0 8096 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1608164981
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1608164981
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1608164981
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1608164981
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608164981
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1608164981
transform 1 0 8740 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_113
timestamp 1608164981
transform 1 0 11500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_105
timestamp 1608164981
transform 1 0 10764 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_114
timestamp 1608164981
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1608164981
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608164981
transform -1 0 11960 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608164981
transform -1 0 11960 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608164981
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608164981
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608164981
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1608164981
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1608164981
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_55
timestamp 1608164981
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_51
timestamp 1608164981
transform 1 0 5796 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1608164981
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp 1608164981
transform 1 0 6348 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_72
timestamp 1608164981
transform 1 0 7728 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1608164981
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608164981
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _102_
timestamp 1608164981
transform 1 0 6808 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp 1608164981
transform 1 0 7452 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_96
timestamp 1608164981
transform 1 0 9936 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_84
timestamp 1608164981
transform 1 0 8832 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_114
timestamp 1608164981
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_108
timestamp 1608164981
transform 1 0 11040 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608164981
transform -1 0 11960 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608164981
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608164981
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608164981
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608164981
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608164981
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608164981
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1608164981
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1608164981
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1608164981
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1608164981
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1608164981
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608164981
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_113
timestamp 1608164981
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_105
timestamp 1608164981
transform 1 0 10764 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608164981
transform -1 0 11960 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1608164981
transform 1 0 2484 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1608164981
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608164981
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_23
timestamp 1608164981
transform 1 0 3220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _162_
timestamp 1608164981
transform 1 0 3404 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1608164981
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1608164981
transform 1 0 5152 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1608164981
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1608164981
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1608164981
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608164981
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1608164981
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1608164981
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_114
timestamp 1608164981
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_110
timestamp 1608164981
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608164981
transform -1 0 11960 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608164981
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608164981
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608164981
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608164981
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1608164981
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608164981
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1608164981
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1608164981
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1608164981
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1608164981
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1608164981
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608164981
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_113
timestamp 1608164981
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_105
timestamp 1608164981
transform 1 0 10764 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608164981
transform -1 0 11960 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608164981
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608164981
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608164981
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1608164981
transform 1 0 4048 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1608164981
transform 1 0 3588 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608164981
transform 1 0 3956 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_56
timestamp 1608164981
transform 1 0 6256 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1608164981
transform 1 0 5152 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1608164981
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_63
timestamp 1608164981
transform 1 0 6900 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608164981
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1608164981
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1608164981
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_92
timestamp 1608164981
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_86
timestamp 1608164981
transform 1 0 9016 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608164981
transform 1 0 9660 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_114
timestamp 1608164981
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1608164981
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608164981
transform -1 0 11960 0 1 12512
box -38 -48 314 592
<< labels >>
rlabel metal2 s 3514 14440 3570 15240 6 cbitin
port 0 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 cbitout
port 1 nsew signal tristate
rlabel metal2 s 2042 14440 2098 15240 6 confclk
port 2 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 confclko
port 3 nsew signal tristate
rlabel metal2 s 9310 0 9366 800 6 dempty
port 4 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 din[0]
port 5 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 din[1]
port 6 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 dout[0]
port 7 nsew signal tristate
rlabel metal2 s 4986 0 5042 800 6 dout[1]
port 8 nsew signal tristate
rlabel metal3 s 0 6264 800 6384 6 hempty
port 9 nsew signal tristate
rlabel metal3 s 12296 8848 13096 8968 6 hempty2
port 10 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 lempty
port 11 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 lin[0]
port 12 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 lin[1]
port 13 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 lout[0]
port 14 nsew signal tristate
rlabel metal3 s 0 1232 800 1352 6 lout[1]
port 15 nsew signal tristate
rlabel metal3 s 12296 6264 13096 6384 6 rempty
port 16 nsew signal input
rlabel metal2 s 662 14440 718 15240 6 reset
port 17 nsew signal input
rlabel metal2 s 662 0 718 800 6 reseto
port 18 nsew signal tristate
rlabel metal3 s 12296 3680 13096 3800 6 rin[0]
port 19 nsew signal input
rlabel metal3 s 12296 1232 13096 1352 6 rin[1]
port 20 nsew signal input
rlabel metal3 s 12296 13880 13096 14000 6 rout[0]
port 21 nsew signal tristate
rlabel metal3 s 12296 11296 13096 11416 6 rout[1]
port 22 nsew signal tristate
rlabel metal2 s 7838 14440 7894 15240 6 uempty
port 23 nsew signal input
rlabel metal2 s 6458 14440 6514 15240 6 uin[0]
port 24 nsew signal input
rlabel metal2 s 4986 14440 5042 15240 6 uin[1]
port 25 nsew signal input
rlabel metal2 s 12254 14440 12310 15240 6 uout[0]
port 26 nsew signal tristate
rlabel metal2 s 10782 14440 10838 15240 6 uout[1]
port 27 nsew signal tristate
rlabel metal2 s 9310 14440 9366 15240 6 vempty
port 28 nsew signal tristate
rlabel metal2 s 7838 0 7894 800 6 vempty2
port 29 nsew signal tristate
rlabel metal4 s 9991 2128 10311 13104 6 vccd1
port 30 nsew power bidirectional
rlabel metal4 s 6372 2128 6692 13104 6 vccd1
port 31 nsew power bidirectional
rlabel metal4 s 2753 2128 3073 13104 6 vccd1
port 32 nsew power bidirectional
rlabel metal4 s 8181 2128 8501 13104 6 vssd1
port 33 nsew ground bidirectional
rlabel metal4 s 4563 2128 4883 13104 6 vssd1
port 34 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 13096 15240
<< end >>
