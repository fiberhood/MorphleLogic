// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

/* Generated by Yosys 0.9+3621 (git sha1 84e9fa7, gcc 8.3.1 -fPIC -Os) */

module mprj_logic_high(vccd1, vssd1, HI);
  output [458:0] HI;
  input vccd1;
  input vssd1;
  sky130_fd_sc_hd__fill_2 FILLER_0_102 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_113 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_117 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_122 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_143 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_147 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_162 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_172 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_176 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_195 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_215 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_226 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_233 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_237 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_242 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_246 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_277 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_292 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_0_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_305 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_309 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_317 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_327 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_334 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_345 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_349 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_362 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_384 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_407 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_41 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_414 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_421 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_432 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_435 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_442 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_446 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_450 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_455 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_463 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_466 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_485 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_49 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_500 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_507 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_528 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_536 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_0_549 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_56 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_568 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_575 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_585 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_60 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_617 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_66 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_73 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_0_92 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_0_94 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_103 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_107 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_115 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_119 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_138 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_145 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_157 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_169 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_173 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_181 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_190 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_202 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_210 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_235 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_242 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_245 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_275 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_287 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_292 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_304 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_306 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_314 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_318 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_322 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_326 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_338 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_350 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_356 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_364 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_367 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_379 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_391 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_400 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_412 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_417 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_425 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_428 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_435 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_443 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_448 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_457 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_469 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_475 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_479 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_487 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_489 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_49 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_501 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_509 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_525 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_531 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_1_543 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_550 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_562 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_1_574 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_583 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_588 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_608 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_1_614 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_618 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_1_62 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_1_70 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_75 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_1_87 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_1_99 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_105 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_109 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_121 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_130 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_142 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_15 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_150 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_154 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_166 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_171 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_183 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_194 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_198 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_206 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_218 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_222 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_227 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_235 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_240 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_247 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_259 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_264 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_269 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_273 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_285 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_292 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_302 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_322 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_330 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_334 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_343 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_353 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_361 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_368 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_374 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_378 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_390 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_396 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_398 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_402 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_406 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_41 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_418 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_433 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_444 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_456 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_459 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_2_467 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_472 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_479 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_491 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_500 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_504 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_508 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_516 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_53 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_535 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_544 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_556 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_567 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_579 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_2_608 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_2_616 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_65 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_2_77 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_83 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_2_87 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_2_91 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_2_93 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_103 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_107 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_111 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_128 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_132 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_139 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_159 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_173 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_180 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_184 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_196 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_200 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_207 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_221 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_240 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_247 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_252 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_260 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_12 FILLER_3_266 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_278 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_280 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_288 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_30 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_8 FILLER_3_300 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_308 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_311 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_317 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_32 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_6 FILLER_3_321 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_327 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_340 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 FILLER_3_354 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_363 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_37 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_371 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_385 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_392 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_419 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_423 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_427 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_435 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_44 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_443 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_447 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_457 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_475 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_483 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_494 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_497 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_505 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_513 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_520 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_534 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_542 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_546 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_553 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_557 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_565 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_570 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_583 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_587 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_60 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_4 FILLER_3_614 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_618 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_2 FILLER_3_69 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__fill_1 FILLER_3_89 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_0 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_1 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_18 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_19 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_2 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_20 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_21 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_22 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_23 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_24 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_25 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_26 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_27 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_28 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_29 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_3 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_30 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_31 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_32 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_33 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_34 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_35 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_36 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_37 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_38 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_39 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_4 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_40 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_41 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_42 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_43 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_44 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_45 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_46 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_47 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_48 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_49 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_5 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_50 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_51 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_52 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_53 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_54 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_55 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_56 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_57 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_58 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_59 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_6 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_60 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_61 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_62 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_63 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_64 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_65 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__decap_3 PHY_7 (
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9 (
    .VGND(vssd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[0]  (
    .HI(HI[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[100]  (
    .HI(HI[100]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[101]  (
    .HI(HI[101]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[102]  (
    .HI(HI[102]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[103]  (
    .HI(HI[103]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[104]  (
    .HI(HI[104]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[105]  (
    .HI(HI[105]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[106]  (
    .HI(HI[106]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[107]  (
    .HI(HI[107]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[108]  (
    .HI(HI[108]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[109]  (
    .HI(HI[109]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[10]  (
    .HI(HI[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[110]  (
    .HI(HI[110]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[111]  (
    .HI(HI[111]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[112]  (
    .HI(HI[112]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[113]  (
    .HI(HI[113]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[114]  (
    .HI(HI[114]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[115]  (
    .HI(HI[115]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[116]  (
    .HI(HI[116]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[117]  (
    .HI(HI[117]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[118]  (
    .HI(HI[118]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[119]  (
    .HI(HI[119]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[11]  (
    .HI(HI[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[120]  (
    .HI(HI[120]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[121]  (
    .HI(HI[121]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[122]  (
    .HI(HI[122]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[123]  (
    .HI(HI[123]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[124]  (
    .HI(HI[124]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[125]  (
    .HI(HI[125]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[126]  (
    .HI(HI[126]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[127]  (
    .HI(HI[127]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[128]  (
    .HI(HI[128]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[129]  (
    .HI(HI[129]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[12]  (
    .HI(HI[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[130]  (
    .HI(HI[130]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[131]  (
    .HI(HI[131]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[132]  (
    .HI(HI[132]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[133]  (
    .HI(HI[133]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[134]  (
    .HI(HI[134]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[135]  (
    .HI(HI[135]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[136]  (
    .HI(HI[136]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[137]  (
    .HI(HI[137]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[138]  (
    .HI(HI[138]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[139]  (
    .HI(HI[139]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[13]  (
    .HI(HI[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[140]  (
    .HI(HI[140]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[141]  (
    .HI(HI[141]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[142]  (
    .HI(HI[142]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[143]  (
    .HI(HI[143]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[144]  (
    .HI(HI[144]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[145]  (
    .HI(HI[145]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[146]  (
    .HI(HI[146]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[147]  (
    .HI(HI[147]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[148]  (
    .HI(HI[148]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[149]  (
    .HI(HI[149]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[14]  (
    .HI(HI[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[150]  (
    .HI(HI[150]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[151]  (
    .HI(HI[151]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[152]  (
    .HI(HI[152]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[153]  (
    .HI(HI[153]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[154]  (
    .HI(HI[154]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[155]  (
    .HI(HI[155]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[156]  (
    .HI(HI[156]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[157]  (
    .HI(HI[157]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[158]  (
    .HI(HI[158]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[159]  (
    .HI(HI[159]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[15]  (
    .HI(HI[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[160]  (
    .HI(HI[160]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[161]  (
    .HI(HI[161]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[162]  (
    .HI(HI[162]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[163]  (
    .HI(HI[163]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[164]  (
    .HI(HI[164]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[165]  (
    .HI(HI[165]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[166]  (
    .HI(HI[166]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[167]  (
    .HI(HI[167]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[168]  (
    .HI(HI[168]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[169]  (
    .HI(HI[169]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[16]  (
    .HI(HI[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[170]  (
    .HI(HI[170]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[171]  (
    .HI(HI[171]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[172]  (
    .HI(HI[172]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[173]  (
    .HI(HI[173]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[174]  (
    .HI(HI[174]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[175]  (
    .HI(HI[175]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[176]  (
    .HI(HI[176]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[177]  (
    .HI(HI[177]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[178]  (
    .HI(HI[178]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[179]  (
    .HI(HI[179]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[17]  (
    .HI(HI[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[180]  (
    .HI(HI[180]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[181]  (
    .HI(HI[181]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[182]  (
    .HI(HI[182]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[183]  (
    .HI(HI[183]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[184]  (
    .HI(HI[184]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[185]  (
    .HI(HI[185]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[186]  (
    .HI(HI[186]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[187]  (
    .HI(HI[187]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[188]  (
    .HI(HI[188]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[189]  (
    .HI(HI[189]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[18]  (
    .HI(HI[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[190]  (
    .HI(HI[190]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[191]  (
    .HI(HI[191]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[192]  (
    .HI(HI[192]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[193]  (
    .HI(HI[193]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[194]  (
    .HI(HI[194]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[195]  (
    .HI(HI[195]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[196]  (
    .HI(HI[196]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[197]  (
    .HI(HI[197]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[198]  (
    .HI(HI[198]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[199]  (
    .HI(HI[199]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[19]  (
    .HI(HI[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[1]  (
    .HI(HI[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[200]  (
    .HI(HI[200]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[201]  (
    .HI(HI[201]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[202]  (
    .HI(HI[202]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[203]  (
    .HI(HI[203]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[204]  (
    .HI(HI[204]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[205]  (
    .HI(HI[205]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[206]  (
    .HI(HI[206]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[207]  (
    .HI(HI[207]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[208]  (
    .HI(HI[208]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[209]  (
    .HI(HI[209]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[20]  (
    .HI(HI[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[210]  (
    .HI(HI[210]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[211]  (
    .HI(HI[211]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[212]  (
    .HI(HI[212]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[213]  (
    .HI(HI[213]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[214]  (
    .HI(HI[214]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[215]  (
    .HI(HI[215]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[216]  (
    .HI(HI[216]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[217]  (
    .HI(HI[217]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[218]  (
    .HI(HI[218]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[219]  (
    .HI(HI[219]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[21]  (
    .HI(HI[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[220]  (
    .HI(HI[220]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[221]  (
    .HI(HI[221]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[222]  (
    .HI(HI[222]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[223]  (
    .HI(HI[223]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[224]  (
    .HI(HI[224]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[225]  (
    .HI(HI[225]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[226]  (
    .HI(HI[226]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[227]  (
    .HI(HI[227]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[228]  (
    .HI(HI[228]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[229]  (
    .HI(HI[229]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[22]  (
    .HI(HI[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[230]  (
    .HI(HI[230]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[231]  (
    .HI(HI[231]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[232]  (
    .HI(HI[232]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[233]  (
    .HI(HI[233]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[234]  (
    .HI(HI[234]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[235]  (
    .HI(HI[235]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[236]  (
    .HI(HI[236]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[237]  (
    .HI(HI[237]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[238]  (
    .HI(HI[238]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[239]  (
    .HI(HI[239]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[23]  (
    .HI(HI[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[240]  (
    .HI(HI[240]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[241]  (
    .HI(HI[241]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[242]  (
    .HI(HI[242]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[243]  (
    .HI(HI[243]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[244]  (
    .HI(HI[244]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[245]  (
    .HI(HI[245]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[246]  (
    .HI(HI[246]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[247]  (
    .HI(HI[247]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[248]  (
    .HI(HI[248]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[249]  (
    .HI(HI[249]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[24]  (
    .HI(HI[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[250]  (
    .HI(HI[250]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[251]  (
    .HI(HI[251]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[252]  (
    .HI(HI[252]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[253]  (
    .HI(HI[253]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[254]  (
    .HI(HI[254]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[255]  (
    .HI(HI[255]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[256]  (
    .HI(HI[256]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[257]  (
    .HI(HI[257]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[258]  (
    .HI(HI[258]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[259]  (
    .HI(HI[259]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[25]  (
    .HI(HI[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[260]  (
    .HI(HI[260]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[261]  (
    .HI(HI[261]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[262]  (
    .HI(HI[262]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[263]  (
    .HI(HI[263]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[264]  (
    .HI(HI[264]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[265]  (
    .HI(HI[265]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[266]  (
    .HI(HI[266]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[267]  (
    .HI(HI[267]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[268]  (
    .HI(HI[268]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[269]  (
    .HI(HI[269]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[26]  (
    .HI(HI[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[270]  (
    .HI(HI[270]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[271]  (
    .HI(HI[271]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[272]  (
    .HI(HI[272]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[273]  (
    .HI(HI[273]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[274]  (
    .HI(HI[274]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[275]  (
    .HI(HI[275]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[276]  (
    .HI(HI[276]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[277]  (
    .HI(HI[277]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[278]  (
    .HI(HI[278]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[279]  (
    .HI(HI[279]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[27]  (
    .HI(HI[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[280]  (
    .HI(HI[280]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[281]  (
    .HI(HI[281]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[282]  (
    .HI(HI[282]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[283]  (
    .HI(HI[283]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[284]  (
    .HI(HI[284]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[285]  (
    .HI(HI[285]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[286]  (
    .HI(HI[286]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[287]  (
    .HI(HI[287]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[288]  (
    .HI(HI[288]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[289]  (
    .HI(HI[289]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[28]  (
    .HI(HI[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[290]  (
    .HI(HI[290]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[291]  (
    .HI(HI[291]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[292]  (
    .HI(HI[292]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[293]  (
    .HI(HI[293]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[294]  (
    .HI(HI[294]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[295]  (
    .HI(HI[295]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[296]  (
    .HI(HI[296]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[297]  (
    .HI(HI[297]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[298]  (
    .HI(HI[298]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[299]  (
    .HI(HI[299]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[29]  (
    .HI(HI[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[2]  (
    .HI(HI[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[300]  (
    .HI(HI[300]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[301]  (
    .HI(HI[301]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[302]  (
    .HI(HI[302]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[303]  (
    .HI(HI[303]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[304]  (
    .HI(HI[304]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[305]  (
    .HI(HI[305]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[306]  (
    .HI(HI[306]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[307]  (
    .HI(HI[307]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[308]  (
    .HI(HI[308]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[309]  (
    .HI(HI[309]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[30]  (
    .HI(HI[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[310]  (
    .HI(HI[310]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[311]  (
    .HI(HI[311]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[312]  (
    .HI(HI[312]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[313]  (
    .HI(HI[313]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[314]  (
    .HI(HI[314]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[315]  (
    .HI(HI[315]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[316]  (
    .HI(HI[316]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[317]  (
    .HI(HI[317]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[318]  (
    .HI(HI[318]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[319]  (
    .HI(HI[319]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[31]  (
    .HI(HI[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[320]  (
    .HI(HI[320]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[321]  (
    .HI(HI[321]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[322]  (
    .HI(HI[322]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[323]  (
    .HI(HI[323]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[324]  (
    .HI(HI[324]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[325]  (
    .HI(HI[325]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[326]  (
    .HI(HI[326]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[327]  (
    .HI(HI[327]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[328]  (
    .HI(HI[328]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[329]  (
    .HI(HI[329]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[32]  (
    .HI(HI[32]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[330]  (
    .HI(HI[330]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[331]  (
    .HI(HI[331]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[332]  (
    .HI(HI[332]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[333]  (
    .HI(HI[333]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[334]  (
    .HI(HI[334]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[335]  (
    .HI(HI[335]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[336]  (
    .HI(HI[336]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[337]  (
    .HI(HI[337]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[338]  (
    .HI(HI[338]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[339]  (
    .HI(HI[339]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[33]  (
    .HI(HI[33]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[340]  (
    .HI(HI[340]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[341]  (
    .HI(HI[341]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[342]  (
    .HI(HI[342]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[343]  (
    .HI(HI[343]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[344]  (
    .HI(HI[344]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[345]  (
    .HI(HI[345]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[346]  (
    .HI(HI[346]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[347]  (
    .HI(HI[347]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[348]  (
    .HI(HI[348]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[349]  (
    .HI(HI[349]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[34]  (
    .HI(HI[34]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[350]  (
    .HI(HI[350]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[351]  (
    .HI(HI[351]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[352]  (
    .HI(HI[352]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[353]  (
    .HI(HI[353]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[354]  (
    .HI(HI[354]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[355]  (
    .HI(HI[355]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[356]  (
    .HI(HI[356]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[357]  (
    .HI(HI[357]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[358]  (
    .HI(HI[358]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[359]  (
    .HI(HI[359]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[35]  (
    .HI(HI[35]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[360]  (
    .HI(HI[360]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[361]  (
    .HI(HI[361]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[362]  (
    .HI(HI[362]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[363]  (
    .HI(HI[363]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[364]  (
    .HI(HI[364]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[365]  (
    .HI(HI[365]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[366]  (
    .HI(HI[366]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[367]  (
    .HI(HI[367]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[368]  (
    .HI(HI[368]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[369]  (
    .HI(HI[369]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[36]  (
    .HI(HI[36]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[370]  (
    .HI(HI[370]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[371]  (
    .HI(HI[371]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[372]  (
    .HI(HI[372]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[373]  (
    .HI(HI[373]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[374]  (
    .HI(HI[374]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[375]  (
    .HI(HI[375]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[376]  (
    .HI(HI[376]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[377]  (
    .HI(HI[377]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[378]  (
    .HI(HI[378]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[379]  (
    .HI(HI[379]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[37]  (
    .HI(HI[37]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[380]  (
    .HI(HI[380]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[381]  (
    .HI(HI[381]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[382]  (
    .HI(HI[382]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[383]  (
    .HI(HI[383]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[384]  (
    .HI(HI[384]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[385]  (
    .HI(HI[385]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[386]  (
    .HI(HI[386]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[387]  (
    .HI(HI[387]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[388]  (
    .HI(HI[388]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[389]  (
    .HI(HI[389]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[38]  (
    .HI(HI[38]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[390]  (
    .HI(HI[390]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[391]  (
    .HI(HI[391]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[392]  (
    .HI(HI[392]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[393]  (
    .HI(HI[393]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[394]  (
    .HI(HI[394]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[395]  (
    .HI(HI[395]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[396]  (
    .HI(HI[396]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[397]  (
    .HI(HI[397]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[398]  (
    .HI(HI[398]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[399]  (
    .HI(HI[399]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[39]  (
    .HI(HI[39]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[3]  (
    .HI(HI[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[400]  (
    .HI(HI[400]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[401]  (
    .HI(HI[401]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[402]  (
    .HI(HI[402]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[403]  (
    .HI(HI[403]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[404]  (
    .HI(HI[404]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[405]  (
    .HI(HI[405]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[406]  (
    .HI(HI[406]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[407]  (
    .HI(HI[407]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[408]  (
    .HI(HI[408]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[409]  (
    .HI(HI[409]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[40]  (
    .HI(HI[40]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[410]  (
    .HI(HI[410]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[411]  (
    .HI(HI[411]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[412]  (
    .HI(HI[412]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[413]  (
    .HI(HI[413]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[414]  (
    .HI(HI[414]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[415]  (
    .HI(HI[415]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[416]  (
    .HI(HI[416]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[417]  (
    .HI(HI[417]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[418]  (
    .HI(HI[418]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[419]  (
    .HI(HI[419]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[41]  (
    .HI(HI[41]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[420]  (
    .HI(HI[420]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[421]  (
    .HI(HI[421]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[422]  (
    .HI(HI[422]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[423]  (
    .HI(HI[423]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[424]  (
    .HI(HI[424]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[425]  (
    .HI(HI[425]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[426]  (
    .HI(HI[426]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[427]  (
    .HI(HI[427]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[428]  (
    .HI(HI[428]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[429]  (
    .HI(HI[429]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[42]  (
    .HI(HI[42]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[430]  (
    .HI(HI[430]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[431]  (
    .HI(HI[431]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[432]  (
    .HI(HI[432]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[433]  (
    .HI(HI[433]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[434]  (
    .HI(HI[434]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[435]  (
    .HI(HI[435]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[436]  (
    .HI(HI[436]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[437]  (
    .HI(HI[437]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[438]  (
    .HI(HI[438]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[439]  (
    .HI(HI[439]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[43]  (
    .HI(HI[43]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[440]  (
    .HI(HI[440]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[441]  (
    .HI(HI[441]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[442]  (
    .HI(HI[442]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[443]  (
    .HI(HI[443]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[444]  (
    .HI(HI[444]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[445]  (
    .HI(HI[445]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[446]  (
    .HI(HI[446]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[447]  (
    .HI(HI[447]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[448]  (
    .HI(HI[448]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[449]  (
    .HI(HI[449]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[44]  (
    .HI(HI[44]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[450]  (
    .HI(HI[450]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[451]  (
    .HI(HI[451]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[452]  (
    .HI(HI[452]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[453]  (
    .HI(HI[453]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[454]  (
    .HI(HI[454]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[455]  (
    .HI(HI[455]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[456]  (
    .HI(HI[456]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[457]  (
    .HI(HI[457]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[458]  (
    .HI(HI[458]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[45]  (
    .HI(HI[45]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[46]  (
    .HI(HI[46]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[47]  (
    .HI(HI[47]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[48]  (
    .HI(HI[48]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[49]  (
    .HI(HI[49]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[4]  (
    .HI(HI[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[50]  (
    .HI(HI[50]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[51]  (
    .HI(HI[51]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[52]  (
    .HI(HI[52]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[53]  (
    .HI(HI[53]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[54]  (
    .HI(HI[54]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[55]  (
    .HI(HI[55]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[56]  (
    .HI(HI[56]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[57]  (
    .HI(HI[57]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[58]  (
    .HI(HI[58]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[59]  (
    .HI(HI[59]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[5]  (
    .HI(HI[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[60]  (
    .HI(HI[60]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[61]  (
    .HI(HI[61]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[62]  (
    .HI(HI[62]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[63]  (
    .HI(HI[63]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[64]  (
    .HI(HI[64]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[65]  (
    .HI(HI[65]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[66]  (
    .HI(HI[66]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[67]  (
    .HI(HI[67]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[68]  (
    .HI(HI[68]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[69]  (
    .HI(HI[69]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[6]  (
    .HI(HI[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[70]  (
    .HI(HI[70]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[71]  (
    .HI(HI[71]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[72]  (
    .HI(HI[72]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[73]  (
    .HI(HI[73]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[74]  (
    .HI(HI[74]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[75]  (
    .HI(HI[75]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[76]  (
    .HI(HI[76]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[77]  (
    .HI(HI[77]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[78]  (
    .HI(HI[78]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[79]  (
    .HI(HI[79]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[7]  (
    .HI(HI[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[80]  (
    .HI(HI[80]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[81]  (
    .HI(HI[81]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[82]  (
    .HI(HI[82]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[83]  (
    .HI(HI[83]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[84]  (
    .HI(HI[84]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[85]  (
    .HI(HI[85]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[86]  (
    .HI(HI[86]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[87]  (
    .HI(HI[87]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[88]  (
    .HI(HI[88]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[89]  (
    .HI(HI[89]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[8]  (
    .HI(HI[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[90]  (
    .HI(HI[90]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[91]  (
    .HI(HI[91]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[92]  (
    .HI(HI[92]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[93]  (
    .HI(HI[93]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[94]  (
    .HI(HI[94]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[95]  (
    .HI(HI[95]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[96]  (
    .HI(HI[96]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[97]  (
    .HI(HI[97]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[98]  (
    .HI(HI[98]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[99]  (
    .HI(HI[99]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
  sky130_fd_sc_hd__conb_1 \insts[9]  (
    .HI(HI[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1)
  );
endmodule
